module cla_52bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add1[19], i_add1[20], i_add1[21], i_add1[22], i_add1[23], i_add1[24], i_add1[25], i_add1[26], i_add1[27], i_add1[28], i_add1[29], i_add1[30], i_add1[31], i_add1[32], i_add1[33], i_add1[34], i_add1[35], i_add1[36], i_add1[37], i_add1[38], i_add1[39], i_add1[40], i_add1[41], i_add1[42], i_add1[43], i_add1[44], i_add1[45], i_add1[46], i_add1[47], i_add1[48], i_add1[49], i_add1[50], i_add1[51], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], i_add2[19], i_add2[20], i_add2[21], i_add2[22], i_add2[23], i_add2[24], i_add2[25], i_add2[26], i_add2[27], i_add2[28], i_add2[29], i_add2[30], i_add2[31], i_add2[32], i_add2[33], i_add2[34], i_add2[35], i_add2[36], i_add2[37], i_add2[38], i_add2[39], i_add2[40], i_add2[41], i_add2[42], i_add2[43], i_add2[44], i_add2[45], i_add2[46], i_add2[47], i_add2[48], i_add2[49], i_add2[50], i_add2[51], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21], o_result[22], o_result[23], o_result[24], o_result[25], o_result[26], o_result[27], o_result[28], o_result[29], o_result[30], o_result[31], o_result[32], o_result[33], o_result[34], o_result[35], o_result[36], o_result[37], o_result[38], o_result[39], o_result[40], o_result[41], o_result[42], o_result[43], o_result[44], o_result[45], o_result[46], o_result[47], o_result[48], o_result[49], o_result[50], o_result[51], o_result[52]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add1[19];
input i_add1[20];
input i_add1[21];
input i_add1[22];
input i_add1[23];
input i_add1[24];
input i_add1[25];
input i_add1[26];
input i_add1[27];
input i_add1[28];
input i_add1[29];
input i_add1[30];
input i_add1[31];
input i_add1[32];
input i_add1[33];
input i_add1[34];
input i_add1[35];
input i_add1[36];
input i_add1[37];
input i_add1[38];
input i_add1[39];
input i_add1[40];
input i_add1[41];
input i_add1[42];
input i_add1[43];
input i_add1[44];
input i_add1[45];
input i_add1[46];
input i_add1[47];
input i_add1[48];
input i_add1[49];
input i_add1[50];
input i_add1[51];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
input i_add2[19];
input i_add2[20];
input i_add2[21];
input i_add2[22];
input i_add2[23];
input i_add2[24];
input i_add2[25];
input i_add2[26];
input i_add2[27];
input i_add2[28];
input i_add2[29];
input i_add2[30];
input i_add2[31];
input i_add2[32];
input i_add2[33];
input i_add2[34];
input i_add2[35];
input i_add2[36];
input i_add2[37];
input i_add2[38];
input i_add2[39];
input i_add2[40];
input i_add2[41];
input i_add2[42];
input i_add2[43];
input i_add2[44];
input i_add2[45];
input i_add2[46];
input i_add2[47];
input i_add2[48];
input i_add2[49];
input i_add2[50];
input i_add2[51];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];
output o_result[22];
output o_result[23];
output o_result[24];
output o_result[25];
output o_result[26];
output o_result[27];
output o_result[28];
output o_result[29];
output o_result[30];
output o_result[31];
output o_result[32];
output o_result[33];
output o_result[34];
output o_result[35];
output o_result[36];
output o_result[37];
output o_result[38];
output o_result[39];
output o_result[40];
output o_result[41];
output o_result[42];
output o_result[43];
output o_result[44];
output o_result[45];
output o_result[46];
output o_result[47];
output o_result[48];
output o_result[49];
output o_result[50];
output o_result[51];
output o_result[52];

INVX1 INVX1_1 ( .A(_127_), .Y(_128_) );
NAND3X1 NAND3X1_1 ( .A(_126_), .B(_128_), .C(_119_), .Y(_129_) );
AND2X2 AND2X2_1 ( .A(_129_), .B(_124_), .Y(_130_) );
INVX1 INVX1_2 ( .A(_130_), .Y(w_C_22_) );
AND2X2 AND2X2_2 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_131_) );
INVX1 INVX1_3 ( .A(_131_), .Y(_132_) );
NAND3X1 NAND3X1_2 ( .A(_124_), .B(_132_), .C(_129_), .Y(_133_) );
OAI21X1 OAI21X1_1 ( .A(i_add2[22]), .B(i_add1[22]), .C(_133_), .Y(_134_) );
INVX1 INVX1_4 ( .A(_134_), .Y(w_C_23_) );
INVX1 INVX1_5 ( .A(i_add2[23]), .Y(_135_) );
INVX1 INVX1_6 ( .A(i_add1[23]), .Y(_136_) );
NOR2X1 NOR2X1_1 ( .A(_135_), .B(_136_), .Y(_137_) );
INVX1 INVX1_7 ( .A(_137_), .Y(_138_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_139_) );
INVX1 INVX1_8 ( .A(_139_), .Y(_140_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_141_) );
INVX1 INVX1_9 ( .A(_141_), .Y(_142_) );
NAND3X1 NAND3X1_3 ( .A(_140_), .B(_142_), .C(_133_), .Y(_143_) );
AND2X2 AND2X2_3 ( .A(_143_), .B(_138_), .Y(_144_) );
INVX1 INVX1_10 ( .A(_144_), .Y(w_C_24_) );
AND2X2 AND2X2_4 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_145_) );
INVX1 INVX1_11 ( .A(_145_), .Y(_146_) );
NAND3X1 NAND3X1_4 ( .A(_138_), .B(_146_), .C(_143_), .Y(_147_) );
OAI21X1 OAI21X1_2 ( .A(i_add2[24]), .B(i_add1[24]), .C(_147_), .Y(_148_) );
INVX1 INVX1_12 ( .A(_148_), .Y(w_C_25_) );
INVX1 INVX1_13 ( .A(i_add2[25]), .Y(_149_) );
INVX1 INVX1_14 ( .A(i_add1[25]), .Y(_150_) );
NOR2X1 NOR2X1_4 ( .A(_149_), .B(_150_), .Y(_151_) );
INVX1 INVX1_15 ( .A(_151_), .Y(_152_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_153_) );
INVX1 INVX1_16 ( .A(_153_), .Y(_154_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_155_) );
INVX1 INVX1_17 ( .A(_155_), .Y(_156_) );
NAND3X1 NAND3X1_5 ( .A(_154_), .B(_156_), .C(_147_), .Y(_157_) );
AND2X2 AND2X2_5 ( .A(_157_), .B(_152_), .Y(_158_) );
INVX1 INVX1_18 ( .A(_158_), .Y(w_C_26_) );
AND2X2 AND2X2_6 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_159_) );
INVX1 INVX1_19 ( .A(_159_), .Y(_160_) );
NAND3X1 NAND3X1_6 ( .A(_152_), .B(_160_), .C(_157_), .Y(_161_) );
OAI21X1 OAI21X1_3 ( .A(i_add2[26]), .B(i_add1[26]), .C(_161_), .Y(_162_) );
INVX1 INVX1_20 ( .A(_162_), .Y(w_C_27_) );
INVX1 INVX1_21 ( .A(i_add2[27]), .Y(_163_) );
INVX1 INVX1_22 ( .A(i_add1[27]), .Y(_164_) );
NOR2X1 NOR2X1_7 ( .A(_163_), .B(_164_), .Y(_165_) );
INVX1 INVX1_23 ( .A(_165_), .Y(_166_) );
BUFX2 BUFX2_1 ( .A(_314__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_314__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_314__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_314__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_314__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_314__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_314__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_314__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_314__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_314__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_314__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_314__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_314__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_314__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_314__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_314__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_314__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_314__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_314__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_314__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_314__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_314__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_314__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_314__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_314__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_314__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_314__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_314__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_314__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_314__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_314__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_314__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_314__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_314__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_314__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_314__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_314__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(_314__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .A(_314__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .A(_314__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .A(_314__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .A(_314__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .A(_314__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .A(_314__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .A(_314__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .A(_314__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .A(_314__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .A(_314__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .A(_314__48_), .Y(o_result[48]) );
BUFX2 BUFX2_50 ( .A(_314__49_), .Y(o_result[49]) );
BUFX2 BUFX2_51 ( .A(_314__50_), .Y(o_result[50]) );
BUFX2 BUFX2_52 ( .A(_314__51_), .Y(o_result[51]) );
BUFX2 BUFX2_53 ( .A(w_C_52_), .Y(o_result[52]) );
INVX1 INVX1_24 ( .A(w_C_4_), .Y(_318_) );
OR2X2 OR2X2_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_319_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_320_) );
NAND3X1 NAND3X1_7 ( .A(_318_), .B(_320_), .C(_319_), .Y(_321_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_315_) );
AND2X2 AND2X2_7 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_316_) );
OAI21X1 OAI21X1_4 ( .A(_315_), .B(_316_), .C(w_C_4_), .Y(_317_) );
NAND2X1 NAND2X1_2 ( .A(_317_), .B(_321_), .Y(_314__4_) );
INVX1 INVX1_25 ( .A(w_C_5_), .Y(_325_) );
OR2X2 OR2X2_2 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_326_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_327_) );
NAND3X1 NAND3X1_8 ( .A(_325_), .B(_327_), .C(_326_), .Y(_328_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_322_) );
AND2X2 AND2X2_8 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_323_) );
OAI21X1 OAI21X1_5 ( .A(_322_), .B(_323_), .C(w_C_5_), .Y(_324_) );
NAND2X1 NAND2X1_4 ( .A(_324_), .B(_328_), .Y(_314__5_) );
INVX1 INVX1_26 ( .A(w_C_6_), .Y(_332_) );
OR2X2 OR2X2_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_333_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_334_) );
NAND3X1 NAND3X1_9 ( .A(_332_), .B(_334_), .C(_333_), .Y(_335_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_329_) );
AND2X2 AND2X2_9 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_330_) );
OAI21X1 OAI21X1_6 ( .A(_329_), .B(_330_), .C(w_C_6_), .Y(_331_) );
NAND2X1 NAND2X1_6 ( .A(_331_), .B(_335_), .Y(_314__6_) );
INVX1 INVX1_27 ( .A(w_C_7_), .Y(_339_) );
OR2X2 OR2X2_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_340_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_341_) );
NAND3X1 NAND3X1_10 ( .A(_339_), .B(_341_), .C(_340_), .Y(_342_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_336_) );
AND2X2 AND2X2_10 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_337_) );
OAI21X1 OAI21X1_7 ( .A(_336_), .B(_337_), .C(w_C_7_), .Y(_338_) );
NAND2X1 NAND2X1_8 ( .A(_338_), .B(_342_), .Y(_314__7_) );
INVX1 INVX1_28 ( .A(w_C_8_), .Y(_346_) );
OR2X2 OR2X2_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_347_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_348_) );
NAND3X1 NAND3X1_11 ( .A(_346_), .B(_348_), .C(_347_), .Y(_349_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_343_) );
AND2X2 AND2X2_11 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_344_) );
OAI21X1 OAI21X1_8 ( .A(_343_), .B(_344_), .C(w_C_8_), .Y(_345_) );
NAND2X1 NAND2X1_10 ( .A(_345_), .B(_349_), .Y(_314__8_) );
INVX1 INVX1_29 ( .A(w_C_9_), .Y(_353_) );
OR2X2 OR2X2_6 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_354_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_355_) );
NAND3X1 NAND3X1_12 ( .A(_353_), .B(_355_), .C(_354_), .Y(_356_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_350_) );
AND2X2 AND2X2_12 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_351_) );
OAI21X1 OAI21X1_9 ( .A(_350_), .B(_351_), .C(w_C_9_), .Y(_352_) );
NAND2X1 NAND2X1_12 ( .A(_352_), .B(_356_), .Y(_314__9_) );
INVX1 INVX1_30 ( .A(w_C_10_), .Y(_360_) );
OR2X2 OR2X2_7 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_361_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_362_) );
NAND3X1 NAND3X1_13 ( .A(_360_), .B(_362_), .C(_361_), .Y(_363_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_357_) );
AND2X2 AND2X2_13 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_358_) );
OAI21X1 OAI21X1_10 ( .A(_357_), .B(_358_), .C(w_C_10_), .Y(_359_) );
NAND2X1 NAND2X1_14 ( .A(_359_), .B(_363_), .Y(_314__10_) );
INVX1 INVX1_31 ( .A(w_C_11_), .Y(_367_) );
OR2X2 OR2X2_8 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_368_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_369_) );
NAND3X1 NAND3X1_14 ( .A(_367_), .B(_369_), .C(_368_), .Y(_370_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_364_) );
AND2X2 AND2X2_14 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_365_) );
OAI21X1 OAI21X1_11 ( .A(_364_), .B(_365_), .C(w_C_11_), .Y(_366_) );
NAND2X1 NAND2X1_16 ( .A(_366_), .B(_370_), .Y(_314__11_) );
INVX1 INVX1_32 ( .A(w_C_12_), .Y(_374_) );
OR2X2 OR2X2_9 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_375_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_376_) );
NAND3X1 NAND3X1_15 ( .A(_374_), .B(_376_), .C(_375_), .Y(_377_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_371_) );
AND2X2 AND2X2_15 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_372_) );
OAI21X1 OAI21X1_12 ( .A(_371_), .B(_372_), .C(w_C_12_), .Y(_373_) );
NAND2X1 NAND2X1_18 ( .A(_373_), .B(_377_), .Y(_314__12_) );
INVX1 INVX1_33 ( .A(w_C_13_), .Y(_381_) );
OR2X2 OR2X2_10 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_382_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_383_) );
NAND3X1 NAND3X1_16 ( .A(_381_), .B(_383_), .C(_382_), .Y(_384_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_378_) );
AND2X2 AND2X2_16 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_379_) );
OAI21X1 OAI21X1_13 ( .A(_378_), .B(_379_), .C(w_C_13_), .Y(_380_) );
NAND2X1 NAND2X1_20 ( .A(_380_), .B(_384_), .Y(_314__13_) );
INVX1 INVX1_34 ( .A(w_C_14_), .Y(_388_) );
OR2X2 OR2X2_11 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_389_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_390_) );
NAND3X1 NAND3X1_17 ( .A(_388_), .B(_390_), .C(_389_), .Y(_391_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_385_) );
AND2X2 AND2X2_17 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_386_) );
OAI21X1 OAI21X1_14 ( .A(_385_), .B(_386_), .C(w_C_14_), .Y(_387_) );
NAND2X1 NAND2X1_22 ( .A(_387_), .B(_391_), .Y(_314__14_) );
INVX1 INVX1_35 ( .A(w_C_15_), .Y(_395_) );
OR2X2 OR2X2_12 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_396_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_397_) );
NAND3X1 NAND3X1_18 ( .A(_395_), .B(_397_), .C(_396_), .Y(_398_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_392_) );
AND2X2 AND2X2_18 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_393_) );
OAI21X1 OAI21X1_15 ( .A(_392_), .B(_393_), .C(w_C_15_), .Y(_394_) );
NAND2X1 NAND2X1_24 ( .A(_394_), .B(_398_), .Y(_314__15_) );
INVX1 INVX1_36 ( .A(w_C_16_), .Y(_402_) );
OR2X2 OR2X2_13 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_403_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_404_) );
NAND3X1 NAND3X1_19 ( .A(_402_), .B(_404_), .C(_403_), .Y(_405_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_399_) );
AND2X2 AND2X2_19 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_400_) );
OAI21X1 OAI21X1_16 ( .A(_399_), .B(_400_), .C(w_C_16_), .Y(_401_) );
NAND2X1 NAND2X1_26 ( .A(_401_), .B(_405_), .Y(_314__16_) );
INVX1 INVX1_37 ( .A(w_C_17_), .Y(_409_) );
OR2X2 OR2X2_14 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_410_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_411_) );
NAND3X1 NAND3X1_20 ( .A(_409_), .B(_411_), .C(_410_), .Y(_412_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_406_) );
AND2X2 AND2X2_20 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_407_) );
OAI21X1 OAI21X1_17 ( .A(_406_), .B(_407_), .C(w_C_17_), .Y(_408_) );
NAND2X1 NAND2X1_28 ( .A(_408_), .B(_412_), .Y(_314__17_) );
INVX1 INVX1_38 ( .A(w_C_18_), .Y(_416_) );
OR2X2 OR2X2_15 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_417_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_418_) );
NAND3X1 NAND3X1_21 ( .A(_416_), .B(_418_), .C(_417_), .Y(_419_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_413_) );
AND2X2 AND2X2_21 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_414_) );
OAI21X1 OAI21X1_18 ( .A(_413_), .B(_414_), .C(w_C_18_), .Y(_415_) );
NAND2X1 NAND2X1_30 ( .A(_415_), .B(_419_), .Y(_314__18_) );
INVX1 INVX1_39 ( .A(w_C_19_), .Y(_423_) );
OR2X2 OR2X2_16 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_424_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_425_) );
NAND3X1 NAND3X1_22 ( .A(_423_), .B(_425_), .C(_424_), .Y(_426_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_420_) );
AND2X2 AND2X2_22 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_421_) );
OAI21X1 OAI21X1_19 ( .A(_420_), .B(_421_), .C(w_C_19_), .Y(_422_) );
NAND2X1 NAND2X1_32 ( .A(_422_), .B(_426_), .Y(_314__19_) );
INVX1 INVX1_40 ( .A(w_C_20_), .Y(_430_) );
OR2X2 OR2X2_17 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_431_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_432_) );
NAND3X1 NAND3X1_23 ( .A(_430_), .B(_432_), .C(_431_), .Y(_433_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_427_) );
AND2X2 AND2X2_23 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_428_) );
OAI21X1 OAI21X1_20 ( .A(_427_), .B(_428_), .C(w_C_20_), .Y(_429_) );
NAND2X1 NAND2X1_34 ( .A(_429_), .B(_433_), .Y(_314__20_) );
INVX1 INVX1_41 ( .A(w_C_21_), .Y(_437_) );
OR2X2 OR2X2_18 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_438_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_439_) );
NAND3X1 NAND3X1_24 ( .A(_437_), .B(_439_), .C(_438_), .Y(_440_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_434_) );
AND2X2 AND2X2_24 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_435_) );
OAI21X1 OAI21X1_21 ( .A(_434_), .B(_435_), .C(w_C_21_), .Y(_436_) );
NAND2X1 NAND2X1_36 ( .A(_436_), .B(_440_), .Y(_314__21_) );
INVX1 INVX1_42 ( .A(w_C_22_), .Y(_444_) );
OR2X2 OR2X2_19 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_445_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_446_) );
NAND3X1 NAND3X1_25 ( .A(_444_), .B(_446_), .C(_445_), .Y(_447_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_441_) );
AND2X2 AND2X2_25 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_442_) );
OAI21X1 OAI21X1_22 ( .A(_441_), .B(_442_), .C(w_C_22_), .Y(_443_) );
NAND2X1 NAND2X1_38 ( .A(_443_), .B(_447_), .Y(_314__22_) );
INVX1 INVX1_43 ( .A(w_C_23_), .Y(_451_) );
OR2X2 OR2X2_20 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_452_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_453_) );
NAND3X1 NAND3X1_26 ( .A(_451_), .B(_453_), .C(_452_), .Y(_454_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_448_) );
AND2X2 AND2X2_26 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_449_) );
OAI21X1 OAI21X1_23 ( .A(_448_), .B(_449_), .C(w_C_23_), .Y(_450_) );
NAND2X1 NAND2X1_40 ( .A(_450_), .B(_454_), .Y(_314__23_) );
INVX1 INVX1_44 ( .A(w_C_24_), .Y(_458_) );
OR2X2 OR2X2_21 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_459_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_460_) );
NAND3X1 NAND3X1_27 ( .A(_458_), .B(_460_), .C(_459_), .Y(_461_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_455_) );
AND2X2 AND2X2_27 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_456_) );
OAI21X1 OAI21X1_24 ( .A(_455_), .B(_456_), .C(w_C_24_), .Y(_457_) );
NAND2X1 NAND2X1_42 ( .A(_457_), .B(_461_), .Y(_314__24_) );
INVX1 INVX1_45 ( .A(w_C_25_), .Y(_465_) );
OR2X2 OR2X2_22 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_466_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_467_) );
NAND3X1 NAND3X1_28 ( .A(_465_), .B(_467_), .C(_466_), .Y(_468_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_462_) );
AND2X2 AND2X2_28 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_463_) );
OAI21X1 OAI21X1_25 ( .A(_462_), .B(_463_), .C(w_C_25_), .Y(_464_) );
NAND2X1 NAND2X1_44 ( .A(_464_), .B(_468_), .Y(_314__25_) );
INVX1 INVX1_46 ( .A(w_C_26_), .Y(_472_) );
OR2X2 OR2X2_23 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_473_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_474_) );
NAND3X1 NAND3X1_29 ( .A(_472_), .B(_474_), .C(_473_), .Y(_475_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_469_) );
AND2X2 AND2X2_29 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_470_) );
OAI21X1 OAI21X1_26 ( .A(_469_), .B(_470_), .C(w_C_26_), .Y(_471_) );
NAND2X1 NAND2X1_46 ( .A(_471_), .B(_475_), .Y(_314__26_) );
INVX1 INVX1_47 ( .A(w_C_27_), .Y(_479_) );
OR2X2 OR2X2_24 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_480_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_481_) );
NAND3X1 NAND3X1_30 ( .A(_479_), .B(_481_), .C(_480_), .Y(_482_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_476_) );
AND2X2 AND2X2_30 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_477_) );
OAI21X1 OAI21X1_27 ( .A(_476_), .B(_477_), .C(w_C_27_), .Y(_478_) );
NAND2X1 NAND2X1_48 ( .A(_478_), .B(_482_), .Y(_314__27_) );
INVX1 INVX1_48 ( .A(w_C_28_), .Y(_486_) );
OR2X2 OR2X2_25 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_487_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_488_) );
NAND3X1 NAND3X1_31 ( .A(_486_), .B(_488_), .C(_487_), .Y(_489_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_483_) );
AND2X2 AND2X2_31 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_484_) );
OAI21X1 OAI21X1_28 ( .A(_483_), .B(_484_), .C(w_C_28_), .Y(_485_) );
NAND2X1 NAND2X1_50 ( .A(_485_), .B(_489_), .Y(_314__28_) );
INVX1 INVX1_49 ( .A(w_C_29_), .Y(_493_) );
OR2X2 OR2X2_26 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_494_) );
NAND2X1 NAND2X1_51 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_495_) );
NAND3X1 NAND3X1_32 ( .A(_493_), .B(_495_), .C(_494_), .Y(_496_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_490_) );
AND2X2 AND2X2_32 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_491_) );
OAI21X1 OAI21X1_29 ( .A(_490_), .B(_491_), .C(w_C_29_), .Y(_492_) );
NAND2X1 NAND2X1_52 ( .A(_492_), .B(_496_), .Y(_314__29_) );
INVX1 INVX1_50 ( .A(w_C_30_), .Y(_500_) );
OR2X2 OR2X2_27 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_501_) );
NAND2X1 NAND2X1_53 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_502_) );
NAND3X1 NAND3X1_33 ( .A(_500_), .B(_502_), .C(_501_), .Y(_503_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_497_) );
AND2X2 AND2X2_33 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_498_) );
OAI21X1 OAI21X1_30 ( .A(_497_), .B(_498_), .C(w_C_30_), .Y(_499_) );
NAND2X1 NAND2X1_54 ( .A(_499_), .B(_503_), .Y(_314__30_) );
INVX1 INVX1_51 ( .A(w_C_31_), .Y(_507_) );
OR2X2 OR2X2_28 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_508_) );
NAND2X1 NAND2X1_55 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_509_) );
NAND3X1 NAND3X1_34 ( .A(_507_), .B(_509_), .C(_508_), .Y(_510_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_504_) );
AND2X2 AND2X2_34 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_505_) );
OAI21X1 OAI21X1_31 ( .A(_504_), .B(_505_), .C(w_C_31_), .Y(_506_) );
NAND2X1 NAND2X1_56 ( .A(_506_), .B(_510_), .Y(_314__31_) );
INVX1 INVX1_52 ( .A(w_C_32_), .Y(_514_) );
OR2X2 OR2X2_29 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_515_) );
NAND2X1 NAND2X1_57 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_516_) );
NAND3X1 NAND3X1_35 ( .A(_514_), .B(_516_), .C(_515_), .Y(_517_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_511_) );
AND2X2 AND2X2_35 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_512_) );
OAI21X1 OAI21X1_32 ( .A(_511_), .B(_512_), .C(w_C_32_), .Y(_513_) );
NAND2X1 NAND2X1_58 ( .A(_513_), .B(_517_), .Y(_314__32_) );
INVX1 INVX1_53 ( .A(w_C_33_), .Y(_521_) );
OR2X2 OR2X2_30 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_522_) );
NAND2X1 NAND2X1_59 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_523_) );
NAND3X1 NAND3X1_36 ( .A(_521_), .B(_523_), .C(_522_), .Y(_524_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_518_) );
AND2X2 AND2X2_36 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_519_) );
OAI21X1 OAI21X1_33 ( .A(_518_), .B(_519_), .C(w_C_33_), .Y(_520_) );
NAND2X1 NAND2X1_60 ( .A(_520_), .B(_524_), .Y(_314__33_) );
INVX1 INVX1_54 ( .A(w_C_34_), .Y(_528_) );
OR2X2 OR2X2_31 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_529_) );
NAND2X1 NAND2X1_61 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_530_) );
NAND3X1 NAND3X1_37 ( .A(_528_), .B(_530_), .C(_529_), .Y(_531_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_525_) );
AND2X2 AND2X2_37 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_526_) );
OAI21X1 OAI21X1_34 ( .A(_525_), .B(_526_), .C(w_C_34_), .Y(_527_) );
NAND2X1 NAND2X1_62 ( .A(_527_), .B(_531_), .Y(_314__34_) );
INVX1 INVX1_55 ( .A(w_C_35_), .Y(_535_) );
OR2X2 OR2X2_32 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_536_) );
NAND2X1 NAND2X1_63 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_537_) );
NAND3X1 NAND3X1_38 ( .A(_535_), .B(_537_), .C(_536_), .Y(_538_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_532_) );
AND2X2 AND2X2_38 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_533_) );
OAI21X1 OAI21X1_35 ( .A(_532_), .B(_533_), .C(w_C_35_), .Y(_534_) );
NAND2X1 NAND2X1_64 ( .A(_534_), .B(_538_), .Y(_314__35_) );
INVX1 INVX1_56 ( .A(w_C_36_), .Y(_542_) );
OR2X2 OR2X2_33 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_543_) );
NAND2X1 NAND2X1_65 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_544_) );
NAND3X1 NAND3X1_39 ( .A(_542_), .B(_544_), .C(_543_), .Y(_545_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_539_) );
AND2X2 AND2X2_39 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_540_) );
OAI21X1 OAI21X1_36 ( .A(_539_), .B(_540_), .C(w_C_36_), .Y(_541_) );
NAND2X1 NAND2X1_66 ( .A(_541_), .B(_545_), .Y(_314__36_) );
INVX1 INVX1_57 ( .A(w_C_37_), .Y(_549_) );
OR2X2 OR2X2_34 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_550_) );
NAND2X1 NAND2X1_67 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_551_) );
NAND3X1 NAND3X1_40 ( .A(_549_), .B(_551_), .C(_550_), .Y(_552_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_546_) );
AND2X2 AND2X2_40 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_547_) );
OAI21X1 OAI21X1_37 ( .A(_546_), .B(_547_), .C(w_C_37_), .Y(_548_) );
NAND2X1 NAND2X1_68 ( .A(_548_), .B(_552_), .Y(_314__37_) );
INVX1 INVX1_58 ( .A(w_C_38_), .Y(_556_) );
OR2X2 OR2X2_35 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_557_) );
NAND2X1 NAND2X1_69 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_558_) );
NAND3X1 NAND3X1_41 ( .A(_556_), .B(_558_), .C(_557_), .Y(_559_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_553_) );
AND2X2 AND2X2_41 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_554_) );
OAI21X1 OAI21X1_38 ( .A(_553_), .B(_554_), .C(w_C_38_), .Y(_555_) );
NAND2X1 NAND2X1_70 ( .A(_555_), .B(_559_), .Y(_314__38_) );
INVX1 INVX1_59 ( .A(w_C_39_), .Y(_563_) );
OR2X2 OR2X2_36 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_564_) );
NAND2X1 NAND2X1_71 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_565_) );
NAND3X1 NAND3X1_42 ( .A(_563_), .B(_565_), .C(_564_), .Y(_566_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_560_) );
AND2X2 AND2X2_42 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_561_) );
OAI21X1 OAI21X1_39 ( .A(_560_), .B(_561_), .C(w_C_39_), .Y(_562_) );
NAND2X1 NAND2X1_72 ( .A(_562_), .B(_566_), .Y(_314__39_) );
INVX1 INVX1_60 ( .A(w_C_40_), .Y(_570_) );
OR2X2 OR2X2_37 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_571_) );
NAND2X1 NAND2X1_73 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_572_) );
NAND3X1 NAND3X1_43 ( .A(_570_), .B(_572_), .C(_571_), .Y(_573_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_567_) );
AND2X2 AND2X2_43 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_568_) );
OAI21X1 OAI21X1_40 ( .A(_567_), .B(_568_), .C(w_C_40_), .Y(_569_) );
NAND2X1 NAND2X1_74 ( .A(_569_), .B(_573_), .Y(_314__40_) );
INVX1 INVX1_61 ( .A(w_C_41_), .Y(_577_) );
OR2X2 OR2X2_38 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_578_) );
NAND2X1 NAND2X1_75 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_579_) );
NAND3X1 NAND3X1_44 ( .A(_577_), .B(_579_), .C(_578_), .Y(_580_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_574_) );
AND2X2 AND2X2_44 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_575_) );
OAI21X1 OAI21X1_41 ( .A(_574_), .B(_575_), .C(w_C_41_), .Y(_576_) );
NAND2X1 NAND2X1_76 ( .A(_576_), .B(_580_), .Y(_314__41_) );
INVX1 INVX1_62 ( .A(w_C_42_), .Y(_584_) );
OR2X2 OR2X2_39 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_585_) );
NAND2X1 NAND2X1_77 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_586_) );
NAND3X1 NAND3X1_45 ( .A(_584_), .B(_586_), .C(_585_), .Y(_587_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_581_) );
AND2X2 AND2X2_45 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_582_) );
OAI21X1 OAI21X1_42 ( .A(_581_), .B(_582_), .C(w_C_42_), .Y(_583_) );
NAND2X1 NAND2X1_78 ( .A(_583_), .B(_587_), .Y(_314__42_) );
INVX1 INVX1_63 ( .A(w_C_43_), .Y(_591_) );
OR2X2 OR2X2_40 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_592_) );
NAND2X1 NAND2X1_79 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_593_) );
NAND3X1 NAND3X1_46 ( .A(_591_), .B(_593_), .C(_592_), .Y(_594_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_588_) );
AND2X2 AND2X2_46 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_589_) );
OAI21X1 OAI21X1_43 ( .A(_588_), .B(_589_), .C(w_C_43_), .Y(_590_) );
NAND2X1 NAND2X1_80 ( .A(_590_), .B(_594_), .Y(_314__43_) );
INVX1 INVX1_64 ( .A(w_C_44_), .Y(_598_) );
OR2X2 OR2X2_41 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_599_) );
NAND2X1 NAND2X1_81 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_600_) );
NAND3X1 NAND3X1_47 ( .A(_598_), .B(_600_), .C(_599_), .Y(_601_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_595_) );
AND2X2 AND2X2_47 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_596_) );
OAI21X1 OAI21X1_44 ( .A(_595_), .B(_596_), .C(w_C_44_), .Y(_597_) );
NAND2X1 NAND2X1_82 ( .A(_597_), .B(_601_), .Y(_314__44_) );
INVX1 INVX1_65 ( .A(w_C_45_), .Y(_605_) );
OR2X2 OR2X2_42 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_606_) );
NAND2X1 NAND2X1_83 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_607_) );
NAND3X1 NAND3X1_48 ( .A(_605_), .B(_607_), .C(_606_), .Y(_608_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_602_) );
AND2X2 AND2X2_48 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_603_) );
OAI21X1 OAI21X1_45 ( .A(_602_), .B(_603_), .C(w_C_45_), .Y(_604_) );
NAND2X1 NAND2X1_84 ( .A(_604_), .B(_608_), .Y(_314__45_) );
INVX1 INVX1_66 ( .A(w_C_46_), .Y(_612_) );
OR2X2 OR2X2_43 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_613_) );
NAND2X1 NAND2X1_85 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_614_) );
NAND3X1 NAND3X1_49 ( .A(_612_), .B(_614_), .C(_613_), .Y(_615_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_609_) );
AND2X2 AND2X2_49 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_610_) );
OAI21X1 OAI21X1_46 ( .A(_609_), .B(_610_), .C(w_C_46_), .Y(_611_) );
NAND2X1 NAND2X1_86 ( .A(_611_), .B(_615_), .Y(_314__46_) );
INVX1 INVX1_67 ( .A(w_C_47_), .Y(_619_) );
OR2X2 OR2X2_44 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_620_) );
NAND2X1 NAND2X1_87 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_621_) );
NAND3X1 NAND3X1_50 ( .A(_619_), .B(_621_), .C(_620_), .Y(_622_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_616_) );
AND2X2 AND2X2_50 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_617_) );
OAI21X1 OAI21X1_47 ( .A(_616_), .B(_617_), .C(w_C_47_), .Y(_618_) );
NAND2X1 NAND2X1_88 ( .A(_618_), .B(_622_), .Y(_314__47_) );
INVX1 INVX1_68 ( .A(w_C_48_), .Y(_626_) );
OR2X2 OR2X2_45 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_627_) );
NAND2X1 NAND2X1_89 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_628_) );
NAND3X1 NAND3X1_51 ( .A(_626_), .B(_628_), .C(_627_), .Y(_629_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_623_) );
AND2X2 AND2X2_51 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_624_) );
OAI21X1 OAI21X1_48 ( .A(_623_), .B(_624_), .C(w_C_48_), .Y(_625_) );
NAND2X1 NAND2X1_90 ( .A(_625_), .B(_629_), .Y(_314__48_) );
INVX1 INVX1_69 ( .A(w_C_49_), .Y(_633_) );
OR2X2 OR2X2_46 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_634_) );
NAND2X1 NAND2X1_91 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_635_) );
NAND3X1 NAND3X1_52 ( .A(_633_), .B(_635_), .C(_634_), .Y(_636_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_630_) );
AND2X2 AND2X2_52 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_631_) );
OAI21X1 OAI21X1_49 ( .A(_630_), .B(_631_), .C(w_C_49_), .Y(_632_) );
NAND2X1 NAND2X1_92 ( .A(_632_), .B(_636_), .Y(_314__49_) );
INVX1 INVX1_70 ( .A(w_C_50_), .Y(_640_) );
OR2X2 OR2X2_47 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_641_) );
NAND2X1 NAND2X1_93 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_642_) );
NAND3X1 NAND3X1_53 ( .A(_640_), .B(_642_), .C(_641_), .Y(_643_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_637_) );
AND2X2 AND2X2_53 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_638_) );
OAI21X1 OAI21X1_50 ( .A(_637_), .B(_638_), .C(w_C_50_), .Y(_639_) );
NAND2X1 NAND2X1_94 ( .A(_639_), .B(_643_), .Y(_314__50_) );
INVX1 INVX1_71 ( .A(w_C_51_), .Y(_647_) );
OR2X2 OR2X2_48 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_648_) );
NAND2X1 NAND2X1_95 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_649_) );
NAND3X1 NAND3X1_54 ( .A(_647_), .B(_649_), .C(_648_), .Y(_650_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_644_) );
AND2X2 AND2X2_54 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_645_) );
OAI21X1 OAI21X1_51 ( .A(_644_), .B(_645_), .C(w_C_51_), .Y(_646_) );
NAND2X1 NAND2X1_96 ( .A(_646_), .B(_650_), .Y(_314__51_) );
INVX1 INVX1_72 ( .A(1'b0), .Y(_654_) );
OR2X2 OR2X2_49 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_655_) );
NAND2X1 NAND2X1_97 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_656_) );
NAND3X1 NAND3X1_55 ( .A(_654_), .B(_656_), .C(_655_), .Y(_657_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_651_) );
AND2X2 AND2X2_55 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_652_) );
OAI21X1 OAI21X1_52 ( .A(_651_), .B(_652_), .C(1'b0), .Y(_653_) );
NAND2X1 NAND2X1_98 ( .A(_653_), .B(_657_), .Y(_314__0_) );
INVX1 INVX1_73 ( .A(w_C_1_), .Y(_661_) );
OR2X2 OR2X2_50 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_662_) );
NAND2X1 NAND2X1_99 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_663_) );
NAND3X1 NAND3X1_56 ( .A(_661_), .B(_663_), .C(_662_), .Y(_664_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_658_) );
AND2X2 AND2X2_56 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_659_) );
OAI21X1 OAI21X1_53 ( .A(_658_), .B(_659_), .C(w_C_1_), .Y(_660_) );
NAND2X1 NAND2X1_100 ( .A(_660_), .B(_664_), .Y(_314__1_) );
INVX1 INVX1_74 ( .A(w_C_2_), .Y(_668_) );
OR2X2 OR2X2_51 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_669_) );
NAND2X1 NAND2X1_101 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_670_) );
NAND3X1 NAND3X1_57 ( .A(_668_), .B(_670_), .C(_669_), .Y(_671_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_665_) );
AND2X2 AND2X2_57 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_666_) );
OAI21X1 OAI21X1_54 ( .A(_665_), .B(_666_), .C(w_C_2_), .Y(_667_) );
NAND2X1 NAND2X1_102 ( .A(_667_), .B(_671_), .Y(_314__2_) );
INVX1 INVX1_75 ( .A(w_C_3_), .Y(_675_) );
OR2X2 OR2X2_52 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_676_) );
NAND2X1 NAND2X1_103 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_677_) );
NAND3X1 NAND3X1_58 ( .A(_675_), .B(_677_), .C(_676_), .Y(_678_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_672_) );
AND2X2 AND2X2_58 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_673_) );
OAI21X1 OAI21X1_55 ( .A(_672_), .B(_673_), .C(w_C_3_), .Y(_674_) );
NAND2X1 NAND2X1_104 ( .A(_674_), .B(_678_), .Y(_314__3_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_167_) );
INVX1 INVX1_76 ( .A(_167_), .Y(_168_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_169_) );
INVX1 INVX1_77 ( .A(_169_), .Y(_170_) );
NAND3X1 NAND3X1_59 ( .A(_168_), .B(_170_), .C(_161_), .Y(_171_) );
AND2X2 AND2X2_59 ( .A(_171_), .B(_166_), .Y(_172_) );
INVX1 INVX1_78 ( .A(_172_), .Y(w_C_28_) );
AND2X2 AND2X2_60 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_173_) );
INVX1 INVX1_79 ( .A(_173_), .Y(_174_) );
NAND3X1 NAND3X1_60 ( .A(_166_), .B(_174_), .C(_171_), .Y(_175_) );
OAI21X1 OAI21X1_56 ( .A(i_add2[28]), .B(i_add1[28]), .C(_175_), .Y(_176_) );
INVX1 INVX1_80 ( .A(_176_), .Y(w_C_29_) );
INVX1 INVX1_81 ( .A(i_add2[29]), .Y(_177_) );
INVX1 INVX1_82 ( .A(i_add1[29]), .Y(_178_) );
NOR2X1 NOR2X1_62 ( .A(_177_), .B(_178_), .Y(_179_) );
INVX1 INVX1_83 ( .A(_179_), .Y(_180_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_181_) );
INVX1 INVX1_84 ( .A(_181_), .Y(_182_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_183_) );
INVX1 INVX1_85 ( .A(_183_), .Y(_184_) );
NAND3X1 NAND3X1_61 ( .A(_182_), .B(_184_), .C(_175_), .Y(_185_) );
AND2X2 AND2X2_61 ( .A(_185_), .B(_180_), .Y(_186_) );
INVX1 INVX1_86 ( .A(_186_), .Y(w_C_30_) );
AND2X2 AND2X2_62 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_187_) );
INVX1 INVX1_87 ( .A(_187_), .Y(_188_) );
NAND3X1 NAND3X1_62 ( .A(_180_), .B(_188_), .C(_185_), .Y(_189_) );
OAI21X1 OAI21X1_57 ( .A(i_add2[30]), .B(i_add1[30]), .C(_189_), .Y(_190_) );
INVX1 INVX1_88 ( .A(_190_), .Y(w_C_31_) );
INVX1 INVX1_89 ( .A(i_add2[31]), .Y(_191_) );
INVX1 INVX1_90 ( .A(i_add1[31]), .Y(_192_) );
NOR2X1 NOR2X1_65 ( .A(_191_), .B(_192_), .Y(_193_) );
INVX1 INVX1_91 ( .A(_193_), .Y(_194_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_195_) );
INVX1 INVX1_92 ( .A(_195_), .Y(_196_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_197_) );
INVX1 INVX1_93 ( .A(_197_), .Y(_198_) );
NAND3X1 NAND3X1_63 ( .A(_196_), .B(_198_), .C(_189_), .Y(_199_) );
AND2X2 AND2X2_63 ( .A(_199_), .B(_194_), .Y(_200_) );
INVX1 INVX1_94 ( .A(_200_), .Y(w_C_32_) );
AND2X2 AND2X2_64 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_201_) );
INVX1 INVX1_95 ( .A(_201_), .Y(_202_) );
NAND3X1 NAND3X1_64 ( .A(_194_), .B(_202_), .C(_199_), .Y(_203_) );
OAI21X1 OAI21X1_58 ( .A(i_add2[32]), .B(i_add1[32]), .C(_203_), .Y(_204_) );
INVX1 INVX1_96 ( .A(_204_), .Y(w_C_33_) );
INVX1 INVX1_97 ( .A(i_add2[33]), .Y(_205_) );
INVX1 INVX1_98 ( .A(i_add1[33]), .Y(_206_) );
NOR2X1 NOR2X1_68 ( .A(_205_), .B(_206_), .Y(_207_) );
INVX1 INVX1_99 ( .A(_207_), .Y(_208_) );
NOR2X1 NOR2X1_69 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_209_) );
INVX1 INVX1_100 ( .A(_209_), .Y(_210_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_211_) );
INVX1 INVX1_101 ( .A(_211_), .Y(_212_) );
NAND3X1 NAND3X1_65 ( .A(_210_), .B(_212_), .C(_203_), .Y(_213_) );
AND2X2 AND2X2_65 ( .A(_213_), .B(_208_), .Y(_214_) );
INVX1 INVX1_102 ( .A(_214_), .Y(w_C_34_) );
AND2X2 AND2X2_66 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_215_) );
INVX1 INVX1_103 ( .A(_215_), .Y(_216_) );
NAND3X1 NAND3X1_66 ( .A(_208_), .B(_216_), .C(_213_), .Y(_217_) );
OAI21X1 OAI21X1_59 ( .A(i_add2[34]), .B(i_add1[34]), .C(_217_), .Y(_218_) );
INVX1 INVX1_104 ( .A(_218_), .Y(w_C_35_) );
INVX1 INVX1_105 ( .A(i_add2[35]), .Y(_219_) );
INVX1 INVX1_106 ( .A(i_add1[35]), .Y(_220_) );
NOR2X1 NOR2X1_71 ( .A(_219_), .B(_220_), .Y(_221_) );
INVX1 INVX1_107 ( .A(_221_), .Y(_222_) );
NOR2X1 NOR2X1_72 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_223_) );
INVX1 INVX1_108 ( .A(_223_), .Y(_224_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_225_) );
INVX1 INVX1_109 ( .A(_225_), .Y(_226_) );
NAND3X1 NAND3X1_67 ( .A(_224_), .B(_226_), .C(_217_), .Y(_227_) );
AND2X2 AND2X2_67 ( .A(_227_), .B(_222_), .Y(_228_) );
INVX1 INVX1_110 ( .A(_228_), .Y(w_C_36_) );
AND2X2 AND2X2_68 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_229_) );
INVX1 INVX1_111 ( .A(_229_), .Y(_230_) );
NAND3X1 NAND3X1_68 ( .A(_222_), .B(_230_), .C(_227_), .Y(_231_) );
OAI21X1 OAI21X1_60 ( .A(i_add2[36]), .B(i_add1[36]), .C(_231_), .Y(_232_) );
INVX1 INVX1_112 ( .A(_232_), .Y(w_C_37_) );
INVX1 INVX1_113 ( .A(i_add2[37]), .Y(_233_) );
INVX1 INVX1_114 ( .A(i_add1[37]), .Y(_234_) );
NOR2X1 NOR2X1_74 ( .A(_233_), .B(_234_), .Y(_235_) );
INVX1 INVX1_115 ( .A(_235_), .Y(_236_) );
NOR2X1 NOR2X1_75 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_237_) );
INVX1 INVX1_116 ( .A(_237_), .Y(_238_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_239_) );
INVX1 INVX1_117 ( .A(_239_), .Y(_240_) );
NAND3X1 NAND3X1_69 ( .A(_238_), .B(_240_), .C(_231_), .Y(_241_) );
AND2X2 AND2X2_69 ( .A(_241_), .B(_236_), .Y(_242_) );
INVX1 INVX1_118 ( .A(_242_), .Y(w_C_38_) );
AND2X2 AND2X2_70 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_243_) );
INVX1 INVX1_119 ( .A(_243_), .Y(_244_) );
NAND3X1 NAND3X1_70 ( .A(_236_), .B(_244_), .C(_241_), .Y(_245_) );
OAI21X1 OAI21X1_61 ( .A(i_add2[38]), .B(i_add1[38]), .C(_245_), .Y(_246_) );
INVX1 INVX1_120 ( .A(_246_), .Y(w_C_39_) );
INVX1 INVX1_121 ( .A(i_add2[39]), .Y(_247_) );
INVX1 INVX1_122 ( .A(i_add1[39]), .Y(_248_) );
NOR2X1 NOR2X1_77 ( .A(_247_), .B(_248_), .Y(_249_) );
INVX1 INVX1_123 ( .A(_249_), .Y(_250_) );
NOR2X1 NOR2X1_78 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_251_) );
INVX1 INVX1_124 ( .A(_251_), .Y(_252_) );
NOR2X1 NOR2X1_79 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_253_) );
INVX1 INVX1_125 ( .A(_253_), .Y(_254_) );
NAND3X1 NAND3X1_71 ( .A(_252_), .B(_254_), .C(_245_), .Y(_255_) );
AND2X2 AND2X2_71 ( .A(_255_), .B(_250_), .Y(_256_) );
INVX1 INVX1_126 ( .A(_256_), .Y(w_C_40_) );
AND2X2 AND2X2_72 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_257_) );
INVX1 INVX1_127 ( .A(_257_), .Y(_258_) );
NAND3X1 NAND3X1_72 ( .A(_250_), .B(_258_), .C(_255_), .Y(_259_) );
OAI21X1 OAI21X1_62 ( .A(i_add2[40]), .B(i_add1[40]), .C(_259_), .Y(_260_) );
INVX1 INVX1_128 ( .A(_260_), .Y(w_C_41_) );
NAND2X1 NAND2X1_105 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_261_) );
NOR2X1 NOR2X1_80 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_262_) );
OAI21X1 OAI21X1_63 ( .A(_262_), .B(_260_), .C(_261_), .Y(w_C_42_) );
OR2X2 OR2X2_53 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_263_) );
NOR2X1 NOR2X1_81 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_264_) );
INVX1 INVX1_129 ( .A(_264_), .Y(_265_) );
INVX1 INVX1_130 ( .A(_262_), .Y(_266_) );
NAND3X1 NAND3X1_73 ( .A(_265_), .B(_266_), .C(_259_), .Y(_267_) );
NAND2X1 NAND2X1_106 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_268_) );
NAND3X1 NAND3X1_74 ( .A(_261_), .B(_268_), .C(_267_), .Y(_269_) );
AND2X2 AND2X2_73 ( .A(_269_), .B(_263_), .Y(w_C_43_) );
INVX1 INVX1_131 ( .A(i_add2[43]), .Y(_270_) );
INVX1 INVX1_132 ( .A(i_add1[43]), .Y(_271_) );
NAND2X1 NAND2X1_107 ( .A(_270_), .B(_271_), .Y(_272_) );
NAND3X1 NAND3X1_75 ( .A(_263_), .B(_272_), .C(_269_), .Y(_273_) );
OAI21X1 OAI21X1_64 ( .A(_270_), .B(_271_), .C(_273_), .Y(w_C_44_) );
INVX1 INVX1_133 ( .A(i_add2[44]), .Y(_274_) );
INVX1 INVX1_134 ( .A(i_add1[44]), .Y(_275_) );
NAND2X1 NAND2X1_108 ( .A(_274_), .B(_275_), .Y(_276_) );
NAND2X1 NAND2X1_109 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_277_) );
NAND2X1 NAND2X1_110 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_278_) );
NAND3X1 NAND3X1_76 ( .A(_277_), .B(_278_), .C(_273_), .Y(_279_) );
AND2X2 AND2X2_74 ( .A(_279_), .B(_276_), .Y(w_C_45_) );
INVX1 INVX1_135 ( .A(i_add2[45]), .Y(_280_) );
INVX1 INVX1_136 ( .A(i_add1[45]), .Y(_281_) );
NAND2X1 NAND2X1_111 ( .A(_280_), .B(_281_), .Y(_282_) );
NAND3X1 NAND3X1_77 ( .A(_276_), .B(_282_), .C(_279_), .Y(_283_) );
OAI21X1 OAI21X1_65 ( .A(_280_), .B(_281_), .C(_283_), .Y(w_C_46_) );
INVX1 INVX1_137 ( .A(i_add2[46]), .Y(_284_) );
INVX1 INVX1_138 ( .A(i_add1[46]), .Y(_285_) );
OAI21X1 OAI21X1_66 ( .A(i_add2[46]), .B(i_add1[46]), .C(w_C_46_), .Y(_286_) );
OAI21X1 OAI21X1_67 ( .A(_284_), .B(_285_), .C(_286_), .Y(w_C_47_) );
NOR2X1 NOR2X1_82 ( .A(_284_), .B(_285_), .Y(_287_) );
INVX1 INVX1_139 ( .A(_287_), .Y(_288_) );
AND2X2 AND2X2_75 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_289_) );
INVX1 INVX1_140 ( .A(_289_), .Y(_290_) );
NAND3X1 NAND3X1_78 ( .A(_288_), .B(_290_), .C(_286_), .Y(_291_) );
OAI21X1 OAI21X1_68 ( .A(i_add2[47]), .B(i_add1[47]), .C(_291_), .Y(_292_) );
INVX1 INVX1_141 ( .A(_292_), .Y(w_C_48_) );
NAND2X1 NAND2X1_112 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_293_) );
NOR2X1 NOR2X1_83 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_294_) );
OAI21X1 OAI21X1_69 ( .A(_294_), .B(_292_), .C(_293_), .Y(w_C_49_) );
NAND2X1 NAND2X1_113 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_295_) );
INVX1 INVX1_142 ( .A(_294_), .Y(_296_) );
NOR2X1 NOR2X1_84 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_297_) );
INVX1 INVX1_143 ( .A(_297_), .Y(_298_) );
NOR2X1 NOR2X1_85 ( .A(_280_), .B(_281_), .Y(_299_) );
INVX1 INVX1_144 ( .A(_299_), .Y(_300_) );
NAND3X1 NAND3X1_79 ( .A(_300_), .B(_288_), .C(_283_), .Y(_301_) );
NOR2X1 NOR2X1_86 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_302_) );
INVX1 INVX1_145 ( .A(_302_), .Y(_303_) );
NAND3X1 NAND3X1_80 ( .A(_298_), .B(_303_), .C(_301_), .Y(_304_) );
NAND3X1 NAND3X1_81 ( .A(_290_), .B(_293_), .C(_304_), .Y(_305_) );
OR2X2 OR2X2_54 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_306_) );
NAND3X1 NAND3X1_82 ( .A(_296_), .B(_306_), .C(_305_), .Y(_307_) );
NAND2X1 NAND2X1_114 ( .A(_295_), .B(_307_), .Y(w_C_50_) );
OR2X2 OR2X2_55 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_308_) );
NAND2X1 NAND2X1_115 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_309_) );
NAND3X1 NAND3X1_83 ( .A(_295_), .B(_309_), .C(_307_), .Y(_310_) );
AND2X2 AND2X2_76 ( .A(_310_), .B(_308_), .Y(w_C_51_) );
NAND2X1 NAND2X1_116 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_311_) );
OR2X2 OR2X2_56 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_312_) );
NAND3X1 NAND3X1_84 ( .A(_308_), .B(_312_), .C(_310_), .Y(_313_) );
NAND2X1 NAND2X1_117 ( .A(_311_), .B(_313_), .Y(w_C_52_) );
NAND2X1 NAND2X1_118 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_146 ( .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_87 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_88 ( .A(_1_), .B(_2_), .Y(w_C_2_) );
NAND2X1 NAND2X1_119 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_3_) );
OAI21X1 OAI21X1_70 ( .A(_1_), .B(_2_), .C(_3_), .Y(_4_) );
OAI21X1 OAI21X1_71 ( .A(i_add2[2]), .B(i_add1[2]), .C(_4_), .Y(_5_) );
INVX1 INVX1_147 ( .A(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_120 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_6_) );
OR2X2 OR2X2_57 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_7_) );
OR2X2 OR2X2_58 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
NAND3X1 NAND3X1_85 ( .A(_7_), .B(_8_), .C(_4_), .Y(_9_) );
NAND2X1 NAND2X1_121 ( .A(_6_), .B(_9_), .Y(w_C_4_) );
NAND2X1 NAND2X1_122 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_10_) );
NAND3X1 NAND3X1_86 ( .A(_6_), .B(_10_), .C(_9_), .Y(_11_) );
OAI21X1 OAI21X1_72 ( .A(i_add2[4]), .B(i_add1[4]), .C(_11_), .Y(_12_) );
INVX1 INVX1_148 ( .A(_12_), .Y(w_C_5_) );
INVX1 INVX1_149 ( .A(i_add2[5]), .Y(_13_) );
INVX1 INVX1_150 ( .A(i_add1[5]), .Y(_14_) );
NOR2X1 NOR2X1_89 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_15_) );
INVX1 INVX1_151 ( .A(_15_), .Y(_16_) );
NOR2X1 NOR2X1_90 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_17_) );
INVX1 INVX1_152 ( .A(_17_), .Y(_18_) );
NAND3X1 NAND3X1_87 ( .A(_16_), .B(_18_), .C(_11_), .Y(_19_) );
OAI21X1 OAI21X1_73 ( .A(_13_), .B(_14_), .C(_19_), .Y(w_C_6_) );
NOR2X1 NOR2X1_91 ( .A(_13_), .B(_14_), .Y(_20_) );
INVX1 INVX1_153 ( .A(_20_), .Y(_21_) );
AND2X2 AND2X2_77 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_154 ( .A(_22_), .Y(_23_) );
NAND3X1 NAND3X1_88 ( .A(_21_), .B(_23_), .C(_19_), .Y(_24_) );
OAI21X1 OAI21X1_74 ( .A(i_add2[6]), .B(i_add1[6]), .C(_24_), .Y(_25_) );
INVX1 INVX1_155 ( .A(_25_), .Y(w_C_7_) );
INVX1 INVX1_156 ( .A(i_add2[7]), .Y(_26_) );
INVX1 INVX1_157 ( .A(i_add1[7]), .Y(_27_) );
NOR2X1 NOR2X1_92 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_28_) );
INVX1 INVX1_158 ( .A(_28_), .Y(_29_) );
NOR2X1 NOR2X1_93 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_30_) );
INVX1 INVX1_159 ( .A(_30_), .Y(_31_) );
NAND3X1 NAND3X1_89 ( .A(_29_), .B(_31_), .C(_24_), .Y(_32_) );
OAI21X1 OAI21X1_75 ( .A(_26_), .B(_27_), .C(_32_), .Y(w_C_8_) );
NOR2X1 NOR2X1_94 ( .A(_26_), .B(_27_), .Y(_33_) );
INVX1 INVX1_160 ( .A(_33_), .Y(_34_) );
AND2X2 AND2X2_78 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_35_) );
INVX1 INVX1_161 ( .A(_35_), .Y(_36_) );
NAND3X1 NAND3X1_90 ( .A(_34_), .B(_36_), .C(_32_), .Y(_37_) );
OAI21X1 OAI21X1_76 ( .A(i_add2[8]), .B(i_add1[8]), .C(_37_), .Y(_38_) );
INVX1 INVX1_162 ( .A(_38_), .Y(w_C_9_) );
INVX1 INVX1_163 ( .A(i_add2[9]), .Y(_39_) );
INVX1 INVX1_164 ( .A(i_add1[9]), .Y(_40_) );
NOR2X1 NOR2X1_95 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_41_) );
INVX1 INVX1_165 ( .A(_41_), .Y(_42_) );
NOR2X1 NOR2X1_96 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_43_) );
INVX1 INVX1_166 ( .A(_43_), .Y(_44_) );
NAND3X1 NAND3X1_91 ( .A(_42_), .B(_44_), .C(_37_), .Y(_45_) );
OAI21X1 OAI21X1_77 ( .A(_39_), .B(_40_), .C(_45_), .Y(w_C_10_) );
NOR2X1 NOR2X1_97 ( .A(_39_), .B(_40_), .Y(_46_) );
INVX1 INVX1_167 ( .A(_46_), .Y(_47_) );
AND2X2 AND2X2_79 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_48_) );
INVX1 INVX1_168 ( .A(_48_), .Y(_49_) );
NAND3X1 NAND3X1_92 ( .A(_47_), .B(_49_), .C(_45_), .Y(_50_) );
OAI21X1 OAI21X1_78 ( .A(i_add2[10]), .B(i_add1[10]), .C(_50_), .Y(_51_) );
INVX1 INVX1_169 ( .A(_51_), .Y(w_C_11_) );
INVX1 INVX1_170 ( .A(i_add2[11]), .Y(_52_) );
INVX1 INVX1_171 ( .A(i_add1[11]), .Y(_53_) );
NOR2X1 NOR2X1_98 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_54_) );
INVX1 INVX1_172 ( .A(_54_), .Y(_55_) );
NOR2X1 NOR2X1_99 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_56_) );
INVX1 INVX1_173 ( .A(_56_), .Y(_57_) );
NAND3X1 NAND3X1_93 ( .A(_55_), .B(_57_), .C(_50_), .Y(_58_) );
OAI21X1 OAI21X1_79 ( .A(_52_), .B(_53_), .C(_58_), .Y(w_C_12_) );
NOR2X1 NOR2X1_100 ( .A(_52_), .B(_53_), .Y(_59_) );
INVX1 INVX1_174 ( .A(_59_), .Y(_60_) );
AND2X2 AND2X2_80 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_61_) );
INVX1 INVX1_175 ( .A(_61_), .Y(_62_) );
NAND3X1 NAND3X1_94 ( .A(_60_), .B(_62_), .C(_58_), .Y(_63_) );
OAI21X1 OAI21X1_80 ( .A(i_add2[12]), .B(i_add1[12]), .C(_63_), .Y(_64_) );
INVX1 INVX1_176 ( .A(_64_), .Y(w_C_13_) );
INVX1 INVX1_177 ( .A(i_add2[13]), .Y(_65_) );
INVX1 INVX1_178 ( .A(i_add1[13]), .Y(_66_) );
NOR2X1 NOR2X1_101 ( .A(_65_), .B(_66_), .Y(_67_) );
INVX1 INVX1_179 ( .A(_67_), .Y(_68_) );
NOR2X1 NOR2X1_102 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_69_) );
INVX1 INVX1_180 ( .A(_69_), .Y(_70_) );
NOR2X1 NOR2X1_103 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_71_) );
INVX1 INVX1_181 ( .A(_71_), .Y(_72_) );
NAND3X1 NAND3X1_95 ( .A(_70_), .B(_72_), .C(_63_), .Y(_73_) );
AND2X2 AND2X2_81 ( .A(_73_), .B(_68_), .Y(_74_) );
INVX1 INVX1_182 ( .A(_74_), .Y(w_C_14_) );
AND2X2 AND2X2_82 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_75_) );
INVX1 INVX1_183 ( .A(_75_), .Y(_76_) );
NAND3X1 NAND3X1_96 ( .A(_68_), .B(_76_), .C(_73_), .Y(_77_) );
OAI21X1 OAI21X1_81 ( .A(i_add2[14]), .B(i_add1[14]), .C(_77_), .Y(_78_) );
INVX1 INVX1_184 ( .A(_78_), .Y(w_C_15_) );
INVX1 INVX1_185 ( .A(i_add2[15]), .Y(_79_) );
INVX1 INVX1_186 ( .A(i_add1[15]), .Y(_80_) );
NOR2X1 NOR2X1_104 ( .A(_79_), .B(_80_), .Y(_81_) );
INVX1 INVX1_187 ( .A(_81_), .Y(_82_) );
NOR2X1 NOR2X1_105 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_83_) );
INVX1 INVX1_188 ( .A(_83_), .Y(_84_) );
NOR2X1 NOR2X1_106 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_85_) );
INVX1 INVX1_189 ( .A(_85_), .Y(_86_) );
NAND3X1 NAND3X1_97 ( .A(_84_), .B(_86_), .C(_77_), .Y(_87_) );
AND2X2 AND2X2_83 ( .A(_87_), .B(_82_), .Y(_88_) );
INVX1 INVX1_190 ( .A(_88_), .Y(w_C_16_) );
AND2X2 AND2X2_84 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_89_) );
INVX1 INVX1_191 ( .A(_89_), .Y(_90_) );
NAND3X1 NAND3X1_98 ( .A(_82_), .B(_90_), .C(_87_), .Y(_91_) );
OAI21X1 OAI21X1_82 ( .A(i_add2[16]), .B(i_add1[16]), .C(_91_), .Y(_92_) );
INVX1 INVX1_192 ( .A(_92_), .Y(w_C_17_) );
INVX1 INVX1_193 ( .A(i_add2[17]), .Y(_93_) );
INVX1 INVX1_194 ( .A(i_add1[17]), .Y(_94_) );
NOR2X1 NOR2X1_107 ( .A(_93_), .B(_94_), .Y(_95_) );
INVX1 INVX1_195 ( .A(_95_), .Y(_96_) );
NOR2X1 NOR2X1_108 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_97_) );
INVX1 INVX1_196 ( .A(_97_), .Y(_98_) );
NOR2X1 NOR2X1_109 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_99_) );
INVX1 INVX1_197 ( .A(_99_), .Y(_100_) );
NAND3X1 NAND3X1_99 ( .A(_98_), .B(_100_), .C(_91_), .Y(_101_) );
AND2X2 AND2X2_85 ( .A(_101_), .B(_96_), .Y(_102_) );
INVX1 INVX1_198 ( .A(_102_), .Y(w_C_18_) );
AND2X2 AND2X2_86 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_103_) );
INVX1 INVX1_199 ( .A(_103_), .Y(_104_) );
NAND3X1 NAND3X1_100 ( .A(_96_), .B(_104_), .C(_101_), .Y(_105_) );
OAI21X1 OAI21X1_83 ( .A(i_add2[18]), .B(i_add1[18]), .C(_105_), .Y(_106_) );
INVX1 INVX1_200 ( .A(_106_), .Y(w_C_19_) );
INVX1 INVX1_201 ( .A(i_add2[19]), .Y(_107_) );
INVX1 INVX1_202 ( .A(i_add1[19]), .Y(_108_) );
NOR2X1 NOR2X1_110 ( .A(_107_), .B(_108_), .Y(_109_) );
INVX1 INVX1_203 ( .A(_109_), .Y(_110_) );
NOR2X1 NOR2X1_111 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_111_) );
INVX1 INVX1_204 ( .A(_111_), .Y(_112_) );
NOR2X1 NOR2X1_112 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_113_) );
INVX1 INVX1_205 ( .A(_113_), .Y(_114_) );
NAND3X1 NAND3X1_101 ( .A(_112_), .B(_114_), .C(_105_), .Y(_115_) );
AND2X2 AND2X2_87 ( .A(_115_), .B(_110_), .Y(_116_) );
INVX1 INVX1_206 ( .A(_116_), .Y(w_C_20_) );
AND2X2 AND2X2_88 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_117_) );
INVX1 INVX1_207 ( .A(_117_), .Y(_118_) );
NAND3X1 NAND3X1_102 ( .A(_110_), .B(_118_), .C(_115_), .Y(_119_) );
OAI21X1 OAI21X1_84 ( .A(i_add2[20]), .B(i_add1[20]), .C(_119_), .Y(_120_) );
INVX1 INVX1_208 ( .A(_120_), .Y(w_C_21_) );
INVX1 INVX1_209 ( .A(i_add2[21]), .Y(_121_) );
INVX1 INVX1_210 ( .A(i_add1[21]), .Y(_122_) );
NOR2X1 NOR2X1_113 ( .A(_121_), .B(_122_), .Y(_123_) );
INVX1 INVX1_211 ( .A(_123_), .Y(_124_) );
NOR2X1 NOR2X1_114 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_125_) );
INVX1 INVX1_212 ( .A(_125_), .Y(_126_) );
NOR2X1 NOR2X1_115 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_127_) );
BUFX2 BUFX2_54 ( .A(w_C_52_), .Y(_314__52_) );
BUFX2 BUFX2_55 ( .A(1'b0), .Y(w_C_0_) );
endmodule
