module csa_30bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output cout;

NAND3X1 NAND3X1_1 ( .A(_382_), .B(_384_), .C(_383_), .Y(_385_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_379_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_380_) );
OAI21X1 OAI21X1_1 ( .A(_379_), .B(_380_), .C(_30__2_), .Y(_381_) );
NAND2X1 NAND2X1_1 ( .A(_381_), .B(_385_), .Y(_28__2_) );
OAI21X1 OAI21X1_2 ( .A(_382_), .B(_379_), .C(_384_), .Y(_30__3_) );
INVX1 INVX1_1 ( .A(_30__3_), .Y(_389_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_390_) );
NAND2X1 NAND2X1_2 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_391_) );
NAND3X1 NAND3X1_2 ( .A(_389_), .B(_391_), .C(_390_), .Y(_392_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_386_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_387_) );
OAI21X1 OAI21X1_3 ( .A(_386_), .B(_387_), .C(_30__3_), .Y(_388_) );
NAND2X1 NAND2X1_3 ( .A(_388_), .B(_392_), .Y(_28__3_) );
OAI21X1 OAI21X1_4 ( .A(_389_), .B(_386_), .C(_391_), .Y(_26_) );
INVX1 INVX1_2 ( .A(1'b0), .Y(_396_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_397_) );
NAND2X1 NAND2X1_4 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_398_) );
NAND3X1 NAND3X1_3 ( .A(_396_), .B(_398_), .C(_397_), .Y(_399_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_393_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_394_) );
OAI21X1 OAI21X1_5 ( .A(_393_), .B(_394_), .C(1'b0), .Y(_395_) );
NAND2X1 NAND2X1_5 ( .A(_395_), .B(_399_), .Y(_33__0_) );
OAI21X1 OAI21X1_6 ( .A(_396_), .B(_393_), .C(_398_), .Y(_35__1_) );
INVX1 INVX1_3 ( .A(_35__1_), .Y(_403_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_404_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_405_) );
NAND3X1 NAND3X1_4 ( .A(_403_), .B(_405_), .C(_404_), .Y(_406_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_400_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_401_) );
OAI21X1 OAI21X1_7 ( .A(_400_), .B(_401_), .C(_35__1_), .Y(_402_) );
NAND2X1 NAND2X1_7 ( .A(_402_), .B(_406_), .Y(_33__1_) );
OAI21X1 OAI21X1_8 ( .A(_403_), .B(_400_), .C(_405_), .Y(_35__2_) );
INVX1 INVX1_4 ( .A(_35__2_), .Y(_410_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_411_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_412_) );
NAND3X1 NAND3X1_5 ( .A(_410_), .B(_412_), .C(_411_), .Y(_413_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_407_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_408_) );
OAI21X1 OAI21X1_9 ( .A(_407_), .B(_408_), .C(_35__2_), .Y(_409_) );
NAND2X1 NAND2X1_9 ( .A(_409_), .B(_413_), .Y(_33__2_) );
OAI21X1 OAI21X1_10 ( .A(_410_), .B(_407_), .C(_412_), .Y(_35__3_) );
INVX1 INVX1_5 ( .A(_35__3_), .Y(_417_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_418_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_419_) );
NAND3X1 NAND3X1_6 ( .A(_417_), .B(_419_), .C(_418_), .Y(_420_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_414_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_415_) );
OAI21X1 OAI21X1_11 ( .A(_414_), .B(_415_), .C(_35__3_), .Y(_416_) );
NAND2X1 NAND2X1_11 ( .A(_416_), .B(_420_), .Y(_33__3_) );
OAI21X1 OAI21X1_12 ( .A(_417_), .B(_414_), .C(_419_), .Y(_31_) );
INVX1 INVX1_6 ( .A(1'b1), .Y(_424_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_425_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_426_) );
NAND3X1 NAND3X1_7 ( .A(_424_), .B(_426_), .C(_425_), .Y(_427_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_421_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_422_) );
OAI21X1 OAI21X1_13 ( .A(_421_), .B(_422_), .C(1'b1), .Y(_423_) );
NAND2X1 NAND2X1_13 ( .A(_423_), .B(_427_), .Y(_34__0_) );
OAI21X1 OAI21X1_14 ( .A(_424_), .B(_421_), .C(_426_), .Y(_36__1_) );
INVX1 INVX1_7 ( .A(_36__1_), .Y(_431_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_432_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_433_) );
NAND3X1 NAND3X1_8 ( .A(_431_), .B(_433_), .C(_432_), .Y(_434_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_428_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_429_) );
OAI21X1 OAI21X1_15 ( .A(_428_), .B(_429_), .C(_36__1_), .Y(_430_) );
NAND2X1 NAND2X1_15 ( .A(_430_), .B(_434_), .Y(_34__1_) );
OAI21X1 OAI21X1_16 ( .A(_431_), .B(_428_), .C(_433_), .Y(_36__2_) );
INVX1 INVX1_8 ( .A(_36__2_), .Y(_438_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_439_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_440_) );
NAND3X1 NAND3X1_9 ( .A(_438_), .B(_440_), .C(_439_), .Y(_441_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_435_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_436_) );
OAI21X1 OAI21X1_17 ( .A(_435_), .B(_436_), .C(_36__2_), .Y(_437_) );
NAND2X1 NAND2X1_17 ( .A(_437_), .B(_441_), .Y(_34__2_) );
OAI21X1 OAI21X1_18 ( .A(_438_), .B(_435_), .C(_440_), .Y(_36__3_) );
INVX1 INVX1_9 ( .A(_36__3_), .Y(_445_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_446_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_447_) );
NAND3X1 NAND3X1_10 ( .A(_445_), .B(_447_), .C(_446_), .Y(_448_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_442_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_443_) );
OAI21X1 OAI21X1_19 ( .A(_442_), .B(_443_), .C(_36__3_), .Y(_444_) );
NAND2X1 NAND2X1_19 ( .A(_444_), .B(_448_), .Y(_34__3_) );
OAI21X1 OAI21X1_20 ( .A(_445_), .B(_442_), .C(_447_), .Y(_32_) );
INVX1 INVX1_10 ( .A(1'b0), .Y(_452_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_453_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_454_) );
NAND3X1 NAND3X1_11 ( .A(_452_), .B(_454_), .C(_453_), .Y(_455_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_449_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_450_) );
OAI21X1 OAI21X1_21 ( .A(_449_), .B(_450_), .C(1'b0), .Y(_451_) );
NAND2X1 NAND2X1_21 ( .A(_451_), .B(_455_), .Y(_39__0_) );
OAI21X1 OAI21X1_22 ( .A(_452_), .B(_449_), .C(_454_), .Y(_41__1_) );
INVX1 INVX1_11 ( .A(_41__1_), .Y(_459_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_460_) );
NAND2X1 NAND2X1_22 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_461_) );
NAND3X1 NAND3X1_12 ( .A(_459_), .B(_461_), .C(_460_), .Y(_462_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_456_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_457_) );
OAI21X1 OAI21X1_23 ( .A(_456_), .B(_457_), .C(_41__1_), .Y(_458_) );
NAND2X1 NAND2X1_23 ( .A(_458_), .B(_462_), .Y(_39__1_) );
OAI21X1 OAI21X1_24 ( .A(_459_), .B(_456_), .C(_461_), .Y(_41__2_) );
INVX1 INVX1_12 ( .A(_41__2_), .Y(_466_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_467_) );
NAND2X1 NAND2X1_24 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_468_) );
NAND3X1 NAND3X1_13 ( .A(_466_), .B(_468_), .C(_467_), .Y(_469_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_463_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_464_) );
OAI21X1 OAI21X1_25 ( .A(_463_), .B(_464_), .C(_41__2_), .Y(_465_) );
NAND2X1 NAND2X1_25 ( .A(_465_), .B(_469_), .Y(_39__2_) );
OAI21X1 OAI21X1_26 ( .A(_466_), .B(_463_), .C(_468_), .Y(_41__3_) );
INVX1 INVX1_13 ( .A(_41__3_), .Y(_473_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_474_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_475_) );
NAND3X1 NAND3X1_14 ( .A(_473_), .B(_475_), .C(_474_), .Y(_476_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_470_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_471_) );
OAI21X1 OAI21X1_27 ( .A(_470_), .B(_471_), .C(_41__3_), .Y(_472_) );
NAND2X1 NAND2X1_27 ( .A(_472_), .B(_476_), .Y(_39__3_) );
OAI21X1 OAI21X1_28 ( .A(_473_), .B(_470_), .C(_475_), .Y(_37_) );
INVX1 INVX1_14 ( .A(1'b1), .Y(_480_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_481_) );
NAND2X1 NAND2X1_28 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_482_) );
NAND3X1 NAND3X1_15 ( .A(_480_), .B(_482_), .C(_481_), .Y(_483_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_477_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_478_) );
OAI21X1 OAI21X1_29 ( .A(_477_), .B(_478_), .C(1'b1), .Y(_479_) );
NAND2X1 NAND2X1_29 ( .A(_479_), .B(_483_), .Y(_40__0_) );
OAI21X1 OAI21X1_30 ( .A(_480_), .B(_477_), .C(_482_), .Y(_42__1_) );
INVX1 INVX1_15 ( .A(_42__1_), .Y(_487_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_488_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_489_) );
NAND3X1 NAND3X1_16 ( .A(_487_), .B(_489_), .C(_488_), .Y(_490_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_484_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_485_) );
OAI21X1 OAI21X1_31 ( .A(_484_), .B(_485_), .C(_42__1_), .Y(_486_) );
NAND2X1 NAND2X1_31 ( .A(_486_), .B(_490_), .Y(_40__1_) );
OAI21X1 OAI21X1_32 ( .A(_487_), .B(_484_), .C(_489_), .Y(_42__2_) );
INVX1 INVX1_16 ( .A(_42__2_), .Y(_494_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_495_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_496_) );
NAND3X1 NAND3X1_17 ( .A(_494_), .B(_496_), .C(_495_), .Y(_497_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_491_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_492_) );
OAI21X1 OAI21X1_33 ( .A(_491_), .B(_492_), .C(_42__2_), .Y(_493_) );
NAND2X1 NAND2X1_33 ( .A(_493_), .B(_497_), .Y(_40__2_) );
OAI21X1 OAI21X1_34 ( .A(_494_), .B(_491_), .C(_496_), .Y(_42__3_) );
INVX1 INVX1_17 ( .A(_42__3_), .Y(_501_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_502_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_503_) );
NAND3X1 NAND3X1_18 ( .A(_501_), .B(_503_), .C(_502_), .Y(_504_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_498_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_499_) );
OAI21X1 OAI21X1_35 ( .A(_498_), .B(_499_), .C(_42__3_), .Y(_500_) );
NAND2X1 NAND2X1_35 ( .A(_500_), .B(_504_), .Y(_40__3_) );
OAI21X1 OAI21X1_36 ( .A(_501_), .B(_498_), .C(_503_), .Y(_38_) );
INVX1 INVX1_18 ( .A(1'b0), .Y(_508_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_509_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_510_) );
NAND3X1 NAND3X1_19 ( .A(_508_), .B(_510_), .C(_509_), .Y(_511_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_505_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_506_) );
OAI21X1 OAI21X1_37 ( .A(_505_), .B(_506_), .C(1'b0), .Y(_507_) );
NAND2X1 NAND2X1_37 ( .A(_507_), .B(_511_), .Y(_0__0_) );
OAI21X1 OAI21X1_38 ( .A(_508_), .B(_505_), .C(_510_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_19 ( .A(rca_inst_w_CARRY_1_), .Y(_515_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_516_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_517_) );
NAND3X1 NAND3X1_20 ( .A(_515_), .B(_517_), .C(_516_), .Y(_518_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_512_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_513_) );
OAI21X1 OAI21X1_39 ( .A(_512_), .B(_513_), .C(rca_inst_w_CARRY_1_), .Y(_514_) );
NAND2X1 NAND2X1_39 ( .A(_514_), .B(_518_), .Y(_0__1_) );
BUFX2 BUFX2_1 ( .A(w_cout_7_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
INVX1 INVX1_20 ( .A(_1_), .Y(_43_) );
NAND2X1 NAND2X1_40 ( .A(_2_), .B(1'b0), .Y(_44_) );
OAI21X1 OAI21X1_40 ( .A(1'b0), .B(_43_), .C(_44_), .Y(w_cout_1_) );
INVX1 INVX1_21 ( .A(_3__0_), .Y(_45_) );
NAND2X1 NAND2X1_41 ( .A(_4__0_), .B(1'b0), .Y(_46_) );
OAI21X1 OAI21X1_41 ( .A(1'b0), .B(_45_), .C(_46_), .Y(_0__2_) );
INVX1 INVX1_22 ( .A(_3__1_), .Y(_47_) );
NAND2X1 NAND2X1_42 ( .A(1'b0), .B(_4__1_), .Y(_48_) );
OAI21X1 OAI21X1_42 ( .A(1'b0), .B(_47_), .C(_48_), .Y(_0__3_) );
INVX1 INVX1_23 ( .A(_3__2_), .Y(_49_) );
NAND2X1 NAND2X1_43 ( .A(1'b0), .B(_4__2_), .Y(_50_) );
OAI21X1 OAI21X1_43 ( .A(1'b0), .B(_49_), .C(_50_), .Y(_0__4_) );
INVX1 INVX1_24 ( .A(_3__3_), .Y(_51_) );
NAND2X1 NAND2X1_44 ( .A(1'b0), .B(_4__3_), .Y(_52_) );
OAI21X1 OAI21X1_44 ( .A(1'b0), .B(_51_), .C(_52_), .Y(_0__5_) );
INVX1 INVX1_25 ( .A(_7_), .Y(_53_) );
NAND2X1 NAND2X1_45 ( .A(_8_), .B(w_cout_1_), .Y(_54_) );
OAI21X1 OAI21X1_45 ( .A(w_cout_1_), .B(_53_), .C(_54_), .Y(w_cout_2_) );
INVX1 INVX1_26 ( .A(_9__0_), .Y(_55_) );
NAND2X1 NAND2X1_46 ( .A(_10__0_), .B(w_cout_1_), .Y(_56_) );
OAI21X1 OAI21X1_46 ( .A(w_cout_1_), .B(_55_), .C(_56_), .Y(_0__6_) );
INVX1 INVX1_27 ( .A(_9__1_), .Y(_57_) );
NAND2X1 NAND2X1_47 ( .A(w_cout_1_), .B(_10__1_), .Y(_58_) );
OAI21X1 OAI21X1_47 ( .A(w_cout_1_), .B(_57_), .C(_58_), .Y(_0__7_) );
INVX1 INVX1_28 ( .A(_9__2_), .Y(_59_) );
NAND2X1 NAND2X1_48 ( .A(w_cout_1_), .B(_10__2_), .Y(_60_) );
OAI21X1 OAI21X1_48 ( .A(w_cout_1_), .B(_59_), .C(_60_), .Y(_0__8_) );
INVX1 INVX1_29 ( .A(_9__3_), .Y(_61_) );
NAND2X1 NAND2X1_49 ( .A(w_cout_1_), .B(_10__3_), .Y(_62_) );
OAI21X1 OAI21X1_49 ( .A(w_cout_1_), .B(_61_), .C(_62_), .Y(_0__9_) );
INVX1 INVX1_30 ( .A(_13_), .Y(_63_) );
NAND2X1 NAND2X1_50 ( .A(_14_), .B(w_cout_2_), .Y(_64_) );
OAI21X1 OAI21X1_50 ( .A(w_cout_2_), .B(_63_), .C(_64_), .Y(w_cout_3_) );
INVX1 INVX1_31 ( .A(_15__0_), .Y(_65_) );
NAND2X1 NAND2X1_51 ( .A(_16__0_), .B(w_cout_2_), .Y(_66_) );
OAI21X1 OAI21X1_51 ( .A(w_cout_2_), .B(_65_), .C(_66_), .Y(_0__10_) );
INVX1 INVX1_32 ( .A(_15__1_), .Y(_67_) );
NAND2X1 NAND2X1_52 ( .A(w_cout_2_), .B(_16__1_), .Y(_68_) );
OAI21X1 OAI21X1_52 ( .A(w_cout_2_), .B(_67_), .C(_68_), .Y(_0__11_) );
INVX1 INVX1_33 ( .A(_15__2_), .Y(_69_) );
NAND2X1 NAND2X1_53 ( .A(w_cout_2_), .B(_16__2_), .Y(_70_) );
OAI21X1 OAI21X1_53 ( .A(w_cout_2_), .B(_69_), .C(_70_), .Y(_0__12_) );
INVX1 INVX1_34 ( .A(_15__3_), .Y(_71_) );
NAND2X1 NAND2X1_54 ( .A(w_cout_2_), .B(_16__3_), .Y(_72_) );
OAI21X1 OAI21X1_54 ( .A(w_cout_2_), .B(_71_), .C(_72_), .Y(_0__13_) );
INVX1 INVX1_35 ( .A(_19_), .Y(_73_) );
NAND2X1 NAND2X1_55 ( .A(_20_), .B(w_cout_3_), .Y(_74_) );
OAI21X1 OAI21X1_55 ( .A(w_cout_3_), .B(_73_), .C(_74_), .Y(w_cout_4_) );
INVX1 INVX1_36 ( .A(_21__0_), .Y(_75_) );
NAND2X1 NAND2X1_56 ( .A(_22__0_), .B(w_cout_3_), .Y(_76_) );
OAI21X1 OAI21X1_56 ( .A(w_cout_3_), .B(_75_), .C(_76_), .Y(_0__14_) );
INVX1 INVX1_37 ( .A(_21__1_), .Y(_77_) );
NAND2X1 NAND2X1_57 ( .A(w_cout_3_), .B(_22__1_), .Y(_78_) );
OAI21X1 OAI21X1_57 ( .A(w_cout_3_), .B(_77_), .C(_78_), .Y(_0__15_) );
INVX1 INVX1_38 ( .A(_21__2_), .Y(_79_) );
NAND2X1 NAND2X1_58 ( .A(w_cout_3_), .B(_22__2_), .Y(_80_) );
OAI21X1 OAI21X1_58 ( .A(w_cout_3_), .B(_79_), .C(_80_), .Y(_0__16_) );
INVX1 INVX1_39 ( .A(_21__3_), .Y(_81_) );
NAND2X1 NAND2X1_59 ( .A(w_cout_3_), .B(_22__3_), .Y(_82_) );
OAI21X1 OAI21X1_59 ( .A(w_cout_3_), .B(_81_), .C(_82_), .Y(_0__17_) );
INVX1 INVX1_40 ( .A(_25_), .Y(_83_) );
NAND2X1 NAND2X1_60 ( .A(_26_), .B(w_cout_4_), .Y(_84_) );
OAI21X1 OAI21X1_60 ( .A(w_cout_4_), .B(_83_), .C(_84_), .Y(w_cout_5_) );
INVX1 INVX1_41 ( .A(_27__0_), .Y(_85_) );
NAND2X1 NAND2X1_61 ( .A(_28__0_), .B(w_cout_4_), .Y(_86_) );
OAI21X1 OAI21X1_61 ( .A(w_cout_4_), .B(_85_), .C(_86_), .Y(_0__18_) );
INVX1 INVX1_42 ( .A(_27__1_), .Y(_87_) );
NAND2X1 NAND2X1_62 ( .A(w_cout_4_), .B(_28__1_), .Y(_88_) );
OAI21X1 OAI21X1_62 ( .A(w_cout_4_), .B(_87_), .C(_88_), .Y(_0__19_) );
INVX1 INVX1_43 ( .A(_27__2_), .Y(_89_) );
NAND2X1 NAND2X1_63 ( .A(w_cout_4_), .B(_28__2_), .Y(_90_) );
OAI21X1 OAI21X1_63 ( .A(w_cout_4_), .B(_89_), .C(_90_), .Y(_0__20_) );
INVX1 INVX1_44 ( .A(_27__3_), .Y(_91_) );
NAND2X1 NAND2X1_64 ( .A(w_cout_4_), .B(_28__3_), .Y(_92_) );
OAI21X1 OAI21X1_64 ( .A(w_cout_4_), .B(_91_), .C(_92_), .Y(_0__21_) );
INVX1 INVX1_45 ( .A(_31_), .Y(_93_) );
NAND2X1 NAND2X1_65 ( .A(_32_), .B(w_cout_5_), .Y(_94_) );
OAI21X1 OAI21X1_65 ( .A(w_cout_5_), .B(_93_), .C(_94_), .Y(w_cout_6_) );
INVX1 INVX1_46 ( .A(_33__0_), .Y(_95_) );
NAND2X1 NAND2X1_66 ( .A(_34__0_), .B(w_cout_5_), .Y(_96_) );
OAI21X1 OAI21X1_66 ( .A(w_cout_5_), .B(_95_), .C(_96_), .Y(_0__22_) );
INVX1 INVX1_47 ( .A(_33__1_), .Y(_97_) );
NAND2X1 NAND2X1_67 ( .A(w_cout_5_), .B(_34__1_), .Y(_98_) );
OAI21X1 OAI21X1_67 ( .A(w_cout_5_), .B(_97_), .C(_98_), .Y(_0__23_) );
INVX1 INVX1_48 ( .A(_33__2_), .Y(_99_) );
NAND2X1 NAND2X1_68 ( .A(w_cout_5_), .B(_34__2_), .Y(_100_) );
OAI21X1 OAI21X1_68 ( .A(w_cout_5_), .B(_99_), .C(_100_), .Y(_0__24_) );
INVX1 INVX1_49 ( .A(_33__3_), .Y(_101_) );
NAND2X1 NAND2X1_69 ( .A(w_cout_5_), .B(_34__3_), .Y(_102_) );
OAI21X1 OAI21X1_69 ( .A(w_cout_5_), .B(_101_), .C(_102_), .Y(_0__25_) );
INVX1 INVX1_50 ( .A(_37_), .Y(_103_) );
NAND2X1 NAND2X1_70 ( .A(_38_), .B(w_cout_6_), .Y(_104_) );
OAI21X1 OAI21X1_70 ( .A(w_cout_6_), .B(_103_), .C(_104_), .Y(w_cout_7_) );
INVX1 INVX1_51 ( .A(_39__0_), .Y(_105_) );
NAND2X1 NAND2X1_71 ( .A(_40__0_), .B(w_cout_6_), .Y(_106_) );
OAI21X1 OAI21X1_71 ( .A(w_cout_6_), .B(_105_), .C(_106_), .Y(_0__26_) );
INVX1 INVX1_52 ( .A(_39__1_), .Y(_107_) );
NAND2X1 NAND2X1_72 ( .A(w_cout_6_), .B(_40__1_), .Y(_108_) );
OAI21X1 OAI21X1_72 ( .A(w_cout_6_), .B(_107_), .C(_108_), .Y(_0__27_) );
INVX1 INVX1_53 ( .A(_39__2_), .Y(_109_) );
NAND2X1 NAND2X1_73 ( .A(w_cout_6_), .B(_40__2_), .Y(_110_) );
OAI21X1 OAI21X1_73 ( .A(w_cout_6_), .B(_109_), .C(_110_), .Y(_0__28_) );
INVX1 INVX1_54 ( .A(_39__3_), .Y(_111_) );
NAND2X1 NAND2X1_74 ( .A(w_cout_6_), .B(_40__3_), .Y(_112_) );
OAI21X1 OAI21X1_74 ( .A(w_cout_6_), .B(_111_), .C(_112_), .Y(_0__29_) );
INVX1 INVX1_55 ( .A(1'b0), .Y(_116_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_117_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_118_) );
NAND3X1 NAND3X1_21 ( .A(_116_), .B(_118_), .C(_117_), .Y(_119_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_113_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_114_) );
OAI21X1 OAI21X1_75 ( .A(_113_), .B(_114_), .C(1'b0), .Y(_115_) );
NAND2X1 NAND2X1_76 ( .A(_115_), .B(_119_), .Y(_3__0_) );
OAI21X1 OAI21X1_76 ( .A(_116_), .B(_113_), .C(_118_), .Y(_5__1_) );
INVX1 INVX1_56 ( .A(_5__1_), .Y(_123_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_124_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_125_) );
NAND3X1 NAND3X1_22 ( .A(_123_), .B(_125_), .C(_124_), .Y(_126_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_120_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_121_) );
OAI21X1 OAI21X1_77 ( .A(_120_), .B(_121_), .C(_5__1_), .Y(_122_) );
NAND2X1 NAND2X1_78 ( .A(_122_), .B(_126_), .Y(_3__1_) );
OAI21X1 OAI21X1_78 ( .A(_123_), .B(_120_), .C(_125_), .Y(_5__2_) );
INVX1 INVX1_57 ( .A(_5__2_), .Y(_130_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_131_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_132_) );
NAND3X1 NAND3X1_23 ( .A(_130_), .B(_132_), .C(_131_), .Y(_133_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_127_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_128_) );
OAI21X1 OAI21X1_79 ( .A(_127_), .B(_128_), .C(_5__2_), .Y(_129_) );
NAND2X1 NAND2X1_80 ( .A(_129_), .B(_133_), .Y(_3__2_) );
OAI21X1 OAI21X1_80 ( .A(_130_), .B(_127_), .C(_132_), .Y(_5__3_) );
INVX1 INVX1_58 ( .A(_5__3_), .Y(_137_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_138_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_139_) );
NAND3X1 NAND3X1_24 ( .A(_137_), .B(_139_), .C(_138_), .Y(_140_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_134_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_135_) );
OAI21X1 OAI21X1_81 ( .A(_134_), .B(_135_), .C(_5__3_), .Y(_136_) );
NAND2X1 NAND2X1_82 ( .A(_136_), .B(_140_), .Y(_3__3_) );
OAI21X1 OAI21X1_82 ( .A(_137_), .B(_134_), .C(_139_), .Y(_1_) );
INVX1 INVX1_59 ( .A(1'b1), .Y(_144_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_145_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_146_) );
NAND3X1 NAND3X1_25 ( .A(_144_), .B(_146_), .C(_145_), .Y(_147_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_141_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_142_) );
OAI21X1 OAI21X1_83 ( .A(_141_), .B(_142_), .C(1'b1), .Y(_143_) );
NAND2X1 NAND2X1_84 ( .A(_143_), .B(_147_), .Y(_4__0_) );
OAI21X1 OAI21X1_84 ( .A(_144_), .B(_141_), .C(_146_), .Y(_6__1_) );
INVX1 INVX1_60 ( .A(_6__1_), .Y(_151_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_152_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_153_) );
NAND3X1 NAND3X1_26 ( .A(_151_), .B(_153_), .C(_152_), .Y(_154_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_148_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_149_) );
OAI21X1 OAI21X1_85 ( .A(_148_), .B(_149_), .C(_6__1_), .Y(_150_) );
NAND2X1 NAND2X1_86 ( .A(_150_), .B(_154_), .Y(_4__1_) );
OAI21X1 OAI21X1_86 ( .A(_151_), .B(_148_), .C(_153_), .Y(_6__2_) );
INVX1 INVX1_61 ( .A(_6__2_), .Y(_158_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_159_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_160_) );
NAND3X1 NAND3X1_27 ( .A(_158_), .B(_160_), .C(_159_), .Y(_161_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_155_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_156_) );
OAI21X1 OAI21X1_87 ( .A(_155_), .B(_156_), .C(_6__2_), .Y(_157_) );
NAND2X1 NAND2X1_88 ( .A(_157_), .B(_161_), .Y(_4__2_) );
OAI21X1 OAI21X1_88 ( .A(_158_), .B(_155_), .C(_160_), .Y(_6__3_) );
INVX1 INVX1_62 ( .A(_6__3_), .Y(_165_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_166_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_167_) );
NAND3X1 NAND3X1_28 ( .A(_165_), .B(_167_), .C(_166_), .Y(_168_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_162_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_163_) );
OAI21X1 OAI21X1_89 ( .A(_162_), .B(_163_), .C(_6__3_), .Y(_164_) );
NAND2X1 NAND2X1_90 ( .A(_164_), .B(_168_), .Y(_4__3_) );
OAI21X1 OAI21X1_90 ( .A(_165_), .B(_162_), .C(_167_), .Y(_2_) );
INVX1 INVX1_63 ( .A(1'b0), .Y(_172_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_173_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_174_) );
NAND3X1 NAND3X1_29 ( .A(_172_), .B(_174_), .C(_173_), .Y(_175_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_169_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_170_) );
OAI21X1 OAI21X1_91 ( .A(_169_), .B(_170_), .C(1'b0), .Y(_171_) );
NAND2X1 NAND2X1_92 ( .A(_171_), .B(_175_), .Y(_9__0_) );
OAI21X1 OAI21X1_92 ( .A(_172_), .B(_169_), .C(_174_), .Y(_11__1_) );
INVX1 INVX1_64 ( .A(_11__1_), .Y(_179_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_180_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_181_) );
NAND3X1 NAND3X1_30 ( .A(_179_), .B(_181_), .C(_180_), .Y(_182_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_176_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_177_) );
OAI21X1 OAI21X1_93 ( .A(_176_), .B(_177_), .C(_11__1_), .Y(_178_) );
NAND2X1 NAND2X1_94 ( .A(_178_), .B(_182_), .Y(_9__1_) );
OAI21X1 OAI21X1_94 ( .A(_179_), .B(_176_), .C(_181_), .Y(_11__2_) );
INVX1 INVX1_65 ( .A(_11__2_), .Y(_186_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_187_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_188_) );
NAND3X1 NAND3X1_31 ( .A(_186_), .B(_188_), .C(_187_), .Y(_189_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_183_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_184_) );
OAI21X1 OAI21X1_95 ( .A(_183_), .B(_184_), .C(_11__2_), .Y(_185_) );
NAND2X1 NAND2X1_96 ( .A(_185_), .B(_189_), .Y(_9__2_) );
OAI21X1 OAI21X1_96 ( .A(_186_), .B(_183_), .C(_188_), .Y(_11__3_) );
INVX1 INVX1_66 ( .A(_11__3_), .Y(_193_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_194_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_195_) );
NAND3X1 NAND3X1_32 ( .A(_193_), .B(_195_), .C(_194_), .Y(_196_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_190_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_191_) );
OAI21X1 OAI21X1_97 ( .A(_190_), .B(_191_), .C(_11__3_), .Y(_192_) );
NAND2X1 NAND2X1_98 ( .A(_192_), .B(_196_), .Y(_9__3_) );
OAI21X1 OAI21X1_98 ( .A(_193_), .B(_190_), .C(_195_), .Y(_7_) );
INVX1 INVX1_67 ( .A(1'b1), .Y(_200_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_201_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_202_) );
NAND3X1 NAND3X1_33 ( .A(_200_), .B(_202_), .C(_201_), .Y(_203_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_197_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_198_) );
OAI21X1 OAI21X1_99 ( .A(_197_), .B(_198_), .C(1'b1), .Y(_199_) );
NAND2X1 NAND2X1_100 ( .A(_199_), .B(_203_), .Y(_10__0_) );
OAI21X1 OAI21X1_100 ( .A(_200_), .B(_197_), .C(_202_), .Y(_12__1_) );
INVX1 INVX1_68 ( .A(_12__1_), .Y(_207_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_208_) );
NAND2X1 NAND2X1_101 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_209_) );
NAND3X1 NAND3X1_34 ( .A(_207_), .B(_209_), .C(_208_), .Y(_210_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_204_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_205_) );
OAI21X1 OAI21X1_101 ( .A(_204_), .B(_205_), .C(_12__1_), .Y(_206_) );
NAND2X1 NAND2X1_102 ( .A(_206_), .B(_210_), .Y(_10__1_) );
OAI21X1 OAI21X1_102 ( .A(_207_), .B(_204_), .C(_209_), .Y(_12__2_) );
INVX1 INVX1_69 ( .A(_12__2_), .Y(_214_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_215_) );
NAND2X1 NAND2X1_103 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_216_) );
NAND3X1 NAND3X1_35 ( .A(_214_), .B(_216_), .C(_215_), .Y(_217_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_211_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_212_) );
OAI21X1 OAI21X1_103 ( .A(_211_), .B(_212_), .C(_12__2_), .Y(_213_) );
NAND2X1 NAND2X1_104 ( .A(_213_), .B(_217_), .Y(_10__2_) );
OAI21X1 OAI21X1_104 ( .A(_214_), .B(_211_), .C(_216_), .Y(_12__3_) );
INVX1 INVX1_70 ( .A(_12__3_), .Y(_221_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_222_) );
NAND2X1 NAND2X1_105 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_223_) );
NAND3X1 NAND3X1_36 ( .A(_221_), .B(_223_), .C(_222_), .Y(_224_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_218_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_219_) );
OAI21X1 OAI21X1_105 ( .A(_218_), .B(_219_), .C(_12__3_), .Y(_220_) );
NAND2X1 NAND2X1_106 ( .A(_220_), .B(_224_), .Y(_10__3_) );
OAI21X1 OAI21X1_106 ( .A(_221_), .B(_218_), .C(_223_), .Y(_8_) );
INVX1 INVX1_71 ( .A(1'b0), .Y(_228_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_229_) );
NAND2X1 NAND2X1_107 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_230_) );
NAND3X1 NAND3X1_37 ( .A(_228_), .B(_230_), .C(_229_), .Y(_231_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_225_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_226_) );
OAI21X1 OAI21X1_107 ( .A(_225_), .B(_226_), .C(1'b0), .Y(_227_) );
NAND2X1 NAND2X1_108 ( .A(_227_), .B(_231_), .Y(_15__0_) );
OAI21X1 OAI21X1_108 ( .A(_228_), .B(_225_), .C(_230_), .Y(_17__1_) );
INVX1 INVX1_72 ( .A(_17__1_), .Y(_235_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_236_) );
NAND2X1 NAND2X1_109 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_237_) );
NAND3X1 NAND3X1_38 ( .A(_235_), .B(_237_), .C(_236_), .Y(_238_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_232_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_233_) );
OAI21X1 OAI21X1_109 ( .A(_232_), .B(_233_), .C(_17__1_), .Y(_234_) );
NAND2X1 NAND2X1_110 ( .A(_234_), .B(_238_), .Y(_15__1_) );
OAI21X1 OAI21X1_110 ( .A(_235_), .B(_232_), .C(_237_), .Y(_17__2_) );
INVX1 INVX1_73 ( .A(_17__2_), .Y(_242_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_243_) );
NAND2X1 NAND2X1_111 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_244_) );
NAND3X1 NAND3X1_39 ( .A(_242_), .B(_244_), .C(_243_), .Y(_245_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_239_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_240_) );
OAI21X1 OAI21X1_111 ( .A(_239_), .B(_240_), .C(_17__2_), .Y(_241_) );
NAND2X1 NAND2X1_112 ( .A(_241_), .B(_245_), .Y(_15__2_) );
OAI21X1 OAI21X1_112 ( .A(_242_), .B(_239_), .C(_244_), .Y(_17__3_) );
INVX1 INVX1_74 ( .A(_17__3_), .Y(_249_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_250_) );
NAND2X1 NAND2X1_113 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_251_) );
NAND3X1 NAND3X1_40 ( .A(_249_), .B(_251_), .C(_250_), .Y(_252_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_246_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_247_) );
OAI21X1 OAI21X1_113 ( .A(_246_), .B(_247_), .C(_17__3_), .Y(_248_) );
NAND2X1 NAND2X1_114 ( .A(_248_), .B(_252_), .Y(_15__3_) );
OAI21X1 OAI21X1_114 ( .A(_249_), .B(_246_), .C(_251_), .Y(_13_) );
INVX1 INVX1_75 ( .A(1'b1), .Y(_256_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_257_) );
NAND2X1 NAND2X1_115 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_258_) );
NAND3X1 NAND3X1_41 ( .A(_256_), .B(_258_), .C(_257_), .Y(_259_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_253_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_254_) );
OAI21X1 OAI21X1_115 ( .A(_253_), .B(_254_), .C(1'b1), .Y(_255_) );
NAND2X1 NAND2X1_116 ( .A(_255_), .B(_259_), .Y(_16__0_) );
OAI21X1 OAI21X1_116 ( .A(_256_), .B(_253_), .C(_258_), .Y(_18__1_) );
INVX1 INVX1_76 ( .A(_18__1_), .Y(_263_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_264_) );
NAND2X1 NAND2X1_117 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_265_) );
NAND3X1 NAND3X1_42 ( .A(_263_), .B(_265_), .C(_264_), .Y(_266_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_260_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_261_) );
OAI21X1 OAI21X1_117 ( .A(_260_), .B(_261_), .C(_18__1_), .Y(_262_) );
NAND2X1 NAND2X1_118 ( .A(_262_), .B(_266_), .Y(_16__1_) );
OAI21X1 OAI21X1_118 ( .A(_263_), .B(_260_), .C(_265_), .Y(_18__2_) );
INVX1 INVX1_77 ( .A(_18__2_), .Y(_270_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_271_) );
NAND2X1 NAND2X1_119 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_272_) );
NAND3X1 NAND3X1_43 ( .A(_270_), .B(_272_), .C(_271_), .Y(_273_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_267_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_268_) );
OAI21X1 OAI21X1_119 ( .A(_267_), .B(_268_), .C(_18__2_), .Y(_269_) );
NAND2X1 NAND2X1_120 ( .A(_269_), .B(_273_), .Y(_16__2_) );
OAI21X1 OAI21X1_120 ( .A(_270_), .B(_267_), .C(_272_), .Y(_18__3_) );
INVX1 INVX1_78 ( .A(_18__3_), .Y(_277_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_278_) );
NAND2X1 NAND2X1_121 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_279_) );
NAND3X1 NAND3X1_44 ( .A(_277_), .B(_279_), .C(_278_), .Y(_280_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_274_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_275_) );
OAI21X1 OAI21X1_121 ( .A(_274_), .B(_275_), .C(_18__3_), .Y(_276_) );
NAND2X1 NAND2X1_122 ( .A(_276_), .B(_280_), .Y(_16__3_) );
OAI21X1 OAI21X1_122 ( .A(_277_), .B(_274_), .C(_279_), .Y(_14_) );
INVX1 INVX1_79 ( .A(1'b0), .Y(_284_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_285_) );
NAND2X1 NAND2X1_123 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_286_) );
NAND3X1 NAND3X1_45 ( .A(_284_), .B(_286_), .C(_285_), .Y(_287_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_281_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_282_) );
OAI21X1 OAI21X1_123 ( .A(_281_), .B(_282_), .C(1'b0), .Y(_283_) );
NAND2X1 NAND2X1_124 ( .A(_283_), .B(_287_), .Y(_21__0_) );
OAI21X1 OAI21X1_124 ( .A(_284_), .B(_281_), .C(_286_), .Y(_23__1_) );
INVX1 INVX1_80 ( .A(_23__1_), .Y(_291_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_292_) );
NAND2X1 NAND2X1_125 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_293_) );
NAND3X1 NAND3X1_46 ( .A(_291_), .B(_293_), .C(_292_), .Y(_294_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_288_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_289_) );
OAI21X1 OAI21X1_125 ( .A(_288_), .B(_289_), .C(_23__1_), .Y(_290_) );
NAND2X1 NAND2X1_126 ( .A(_290_), .B(_294_), .Y(_21__1_) );
OAI21X1 OAI21X1_126 ( .A(_291_), .B(_288_), .C(_293_), .Y(_23__2_) );
INVX1 INVX1_81 ( .A(_23__2_), .Y(_298_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_299_) );
NAND2X1 NAND2X1_127 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_300_) );
NAND3X1 NAND3X1_47 ( .A(_298_), .B(_300_), .C(_299_), .Y(_301_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_295_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_296_) );
OAI21X1 OAI21X1_127 ( .A(_295_), .B(_296_), .C(_23__2_), .Y(_297_) );
NAND2X1 NAND2X1_128 ( .A(_297_), .B(_301_), .Y(_21__2_) );
OAI21X1 OAI21X1_128 ( .A(_298_), .B(_295_), .C(_300_), .Y(_23__3_) );
INVX1 INVX1_82 ( .A(_23__3_), .Y(_305_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_306_) );
NAND2X1 NAND2X1_129 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_307_) );
NAND3X1 NAND3X1_48 ( .A(_305_), .B(_307_), .C(_306_), .Y(_308_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_302_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_303_) );
OAI21X1 OAI21X1_129 ( .A(_302_), .B(_303_), .C(_23__3_), .Y(_304_) );
NAND2X1 NAND2X1_130 ( .A(_304_), .B(_308_), .Y(_21__3_) );
OAI21X1 OAI21X1_130 ( .A(_305_), .B(_302_), .C(_307_), .Y(_19_) );
INVX1 INVX1_83 ( .A(1'b1), .Y(_312_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_313_) );
NAND2X1 NAND2X1_131 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_314_) );
NAND3X1 NAND3X1_49 ( .A(_312_), .B(_314_), .C(_313_), .Y(_315_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_309_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_310_) );
OAI21X1 OAI21X1_131 ( .A(_309_), .B(_310_), .C(1'b1), .Y(_311_) );
NAND2X1 NAND2X1_132 ( .A(_311_), .B(_315_), .Y(_22__0_) );
OAI21X1 OAI21X1_132 ( .A(_312_), .B(_309_), .C(_314_), .Y(_24__1_) );
INVX1 INVX1_84 ( .A(_24__1_), .Y(_319_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_320_) );
NAND2X1 NAND2X1_133 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_321_) );
NAND3X1 NAND3X1_50 ( .A(_319_), .B(_321_), .C(_320_), .Y(_322_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_316_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_317_) );
OAI21X1 OAI21X1_133 ( .A(_316_), .B(_317_), .C(_24__1_), .Y(_318_) );
NAND2X1 NAND2X1_134 ( .A(_318_), .B(_322_), .Y(_22__1_) );
OAI21X1 OAI21X1_134 ( .A(_319_), .B(_316_), .C(_321_), .Y(_24__2_) );
INVX1 INVX1_85 ( .A(_24__2_), .Y(_326_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_327_) );
NAND2X1 NAND2X1_135 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_328_) );
NAND3X1 NAND3X1_51 ( .A(_326_), .B(_328_), .C(_327_), .Y(_329_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_323_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_324_) );
OAI21X1 OAI21X1_135 ( .A(_323_), .B(_324_), .C(_24__2_), .Y(_325_) );
NAND2X1 NAND2X1_136 ( .A(_325_), .B(_329_), .Y(_22__2_) );
OAI21X1 OAI21X1_136 ( .A(_326_), .B(_323_), .C(_328_), .Y(_24__3_) );
INVX1 INVX1_86 ( .A(_24__3_), .Y(_333_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_334_) );
NAND2X1 NAND2X1_137 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_335_) );
NAND3X1 NAND3X1_52 ( .A(_333_), .B(_335_), .C(_334_), .Y(_336_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_330_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_331_) );
OAI21X1 OAI21X1_137 ( .A(_330_), .B(_331_), .C(_24__3_), .Y(_332_) );
NAND2X1 NAND2X1_138 ( .A(_332_), .B(_336_), .Y(_22__3_) );
OAI21X1 OAI21X1_138 ( .A(_333_), .B(_330_), .C(_335_), .Y(_20_) );
INVX1 INVX1_87 ( .A(1'b0), .Y(_340_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_341_) );
NAND2X1 NAND2X1_139 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_342_) );
NAND3X1 NAND3X1_53 ( .A(_340_), .B(_342_), .C(_341_), .Y(_343_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_337_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_338_) );
OAI21X1 OAI21X1_139 ( .A(_337_), .B(_338_), .C(1'b0), .Y(_339_) );
NAND2X1 NAND2X1_140 ( .A(_339_), .B(_343_), .Y(_27__0_) );
OAI21X1 OAI21X1_140 ( .A(_340_), .B(_337_), .C(_342_), .Y(_29__1_) );
INVX1 INVX1_88 ( .A(_29__1_), .Y(_347_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_348_) );
NAND2X1 NAND2X1_141 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_349_) );
NAND3X1 NAND3X1_54 ( .A(_347_), .B(_349_), .C(_348_), .Y(_350_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_344_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_345_) );
OAI21X1 OAI21X1_141 ( .A(_344_), .B(_345_), .C(_29__1_), .Y(_346_) );
NAND2X1 NAND2X1_142 ( .A(_346_), .B(_350_), .Y(_27__1_) );
OAI21X1 OAI21X1_142 ( .A(_347_), .B(_344_), .C(_349_), .Y(_29__2_) );
INVX1 INVX1_89 ( .A(_29__2_), .Y(_354_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_355_) );
NAND2X1 NAND2X1_143 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_356_) );
NAND3X1 NAND3X1_55 ( .A(_354_), .B(_356_), .C(_355_), .Y(_357_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_351_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_352_) );
OAI21X1 OAI21X1_143 ( .A(_351_), .B(_352_), .C(_29__2_), .Y(_353_) );
NAND2X1 NAND2X1_144 ( .A(_353_), .B(_357_), .Y(_27__2_) );
OAI21X1 OAI21X1_144 ( .A(_354_), .B(_351_), .C(_356_), .Y(_29__3_) );
INVX1 INVX1_90 ( .A(_29__3_), .Y(_361_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_362_) );
NAND2X1 NAND2X1_145 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_363_) );
NAND3X1 NAND3X1_56 ( .A(_361_), .B(_363_), .C(_362_), .Y(_364_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_358_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_359_) );
OAI21X1 OAI21X1_145 ( .A(_358_), .B(_359_), .C(_29__3_), .Y(_360_) );
NAND2X1 NAND2X1_146 ( .A(_360_), .B(_364_), .Y(_27__3_) );
OAI21X1 OAI21X1_146 ( .A(_361_), .B(_358_), .C(_363_), .Y(_25_) );
INVX1 INVX1_91 ( .A(1'b1), .Y(_368_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_369_) );
NAND2X1 NAND2X1_147 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_370_) );
NAND3X1 NAND3X1_57 ( .A(_368_), .B(_370_), .C(_369_), .Y(_371_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_365_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_366_) );
OAI21X1 OAI21X1_147 ( .A(_365_), .B(_366_), .C(1'b1), .Y(_367_) );
NAND2X1 NAND2X1_148 ( .A(_367_), .B(_371_), .Y(_28__0_) );
OAI21X1 OAI21X1_148 ( .A(_368_), .B(_365_), .C(_370_), .Y(_30__1_) );
INVX1 INVX1_92 ( .A(_30__1_), .Y(_375_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_376_) );
NAND2X1 NAND2X1_149 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_377_) );
NAND3X1 NAND3X1_58 ( .A(_375_), .B(_377_), .C(_376_), .Y(_378_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_372_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_373_) );
OAI21X1 OAI21X1_149 ( .A(_372_), .B(_373_), .C(_30__1_), .Y(_374_) );
NAND2X1 NAND2X1_150 ( .A(_374_), .B(_378_), .Y(_28__1_) );
OAI21X1 OAI21X1_150 ( .A(_375_), .B(_372_), .C(_377_), .Y(_30__2_) );
INVX1 INVX1_93 ( .A(_30__2_), .Y(_382_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_383_) );
NAND2X1 NAND2X1_151 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_384_) );
BUFX2 BUFX2_32 ( .A(1'b0), .Y(_5__0_) );
BUFX2 BUFX2_33 ( .A(_1_), .Y(_5__4_) );
BUFX2 BUFX2_34 ( .A(1'b1), .Y(_6__0_) );
BUFX2 BUFX2_35 ( .A(_2_), .Y(_6__4_) );
BUFX2 BUFX2_36 ( .A(1'b0), .Y(_11__0_) );
BUFX2 BUFX2_37 ( .A(_7_), .Y(_11__4_) );
BUFX2 BUFX2_38 ( .A(1'b1), .Y(_12__0_) );
BUFX2 BUFX2_39 ( .A(_8_), .Y(_12__4_) );
BUFX2 BUFX2_40 ( .A(1'b0), .Y(_17__0_) );
BUFX2 BUFX2_41 ( .A(_13_), .Y(_17__4_) );
BUFX2 BUFX2_42 ( .A(1'b1), .Y(_18__0_) );
BUFX2 BUFX2_43 ( .A(_14_), .Y(_18__4_) );
BUFX2 BUFX2_44 ( .A(1'b0), .Y(_23__0_) );
BUFX2 BUFX2_45 ( .A(_19_), .Y(_23__4_) );
BUFX2 BUFX2_46 ( .A(1'b1), .Y(_24__0_) );
BUFX2 BUFX2_47 ( .A(_20_), .Y(_24__4_) );
BUFX2 BUFX2_48 ( .A(1'b0), .Y(_29__0_) );
BUFX2 BUFX2_49 ( .A(_25_), .Y(_29__4_) );
BUFX2 BUFX2_50 ( .A(1'b1), .Y(_30__0_) );
BUFX2 BUFX2_51 ( .A(_26_), .Y(_30__4_) );
BUFX2 BUFX2_52 ( .A(1'b0), .Y(_35__0_) );
BUFX2 BUFX2_53 ( .A(_31_), .Y(_35__4_) );
BUFX2 BUFX2_54 ( .A(1'b1), .Y(_36__0_) );
BUFX2 BUFX2_55 ( .A(_32_), .Y(_36__4_) );
BUFX2 BUFX2_56 ( .A(1'b0), .Y(_41__0_) );
BUFX2 BUFX2_57 ( .A(_37_), .Y(_41__4_) );
BUFX2 BUFX2_58 ( .A(1'b1), .Y(_42__0_) );
BUFX2 BUFX2_59 ( .A(_38_), .Y(_42__4_) );
BUFX2 BUFX2_60 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_61 ( .A(1'b0), .Y(w_cout_0_) );
endmodule
