module cla_62bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [61:0] i_add1;
input [61:0] i_add2;
output [62:0] o_result;

NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_213_), .C(_209_), .Y(_214_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .C(_214_), .Y(_215_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_215_), .Y(w_C_37_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .Y(_216_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add1[37]), .Y(_217_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_218_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_218_), .Y(_219_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_220_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_220_), .Y(_221_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_221_), .C(_214_), .Y(_222_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_217_), .C(_222_), .Y(w_C_38_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_217_), .Y(_223_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_223_), .Y(_224_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_225_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_225_), .Y(_226_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_226_), .C(_222_), .Y(_227_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .C(_227_), .Y(_228_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_228_), .Y(w_C_39_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .Y(_229_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add1[39]), .Y(_230_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_231_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_231_), .Y(_232_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_233_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_233_), .Y(_234_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_234_), .C(_227_), .Y(_235_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_230_), .C(_235_), .Y(w_C_40_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_230_), .Y(_236_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_236_), .Y(_237_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_238_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_238_), .Y(_239_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_239_), .C(_235_), .Y(_240_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .C(_240_), .Y(_241_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_241_), .Y(w_C_41_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .Y(_242_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add1[41]), .Y(_243_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_244_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_244_), .Y(_245_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_246_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_246_), .Y(_247_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_247_), .C(_240_), .Y(_248_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_243_), .C(_248_), .Y(w_C_42_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_243_), .Y(_249_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_249_), .Y(_250_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_251_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_251_), .Y(_252_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_252_), .C(_248_), .Y(_253_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .C(_253_), .Y(_254_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_254_), .Y(w_C_43_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .Y(_255_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add1[43]), .Y(_256_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_257_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_257_), .Y(_258_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_259_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_259_), .Y(_260_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_260_), .C(_253_), .Y(_261_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_256_), .C(_261_), .Y(w_C_44_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_256_), .Y(_262_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_262_), .Y(_263_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_264_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_264_), .Y(_265_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_265_), .C(_261_), .Y(_266_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .C(_266_), .Y(_267_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_267_), .Y(w_C_45_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .Y(_268_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add1[45]), .Y(_269_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_270_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_270_), .Y(_271_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_272_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_272_), .Y(_273_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_273_), .C(_266_), .Y(_274_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_269_), .C(_274_), .Y(w_C_46_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_269_), .Y(_275_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_275_), .Y(_276_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_277_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_277_), .Y(_278_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_278_), .C(_274_), .Y(_279_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .C(_279_), .Y(_280_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_280_), .Y(w_C_47_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .Y(_281_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add1[47]), .Y(_282_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_283_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_283_), .Y(_284_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_285_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_285_), .Y(_286_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_286_), .C(_279_), .Y(_287_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_282_), .C(_287_), .Y(w_C_48_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_282_), .Y(_288_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_288_), .Y(_289_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_290_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_290_), .Y(_291_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_291_), .C(_287_), .Y(_292_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .C(_292_), .Y(_293_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_293_), .Y(w_C_49_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .Y(_294_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add1[49]), .Y(_295_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_296_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_296_), .Y(_297_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_298_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_298_), .Y(_299_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_299_), .C(_292_), .Y(_300_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_295_), .C(_300_), .Y(w_C_50_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_301_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_301_), .Y(_302_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_295_), .Y(_303_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_303_), .Y(_304_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_305_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_305_), .C(_300_), .Y(_306_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_302_), .Y(w_C_51_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .Y(_307_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add1[51]), .Y(_308_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_308_), .Y(_309_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_309_), .C(_306_), .Y(_310_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_308_), .C(_310_), .Y(w_C_52_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .Y(_311_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add1[52]), .Y(_312_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .C(w_C_52_), .Y(_313_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_312_), .C(_313_), .Y(w_C_53_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .Y(_314_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add1[53]), .Y(_315_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_315_), .Y(_316_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(w_C_53_), .B(_316_), .Y(_317_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .C(_317_), .Y(_318_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_318_), .Y(w_C_54_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_319_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_320_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_318_), .C(_319_), .Y(w_C_55_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .Y(_321_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add1[55]), .Y(_322_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_320_), .Y(_323_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_316_), .Y(_324_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_312_), .Y(_325_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_326_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_327_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_327_), .C(_310_), .Y(_328_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_315_), .Y(_329_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_329_), .C(_328_), .Y(_330_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_319_), .C(_330_), .Y(_331_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_322_), .Y(_332_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_332_), .C(_331_), .Y(_333_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_322_), .C(_333_), .Y(w_C_56_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .Y(_334_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add1[56]), .Y(_335_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .C(w_C_56_), .Y(_336_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_335_), .C(_336_), .Y(w_C_57_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_335_), .Y(_337_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_337_), .Y(_338_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_339_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_339_), .Y(_340_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_340_), .C(_336_), .Y(_341_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .C(_341_), .Y(_342_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_342_), .Y(w_C_58_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_343_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_344_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_342_), .C(_343_), .Y(w_C_59_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_345_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_344_), .Y(_346_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_347_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_347_), .Y(_348_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_322_), .Y(_349_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_349_), .Y(_350_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_338_), .C(_333_), .Y(_351_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_352_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_352_), .Y(_353_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_353_), .C(_351_), .Y(_354_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_343_), .C(_354_), .Y(_355_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_356_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_356_), .C(_355_), .Y(_357_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_357_), .Y(w_C_60_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[60]), .B(i_add1[60]), .Y(_358_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[60]), .B(i_add1[60]), .Y(_359_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_359_), .C(_357_), .Y(_360_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_358_), .Y(w_C_61_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[61]), .B(i_add1[61]), .Y(_361_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[61]), .B(i_add1[61]), .Y(_362_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_358_), .B(_362_), .C(_360_), .Y(_363_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_363_), .Y(w_C_62_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_2_), .Y(w_C_2_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .Y(_3_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add1[2]), .Y(_4_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_2_), .C(_6_), .Y(_7_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_9_), .C(_7_), .Y(_10_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_10_), .Y(w_C_4_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(_12_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_13_), .C(_10_), .Y(_14_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_12_), .Y(w_C_5_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .Y(_15_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add1[5]), .Y(_16_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_17_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_17_), .Y(_18_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_18_), .C(_14_), .Y(_19_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_16_), .C(_19_), .Y(w_C_6_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_20_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_20_), .Y(_21_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_16_), .Y(_22_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_23_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_24_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(_24_), .Y(_25_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_25_), .C(_19_), .Y(_26_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_21_), .Y(w_C_7_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .Y(_27_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add1[7]), .Y(_28_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_29_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_29_), .Y(_30_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_30_), .C(_26_), .Y(_31_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_28_), .C(_31_), .Y(w_C_8_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_32_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_32_), .Y(_33_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_28_), .Y(_34_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(_34_), .Y(_35_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_36_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_36_), .Y(_37_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_37_), .C(_31_), .Y(_38_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_33_), .Y(w_C_9_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_39_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_364__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_364__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_364__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_364__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_364__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_364__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_364__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_364__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_364__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_364__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_364__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_364__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_364__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_364__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_364__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_364__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_364__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_364__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_364__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_364__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_364__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_364__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_364__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_364__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_364__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_364__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_364__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_364__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_364__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_364__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_364__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_364__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_364__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_364__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_364__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_364__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_364__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_364__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_364__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_364__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_364__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_364__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_364__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_364__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_364__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_364__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_364__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_364__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_364__48_), .Y(o_result[48]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_364__49_), .Y(o_result[49]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_364__50_), .Y(o_result[50]) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_364__51_), .Y(o_result[51]) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(_364__52_), .Y(o_result[52]) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(_364__53_), .Y(o_result[53]) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(_364__54_), .Y(o_result[54]) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_364__55_), .Y(o_result[55]) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_364__56_), .Y(o_result[56]) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_364__57_), .Y(o_result[57]) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_364__58_), .Y(o_result[58]) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(_364__59_), .Y(o_result[59]) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(_364__60_), .Y(o_result[60]) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(_364__61_), .Y(o_result[61]) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(w_C_62_), .Y(o_result[62]) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_368_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_369_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_370_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_370_), .C(_369_), .Y(_371_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_365_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_366_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_365_), .B(_366_), .C(w_C_4_), .Y(_367_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_371_), .Y(_364__4_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_375_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_376_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_377_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_377_), .C(_376_), .Y(_378_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_372_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_373_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_373_), .C(w_C_5_), .Y(_374_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_378_), .Y(_364__5_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_382_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_383_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_384_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_382_), .B(_384_), .C(_383_), .Y(_385_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_379_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_380_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_380_), .C(w_C_6_), .Y(_381_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_385_), .Y(_364__6_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_389_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_390_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_391_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_391_), .C(_390_), .Y(_392_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_386_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_387_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_387_), .C(w_C_7_), .Y(_388_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(_392_), .Y(_364__7_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_396_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_397_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_398_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_398_), .C(_397_), .Y(_399_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_393_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_394_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_394_), .C(w_C_8_), .Y(_395_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_399_), .Y(_364__8_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_403_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_404_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_405_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_405_), .C(_404_), .Y(_406_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_400_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_401_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_400_), .B(_401_), .C(w_C_9_), .Y(_402_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_406_), .Y(_364__9_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_410_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_411_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_412_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(_412_), .C(_411_), .Y(_413_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_407_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_408_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_408_), .C(w_C_10_), .Y(_409_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_413_), .Y(_364__10_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_417_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_418_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_419_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_419_), .C(_418_), .Y(_420_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_414_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_415_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_414_), .B(_415_), .C(w_C_11_), .Y(_416_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_420_), .Y(_364__11_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(w_C_12_), .Y(_424_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_425_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_426_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_426_), .C(_425_), .Y(_427_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_421_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_422_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_422_), .C(w_C_12_), .Y(_423_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_427_), .Y(_364__12_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(w_C_13_), .Y(_431_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_432_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_433_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_433_), .C(_432_), .Y(_434_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_428_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_429_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_429_), .C(w_C_13_), .Y(_430_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_434_), .Y(_364__13_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(w_C_14_), .Y(_438_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_439_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_440_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_440_), .C(_439_), .Y(_441_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_435_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_436_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_436_), .C(w_C_14_), .Y(_437_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_441_), .Y(_364__14_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(_445_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_446_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_447_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_445_), .B(_447_), .C(_446_), .Y(_448_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_442_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_443_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_443_), .C(w_C_15_), .Y(_444_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_448_), .Y(_364__15_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(w_C_16_), .Y(_452_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_453_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_454_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_454_), .C(_453_), .Y(_455_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_449_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_450_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_450_), .C(w_C_16_), .Y(_451_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_455_), .Y(_364__16_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(w_C_17_), .Y(_459_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_460_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_461_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_461_), .C(_460_), .Y(_462_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_456_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_457_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_456_), .B(_457_), .C(w_C_17_), .Y(_458_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_462_), .Y(_364__17_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(w_C_18_), .Y(_466_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_467_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_468_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_466_), .B(_468_), .C(_467_), .Y(_469_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_463_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_464_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_464_), .C(w_C_18_), .Y(_465_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_469_), .Y(_364__18_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(w_C_19_), .Y(_473_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_474_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_475_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_475_), .C(_474_), .Y(_476_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_470_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_471_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_470_), .B(_471_), .C(w_C_19_), .Y(_472_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_476_), .Y(_364__19_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(w_C_20_), .Y(_480_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_481_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_482_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_482_), .C(_481_), .Y(_483_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_477_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_478_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_477_), .B(_478_), .C(w_C_20_), .Y(_479_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_483_), .Y(_364__20_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(w_C_21_), .Y(_487_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_488_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_489_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_489_), .C(_488_), .Y(_490_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_484_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_485_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_484_), .B(_485_), .C(w_C_21_), .Y(_486_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_490_), .Y(_364__21_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(w_C_22_), .Y(_494_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_495_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_496_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_496_), .C(_495_), .Y(_497_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_491_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_492_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_492_), .C(w_C_22_), .Y(_493_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_497_), .Y(_364__22_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(w_C_23_), .Y(_501_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_502_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_503_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_501_), .B(_503_), .C(_502_), .Y(_504_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_498_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_499_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_499_), .C(w_C_23_), .Y(_500_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_504_), .Y(_364__23_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(w_C_24_), .Y(_508_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_509_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_510_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_510_), .C(_509_), .Y(_511_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_505_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_506_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(_506_), .C(w_C_24_), .Y(_507_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_511_), .Y(_364__24_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(w_C_25_), .Y(_515_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_516_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_517_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_517_), .C(_516_), .Y(_518_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_512_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_513_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_513_), .C(w_C_25_), .Y(_514_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_518_), .Y(_364__25_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(w_C_26_), .Y(_522_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_523_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_524_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_522_), .B(_524_), .C(_523_), .Y(_525_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_519_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_520_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_520_), .C(w_C_26_), .Y(_521_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_525_), .Y(_364__26_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(w_C_27_), .Y(_529_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_530_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_531_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_531_), .C(_530_), .Y(_532_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_526_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_527_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_527_), .C(w_C_27_), .Y(_528_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_532_), .Y(_364__27_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(w_C_28_), .Y(_536_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_537_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_538_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_536_), .B(_538_), .C(_537_), .Y(_539_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_533_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_534_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_534_), .C(w_C_28_), .Y(_535_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_539_), .Y(_364__28_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(w_C_29_), .Y(_543_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_544_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_545_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_545_), .C(_544_), .Y(_546_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_540_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_541_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_541_), .C(w_C_29_), .Y(_542_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_542_), .B(_546_), .Y(_364__29_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(w_C_30_), .Y(_550_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_551_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_552_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_550_), .B(_552_), .C(_551_), .Y(_553_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_547_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_548_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_548_), .C(w_C_30_), .Y(_549_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(_553_), .Y(_364__30_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(w_C_31_), .Y(_557_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_558_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_559_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_557_), .B(_559_), .C(_558_), .Y(_560_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_554_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_555_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_555_), .C(w_C_31_), .Y(_556_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_556_), .B(_560_), .Y(_364__31_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(w_C_32_), .Y(_564_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_565_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_566_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_564_), .B(_566_), .C(_565_), .Y(_567_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_561_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_562_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_562_), .C(w_C_32_), .Y(_563_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(_567_), .Y(_364__32_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(w_C_33_), .Y(_571_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_572_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_573_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_573_), .C(_572_), .Y(_574_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_568_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_569_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_569_), .C(w_C_33_), .Y(_570_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_574_), .Y(_364__33_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(w_C_34_), .Y(_578_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_579_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_580_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_578_), .B(_580_), .C(_579_), .Y(_581_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_575_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_576_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_576_), .C(w_C_34_), .Y(_577_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_581_), .Y(_364__34_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(w_C_35_), .Y(_585_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_586_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_587_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_585_), .B(_587_), .C(_586_), .Y(_588_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_582_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_583_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_583_), .C(w_C_35_), .Y(_584_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_588_), .Y(_364__35_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(w_C_36_), .Y(_592_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_593_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_594_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_592_), .B(_594_), .C(_593_), .Y(_595_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_589_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_590_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_589_), .B(_590_), .C(w_C_36_), .Y(_591_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_595_), .Y(_364__36_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(w_C_37_), .Y(_599_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_600_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_601_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_599_), .B(_601_), .C(_600_), .Y(_602_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_596_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_597_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_597_), .C(w_C_37_), .Y(_598_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_598_), .B(_602_), .Y(_364__37_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(w_C_38_), .Y(_606_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_607_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_608_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_608_), .C(_607_), .Y(_609_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_603_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_604_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_603_), .B(_604_), .C(w_C_38_), .Y(_605_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_609_), .Y(_364__38_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(w_C_39_), .Y(_613_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_614_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_615_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_613_), .B(_615_), .C(_614_), .Y(_616_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_610_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_611_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_611_), .C(w_C_39_), .Y(_612_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_612_), .B(_616_), .Y(_364__39_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(w_C_40_), .Y(_620_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_621_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_622_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_622_), .C(_621_), .Y(_623_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_617_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_618_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_617_), .B(_618_), .C(w_C_40_), .Y(_619_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_623_), .Y(_364__40_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(w_C_41_), .Y(_627_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_628_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_629_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(_629_), .C(_628_), .Y(_630_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_624_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_625_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_624_), .B(_625_), .C(w_C_41_), .Y(_626_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_630_), .Y(_364__41_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(w_C_42_), .Y(_634_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_635_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_636_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_634_), .B(_636_), .C(_635_), .Y(_637_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_631_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_632_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_631_), .B(_632_), .C(w_C_42_), .Y(_633_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_637_), .Y(_364__42_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(w_C_43_), .Y(_641_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_642_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_643_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_641_), .B(_643_), .C(_642_), .Y(_644_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_638_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_639_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_639_), .C(w_C_43_), .Y(_640_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(_644_), .Y(_364__43_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(w_C_44_), .Y(_648_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_649_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_650_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_650_), .C(_649_), .Y(_651_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_645_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_646_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_645_), .B(_646_), .C(w_C_44_), .Y(_647_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_647_), .B(_651_), .Y(_364__44_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(w_C_45_), .Y(_655_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_656_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_657_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_657_), .C(_656_), .Y(_658_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_652_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_653_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_653_), .C(w_C_45_), .Y(_654_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_658_), .Y(_364__45_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(w_C_46_), .Y(_662_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_663_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_664_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_664_), .C(_663_), .Y(_665_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_659_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_660_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(_660_), .C(w_C_46_), .Y(_661_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_661_), .B(_665_), .Y(_364__46_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(w_C_47_), .Y(_669_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_670_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_671_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_669_), .B(_671_), .C(_670_), .Y(_672_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_666_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_667_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_666_), .B(_667_), .C(w_C_47_), .Y(_668_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_672_), .Y(_364__47_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(w_C_48_), .Y(_676_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_677_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_678_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_676_), .B(_678_), .C(_677_), .Y(_679_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_673_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_674_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(_674_), .C(w_C_48_), .Y(_675_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_679_), .Y(_364__48_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(w_C_49_), .Y(_683_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_684_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_685_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_683_), .B(_685_), .C(_684_), .Y(_686_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_680_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_681_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_680_), .B(_681_), .C(w_C_49_), .Y(_682_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_682_), .B(_686_), .Y(_364__49_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(w_C_50_), .Y(_690_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_691_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_692_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_690_), .B(_692_), .C(_691_), .Y(_693_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_687_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_688_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_687_), .B(_688_), .C(w_C_50_), .Y(_689_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_693_), .Y(_364__50_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(w_C_51_), .Y(_697_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_698_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_699_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_697_), .B(_699_), .C(_698_), .Y(_700_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_694_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_695_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_695_), .C(w_C_51_), .Y(_696_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_700_), .Y(_364__51_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(w_C_52_), .Y(_704_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_705_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_706_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_706_), .C(_705_), .Y(_707_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_701_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_702_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_701_), .B(_702_), .C(w_C_52_), .Y(_703_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_707_), .Y(_364__52_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(w_C_53_), .Y(_711_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_712_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_713_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_713_), .C(_712_), .Y(_714_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_708_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_709_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_708_), .B(_709_), .C(w_C_53_), .Y(_710_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_710_), .B(_714_), .Y(_364__53_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(w_C_54_), .Y(_718_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_719_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_720_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_718_), .B(_720_), .C(_719_), .Y(_721_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_715_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_716_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(_716_), .C(w_C_54_), .Y(_717_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_717_), .B(_721_), .Y(_364__54_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(w_C_55_), .Y(_725_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_726_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_727_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(_727_), .C(_726_), .Y(_728_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_722_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_723_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_722_), .B(_723_), .C(w_C_55_), .Y(_724_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_724_), .B(_728_), .Y(_364__55_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(w_C_56_), .Y(_732_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_733_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_734_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_734_), .C(_733_), .Y(_735_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_729_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_730_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_730_), .C(w_C_56_), .Y(_731_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_731_), .B(_735_), .Y(_364__56_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(w_C_57_), .Y(_739_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_740_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_741_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_739_), .B(_741_), .C(_740_), .Y(_742_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_736_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_737_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_736_), .B(_737_), .C(w_C_57_), .Y(_738_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_738_), .B(_742_), .Y(_364__57_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(w_C_58_), .Y(_746_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_747_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_748_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_748_), .C(_747_), .Y(_749_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_743_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_744_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_743_), .B(_744_), .C(w_C_58_), .Y(_745_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_745_), .B(_749_), .Y(_364__58_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(w_C_59_), .Y(_753_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_754_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_755_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_753_), .B(_755_), .C(_754_), .Y(_756_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_750_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_751_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_750_), .B(_751_), .C(w_C_59_), .Y(_752_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(_756_), .Y(_364__59_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(w_C_60_), .Y(_760_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[60]), .B(i_add1[60]), .Y(_761_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(i_add2[60]), .B(i_add1[60]), .Y(_762_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_760_), .B(_762_), .C(_761_), .Y(_763_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[60]), .B(i_add1[60]), .Y(_757_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[60]), .B(i_add1[60]), .Y(_758_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_757_), .B(_758_), .C(w_C_60_), .Y(_759_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_759_), .B(_763_), .Y(_364__60_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(w_C_61_), .Y(_767_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[61]), .B(i_add1[61]), .Y(_768_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(i_add2[61]), .B(i_add1[61]), .Y(_769_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_767_), .B(_769_), .C(_768_), .Y(_770_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add2[61]), .B(i_add1[61]), .Y(_764_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[61]), .B(i_add1[61]), .Y(_765_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_764_), .B(_765_), .C(w_C_61_), .Y(_766_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_766_), .B(_770_), .Y(_364__61_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_774_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_775_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_776_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_774_), .B(_776_), .C(_775_), .Y(_777_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_771_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_772_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_771_), .B(_772_), .C(gnd), .Y(_773_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_777_), .Y(_364__0_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_781_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_782_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_783_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_781_), .B(_783_), .C(_782_), .Y(_784_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_778_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_779_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(_779_), .C(w_C_1_), .Y(_780_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_780_), .B(_784_), .Y(_364__1_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_788_) );
OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_789_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_790_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_790_), .C(_789_), .Y(_791_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_785_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_786_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_786_), .C(w_C_2_), .Y(_787_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_791_), .Y(_364__2_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_795_) );
OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_796_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_797_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_795_), .B(_797_), .C(_796_), .Y(_798_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_792_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_793_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_792_), .B(_793_), .C(w_C_3_), .Y(_794_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_798_), .Y(_364__3_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(_39_), .Y(_40_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_41_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(_41_), .Y(_42_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_42_), .C(_38_), .Y(_43_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_40_), .Y(_44_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(_44_), .Y(w_C_10_) );
AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_45_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(_45_), .Y(_46_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_47_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_44_), .C(_46_), .Y(w_C_11_) );
AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_48_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(_48_), .Y(_49_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(_47_), .Y(_50_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_46_), .C(_43_), .Y(_51_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_52_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(_52_), .Y(_53_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_53_), .C(_51_), .Y(_54_) );
AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_49_), .Y(_55_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(_55_), .Y(w_C_12_) );
AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_56_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(_56_), .Y(_57_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_57_), .C(_54_), .Y(_58_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .C(_58_), .Y(_59_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(_59_), .Y(w_C_13_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .Y(_60_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(i_add1[13]), .Y(_61_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_62_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(_62_), .Y(_63_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_64_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(_64_), .Y(_65_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_65_), .C(_58_), .Y(_66_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_61_), .C(_66_), .Y(w_C_14_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_61_), .Y(_67_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(_67_), .Y(_68_) );
AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_69_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(_70_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_70_), .C(_66_), .Y(_71_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .C(_71_), .Y(_72_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(_72_), .Y(w_C_15_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .Y(_73_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(i_add1[15]), .Y(_74_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_75_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(_75_), .Y(_76_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_77_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(_78_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_78_), .C(_71_), .Y(_79_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_74_), .C(_79_), .Y(w_C_16_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_74_), .Y(_80_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(_80_), .Y(_81_) );
AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_82_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(_82_), .Y(_83_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_83_), .C(_79_), .Y(_84_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .C(_84_), .Y(_85_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(_85_), .Y(w_C_17_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .Y(_86_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(i_add1[17]), .Y(_87_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_88_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(_88_), .Y(_89_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_90_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(_90_), .Y(_91_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_91_), .C(_84_), .Y(_92_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_87_), .C(_92_), .Y(w_C_18_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_87_), .Y(_93_) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(_93_), .Y(_94_) );
AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_95_) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(_95_), .Y(_96_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_96_), .C(_92_), .Y(_97_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .C(_97_), .Y(_98_) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(_98_), .Y(w_C_19_) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .Y(_99_) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(i_add1[19]), .Y(_100_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_101_) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(_101_), .Y(_102_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_103_) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(_103_), .Y(_104_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_104_), .C(_97_), .Y(_105_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_100_), .C(_105_), .Y(w_C_20_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_100_), .Y(_106_) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(_106_), .Y(_107_) );
AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_108_) );
INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(_108_), .Y(_109_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_109_), .C(_105_), .Y(_110_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .C(_110_), .Y(_111_) );
INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(_111_), .Y(w_C_21_) );
INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .Y(_112_) );
INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(i_add1[21]), .Y(_113_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_114_) );
INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(_114_), .Y(_115_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_116_) );
INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(_116_), .Y(_117_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_117_), .C(_110_), .Y(_118_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_113_), .C(_118_), .Y(w_C_22_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_113_), .Y(_119_) );
INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(_119_), .Y(_120_) );
AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_121_) );
INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(_121_), .Y(_122_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_122_), .C(_118_), .Y(_123_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .C(_123_), .Y(_124_) );
INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(_124_), .Y(w_C_23_) );
INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .Y(_125_) );
INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(i_add1[23]), .Y(_126_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_127_) );
INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(_127_), .Y(_128_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_129_) );
INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(_129_), .Y(_130_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_130_), .C(_123_), .Y(_131_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_126_), .C(_131_), .Y(w_C_24_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_126_), .Y(_132_) );
INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(_132_), .Y(_133_) );
AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_134_) );
INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(_134_), .Y(_135_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_135_), .C(_131_), .Y(_136_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .C(_136_), .Y(_137_) );
INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(_137_), .Y(w_C_25_) );
INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .Y(_138_) );
INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(i_add1[25]), .Y(_139_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_140_) );
INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(_140_), .Y(_141_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_142_) );
INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(_142_), .Y(_143_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_143_), .C(_136_), .Y(_144_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_139_), .C(_144_), .Y(w_C_26_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_139_), .Y(_145_) );
INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(_145_), .Y(_146_) );
AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_147_) );
INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(_147_), .Y(_148_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_148_), .C(_144_), .Y(_149_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .C(_149_), .Y(_150_) );
INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(_150_), .Y(w_C_27_) );
INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .Y(_151_) );
INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(i_add1[27]), .Y(_152_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_153_) );
INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(_153_), .Y(_154_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_155_) );
INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(_156_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_156_), .C(_149_), .Y(_157_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_152_), .C(_157_), .Y(w_C_28_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_152_), .Y(_158_) );
INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(_158_), .Y(_159_) );
AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_160_) );
INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(_160_), .Y(_161_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_159_), .B(_161_), .C(_157_), .Y(_162_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .C(_162_), .Y(_163_) );
INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(_163_), .Y(w_C_29_) );
INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .Y(_164_) );
INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(i_add1[29]), .Y(_165_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_166_) );
INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(_166_), .Y(_167_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_168_) );
INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(_168_), .Y(_169_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_169_), .C(_162_), .Y(_170_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_165_), .C(_170_), .Y(w_C_30_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_165_), .Y(_171_) );
INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(_171_), .Y(_172_) );
AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_173_) );
INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(_173_), .Y(_174_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_174_), .C(_170_), .Y(_175_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .C(_175_), .Y(_176_) );
INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(_176_), .Y(w_C_31_) );
INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .Y(_177_) );
INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(i_add1[31]), .Y(_178_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_179_) );
INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(_179_), .Y(_180_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_181_) );
INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(_181_), .Y(_182_) );
NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_182_), .C(_175_), .Y(_183_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_178_), .C(_183_), .Y(w_C_32_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_178_), .Y(_184_) );
INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(_184_), .Y(_185_) );
AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_186_) );
INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(_186_), .Y(_187_) );
NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_187_), .C(_183_), .Y(_188_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .C(_188_), .Y(_189_) );
INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(_189_), .Y(w_C_33_) );
INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .Y(_190_) );
INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(i_add1[33]), .Y(_191_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_192_) );
INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(_192_), .Y(_193_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_194_) );
INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(_194_), .Y(_195_) );
NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_195_), .C(_188_), .Y(_196_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_191_), .C(_196_), .Y(w_C_34_) );
NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_191_), .Y(_197_) );
INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(_197_), .Y(_198_) );
AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_199_) );
INVX1 INVX1_233 ( .gnd(gnd), .vdd(vdd), .A(_199_), .Y(_200_) );
NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_200_), .C(_196_), .Y(_201_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .C(_201_), .Y(_202_) );
INVX1 INVX1_234 ( .gnd(gnd), .vdd(vdd), .A(_202_), .Y(w_C_35_) );
INVX1 INVX1_235 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .Y(_203_) );
INVX1 INVX1_236 ( .gnd(gnd), .vdd(vdd), .A(i_add1[35]), .Y(_204_) );
NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_205_) );
INVX1 INVX1_237 ( .gnd(gnd), .vdd(vdd), .A(_205_), .Y(_206_) );
NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_207_) );
INVX1 INVX1_238 ( .gnd(gnd), .vdd(vdd), .A(_207_), .Y(_208_) );
NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_208_), .C(_201_), .Y(_209_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_204_), .C(_209_), .Y(w_C_36_) );
NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_204_), .Y(_210_) );
INVX1 INVX1_239 ( .gnd(gnd), .vdd(vdd), .A(_210_), .Y(_211_) );
AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_212_) );
INVX1 INVX1_240 ( .gnd(gnd), .vdd(vdd), .A(_212_), .Y(_213_) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(w_C_62_), .Y(_364__62_) );
BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
