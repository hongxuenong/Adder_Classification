module cla_32bit (i_add1, i_add2, o_result);

input [31:0] i_add1;
input [31:0] i_add2;
output [32:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_176_) );
INVX1 INVX1_1 ( .A(_176_), .Y(w_C_1_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_177_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_0_) );
NOR2X1 NOR2X1_2 ( .A(_177_), .B(_0_), .Y(w_C_2_) );
INVX1 INVX1_2 ( .A(i_add2[2]), .Y(_1_) );
INVX1 INVX1_3 ( .A(i_add1[2]), .Y(_2_) );
NAND2X1 NAND2X1_2 ( .A(_1_), .B(_2_), .Y(_3_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OAI21X1 OAI21X1_1 ( .A(_177_), .B(_0_), .C(_4_), .Y(_5_) );
AND2X2 AND2X2_1 ( .A(_5_), .B(_3_), .Y(w_C_3_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_6_) );
OR2X2 OR2X2_1 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_7_) );
NAND3X1 NAND3X1_1 ( .A(_3_), .B(_7_), .C(_5_), .Y(_8_) );
NAND2X1 NAND2X1_5 ( .A(_6_), .B(_8_), .Y(w_C_4_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_9_) );
INVX1 INVX1_4 ( .A(_9_), .Y(_10_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
NAND3X1 NAND3X1_2 ( .A(_6_), .B(_11_), .C(_8_), .Y(_12_) );
AND2X2 AND2X2_2 ( .A(_12_), .B(_10_), .Y(w_C_5_) );
INVX1 INVX1_5 ( .A(i_add2[5]), .Y(_13_) );
INVX1 INVX1_6 ( .A(i_add1[5]), .Y(_14_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_15_) );
INVX1 INVX1_7 ( .A(_15_), .Y(_16_) );
NAND3X1 NAND3X1_3 ( .A(_10_), .B(_16_), .C(_12_), .Y(_17_) );
OAI21X1 OAI21X1_2 ( .A(_13_), .B(_14_), .C(_17_), .Y(w_C_6_) );
NOR2X1 NOR2X1_5 ( .A(_13_), .B(_14_), .Y(_18_) );
INVX1 INVX1_8 ( .A(_18_), .Y(_19_) );
AND2X2 AND2X2_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_20_) );
INVX1 INVX1_9 ( .A(_20_), .Y(_21_) );
NAND3X1 NAND3X1_4 ( .A(_19_), .B(_21_), .C(_17_), .Y(_22_) );
OAI21X1 OAI21X1_3 ( .A(i_add2[6]), .B(i_add1[6]), .C(_22_), .Y(_23_) );
INVX1 INVX1_10 ( .A(_23_), .Y(w_C_7_) );
INVX1 INVX1_11 ( .A(i_add2[7]), .Y(_24_) );
INVX1 INVX1_12 ( .A(i_add1[7]), .Y(_25_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_26_) );
INVX1 INVX1_13 ( .A(_26_), .Y(_27_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_28_) );
INVX1 INVX1_14 ( .A(_28_), .Y(_29_) );
NAND3X1 NAND3X1_5 ( .A(_27_), .B(_29_), .C(_22_), .Y(_30_) );
OAI21X1 OAI21X1_4 ( .A(_24_), .B(_25_), .C(_30_), .Y(w_C_8_) );
NOR2X1 NOR2X1_8 ( .A(_24_), .B(_25_), .Y(_31_) );
INVX1 INVX1_15 ( .A(_31_), .Y(_32_) );
AND2X2 AND2X2_4 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_33_) );
INVX1 INVX1_16 ( .A(_33_), .Y(_34_) );
NAND3X1 NAND3X1_6 ( .A(_32_), .B(_34_), .C(_30_), .Y(_35_) );
OAI21X1 OAI21X1_5 ( .A(i_add2[8]), .B(i_add1[8]), .C(_35_), .Y(_36_) );
INVX1 INVX1_17 ( .A(_36_), .Y(w_C_9_) );
INVX1 INVX1_18 ( .A(i_add2[9]), .Y(_37_) );
INVX1 INVX1_19 ( .A(i_add1[9]), .Y(_38_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_39_) );
INVX1 INVX1_20 ( .A(_39_), .Y(_40_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_41_) );
INVX1 INVX1_21 ( .A(_41_), .Y(_42_) );
NAND3X1 NAND3X1_7 ( .A(_40_), .B(_42_), .C(_35_), .Y(_43_) );
OAI21X1 OAI21X1_6 ( .A(_37_), .B(_38_), .C(_43_), .Y(w_C_10_) );
NOR2X1 NOR2X1_11 ( .A(_37_), .B(_38_), .Y(_44_) );
INVX1 INVX1_22 ( .A(_44_), .Y(_45_) );
AND2X2 AND2X2_5 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_46_) );
INVX1 INVX1_23 ( .A(_46_), .Y(_47_) );
NAND3X1 NAND3X1_8 ( .A(_45_), .B(_47_), .C(_43_), .Y(_48_) );
OAI21X1 OAI21X1_7 ( .A(i_add2[10]), .B(i_add1[10]), .C(_48_), .Y(_49_) );
INVX1 INVX1_24 ( .A(_49_), .Y(w_C_11_) );
INVX1 INVX1_25 ( .A(i_add2[11]), .Y(_50_) );
INVX1 INVX1_26 ( .A(i_add1[11]), .Y(_51_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_52_) );
INVX1 INVX1_27 ( .A(_52_), .Y(_53_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_54_) );
INVX1 INVX1_28 ( .A(_54_), .Y(_55_) );
NAND3X1 NAND3X1_9 ( .A(_53_), .B(_55_), .C(_48_), .Y(_56_) );
OAI21X1 OAI21X1_8 ( .A(_50_), .B(_51_), .C(_56_), .Y(w_C_12_) );
NOR2X1 NOR2X1_14 ( .A(_50_), .B(_51_), .Y(_57_) );
INVX1 INVX1_29 ( .A(_57_), .Y(_58_) );
AND2X2 AND2X2_6 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_59_) );
INVX1 INVX1_30 ( .A(_59_), .Y(_60_) );
NAND3X1 NAND3X1_10 ( .A(_58_), .B(_60_), .C(_56_), .Y(_61_) );
OAI21X1 OAI21X1_9 ( .A(i_add2[12]), .B(i_add1[12]), .C(_61_), .Y(_62_) );
INVX1 INVX1_31 ( .A(_62_), .Y(w_C_13_) );
INVX1 INVX1_32 ( .A(i_add2[13]), .Y(_63_) );
INVX1 INVX1_33 ( .A(i_add1[13]), .Y(_64_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_65_) );
INVX1 INVX1_34 ( .A(_65_), .Y(_66_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_67_) );
INVX1 INVX1_35 ( .A(_67_), .Y(_68_) );
NAND3X1 NAND3X1_11 ( .A(_66_), .B(_68_), .C(_61_), .Y(_69_) );
OAI21X1 OAI21X1_10 ( .A(_63_), .B(_64_), .C(_69_), .Y(w_C_14_) );
NOR2X1 NOR2X1_17 ( .A(_63_), .B(_64_), .Y(_70_) );
INVX1 INVX1_36 ( .A(_70_), .Y(_71_) );
AND2X2 AND2X2_7 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_72_) );
INVX1 INVX1_37 ( .A(_72_), .Y(_73_) );
NAND3X1 NAND3X1_12 ( .A(_71_), .B(_73_), .C(_69_), .Y(_74_) );
OAI21X1 OAI21X1_11 ( .A(i_add2[14]), .B(i_add1[14]), .C(_74_), .Y(_75_) );
INVX1 INVX1_38 ( .A(_75_), .Y(w_C_15_) );
INVX1 INVX1_39 ( .A(i_add2[15]), .Y(_76_) );
INVX1 INVX1_40 ( .A(i_add1[15]), .Y(_77_) );
NOR2X1 NOR2X1_18 ( .A(_76_), .B(_77_), .Y(_78_) );
INVX1 INVX1_41 ( .A(_78_), .Y(_79_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_80_) );
INVX1 INVX1_42 ( .A(_80_), .Y(_81_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_82_) );
INVX1 INVX1_43 ( .A(_82_), .Y(_83_) );
NAND3X1 NAND3X1_13 ( .A(_81_), .B(_83_), .C(_74_), .Y(_84_) );
AND2X2 AND2X2_8 ( .A(_84_), .B(_79_), .Y(_85_) );
INVX1 INVX1_44 ( .A(_85_), .Y(w_C_16_) );
AND2X2 AND2X2_9 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_86_) );
INVX1 INVX1_45 ( .A(_86_), .Y(_87_) );
NAND3X1 NAND3X1_14 ( .A(_79_), .B(_87_), .C(_84_), .Y(_88_) );
OAI21X1 OAI21X1_12 ( .A(i_add2[16]), .B(i_add1[16]), .C(_88_), .Y(_89_) );
INVX1 INVX1_46 ( .A(_89_), .Y(w_C_17_) );
INVX1 INVX1_47 ( .A(i_add2[17]), .Y(_90_) );
INVX1 INVX1_48 ( .A(i_add1[17]), .Y(_91_) );
NOR2X1 NOR2X1_21 ( .A(_90_), .B(_91_), .Y(_92_) );
INVX1 INVX1_49 ( .A(_92_), .Y(_93_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_94_) );
INVX1 INVX1_50 ( .A(_94_), .Y(_95_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_96_) );
INVX1 INVX1_51 ( .A(_96_), .Y(_97_) );
NAND3X1 NAND3X1_15 ( .A(_95_), .B(_97_), .C(_88_), .Y(_98_) );
AND2X2 AND2X2_10 ( .A(_98_), .B(_93_), .Y(_99_) );
INVX1 INVX1_52 ( .A(_99_), .Y(w_C_18_) );
AND2X2 AND2X2_11 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_100_) );
INVX1 INVX1_53 ( .A(_100_), .Y(_101_) );
NAND3X1 NAND3X1_16 ( .A(_93_), .B(_101_), .C(_98_), .Y(_102_) );
OAI21X1 OAI21X1_13 ( .A(i_add2[18]), .B(i_add1[18]), .C(_102_), .Y(_103_) );
INVX1 INVX1_54 ( .A(_103_), .Y(w_C_19_) );
INVX1 INVX1_55 ( .A(i_add2[19]), .Y(_104_) );
INVX1 INVX1_56 ( .A(i_add1[19]), .Y(_105_) );
NOR2X1 NOR2X1_24 ( .A(_104_), .B(_105_), .Y(_106_) );
INVX1 INVX1_57 ( .A(_106_), .Y(_107_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_108_) );
INVX1 INVX1_58 ( .A(_108_), .Y(_109_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_110_) );
INVX1 INVX1_59 ( .A(_110_), .Y(_111_) );
NAND3X1 NAND3X1_17 ( .A(_109_), .B(_111_), .C(_102_), .Y(_112_) );
AND2X2 AND2X2_12 ( .A(_112_), .B(_107_), .Y(_113_) );
INVX1 INVX1_60 ( .A(_113_), .Y(w_C_20_) );
AND2X2 AND2X2_13 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_114_) );
INVX1 INVX1_61 ( .A(_114_), .Y(_115_) );
NAND3X1 NAND3X1_18 ( .A(_107_), .B(_115_), .C(_112_), .Y(_116_) );
OAI21X1 OAI21X1_14 ( .A(i_add2[20]), .B(i_add1[20]), .C(_116_), .Y(_117_) );
INVX1 INVX1_62 ( .A(_117_), .Y(w_C_21_) );
INVX1 INVX1_63 ( .A(i_add2[21]), .Y(_118_) );
INVX1 INVX1_64 ( .A(i_add1[21]), .Y(_119_) );
NOR2X1 NOR2X1_27 ( .A(_118_), .B(_119_), .Y(_120_) );
INVX1 INVX1_65 ( .A(_120_), .Y(_121_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_122_) );
INVX1 INVX1_66 ( .A(_122_), .Y(_123_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_124_) );
INVX1 INVX1_67 ( .A(_124_), .Y(_125_) );
NAND3X1 NAND3X1_19 ( .A(_123_), .B(_125_), .C(_116_), .Y(_126_) );
AND2X2 AND2X2_14 ( .A(_126_), .B(_121_), .Y(_127_) );
INVX1 INVX1_68 ( .A(_127_), .Y(w_C_22_) );
AND2X2 AND2X2_15 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_128_) );
INVX1 INVX1_69 ( .A(_128_), .Y(_129_) );
NAND3X1 NAND3X1_20 ( .A(_121_), .B(_129_), .C(_126_), .Y(_130_) );
OAI21X1 OAI21X1_15 ( .A(i_add2[22]), .B(i_add1[22]), .C(_130_), .Y(_131_) );
INVX1 INVX1_70 ( .A(_131_), .Y(w_C_23_) );
INVX1 INVX1_71 ( .A(i_add2[23]), .Y(_132_) );
INVX1 INVX1_72 ( .A(i_add1[23]), .Y(_133_) );
NOR2X1 NOR2X1_30 ( .A(_132_), .B(_133_), .Y(_134_) );
INVX1 INVX1_73 ( .A(_134_), .Y(_135_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_136_) );
INVX1 INVX1_74 ( .A(_136_), .Y(_137_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_138_) );
INVX1 INVX1_75 ( .A(_138_), .Y(_139_) );
NAND3X1 NAND3X1_21 ( .A(_137_), .B(_139_), .C(_130_), .Y(_140_) );
AND2X2 AND2X2_16 ( .A(_140_), .B(_135_), .Y(_141_) );
INVX1 INVX1_76 ( .A(_141_), .Y(w_C_24_) );
AND2X2 AND2X2_17 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_142_) );
INVX1 INVX1_77 ( .A(_142_), .Y(_143_) );
NAND3X1 NAND3X1_22 ( .A(_135_), .B(_143_), .C(_140_), .Y(_144_) );
OAI21X1 OAI21X1_16 ( .A(i_add2[24]), .B(i_add1[24]), .C(_144_), .Y(_145_) );
INVX1 INVX1_78 ( .A(_145_), .Y(w_C_25_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_146_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_147_) );
OAI21X1 OAI21X1_17 ( .A(_147_), .B(_145_), .C(_146_), .Y(w_C_26_) );
OR2X2 OR2X2_2 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_148_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_149_) );
INVX1 INVX1_79 ( .A(_149_), .Y(_150_) );
INVX1 INVX1_80 ( .A(_147_), .Y(_151_) );
NAND3X1 NAND3X1_23 ( .A(_150_), .B(_151_), .C(_144_), .Y(_152_) );
NAND2X1 NAND2X1_8 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_153_) );
NAND3X1 NAND3X1_24 ( .A(_146_), .B(_153_), .C(_152_), .Y(_154_) );
AND2X2 AND2X2_18 ( .A(_154_), .B(_148_), .Y(w_C_27_) );
INVX1 INVX1_81 ( .A(i_add2[27]), .Y(_155_) );
INVX1 INVX1_82 ( .A(i_add1[27]), .Y(_156_) );
NAND2X1 NAND2X1_9 ( .A(_155_), .B(_156_), .Y(_157_) );
NAND3X1 NAND3X1_25 ( .A(_148_), .B(_157_), .C(_154_), .Y(_158_) );
OAI21X1 OAI21X1_18 ( .A(_155_), .B(_156_), .C(_158_), .Y(w_C_28_) );
INVX1 INVX1_83 ( .A(i_add2[28]), .Y(_159_) );
INVX1 INVX1_84 ( .A(i_add1[28]), .Y(_160_) );
NAND2X1 NAND2X1_10 ( .A(_159_), .B(_160_), .Y(_161_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_162_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_163_) );
NAND3X1 NAND3X1_26 ( .A(_162_), .B(_163_), .C(_158_), .Y(_164_) );
AND2X2 AND2X2_19 ( .A(_164_), .B(_161_), .Y(w_C_29_) );
INVX1 INVX1_85 ( .A(i_add2[29]), .Y(_165_) );
INVX1 INVX1_86 ( .A(i_add1[29]), .Y(_166_) );
NAND2X1 NAND2X1_13 ( .A(_165_), .B(_166_), .Y(_167_) );
NAND3X1 NAND3X1_27 ( .A(_161_), .B(_167_), .C(_164_), .Y(_168_) );
OAI21X1 OAI21X1_19 ( .A(_165_), .B(_166_), .C(_168_), .Y(w_C_30_) );
OR2X2 OR2X2_3 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_169_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_170_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_171_) );
NAND3X1 NAND3X1_28 ( .A(_170_), .B(_171_), .C(_168_), .Y(_172_) );
AND2X2 AND2X2_20 ( .A(_172_), .B(_169_), .Y(w_C_31_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_173_) );
OR2X2 OR2X2_4 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_174_) );
NAND3X1 NAND3X1_29 ( .A(_169_), .B(_174_), .C(_172_), .Y(_175_) );
NAND2X1 NAND2X1_17 ( .A(_173_), .B(_175_), .Y(w_C_32_) );
BUFX2 BUFX2_1 ( .A(_178__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_178__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_178__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_178__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_178__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_178__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_178__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_178__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_178__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_178__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_178__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_178__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_178__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_178__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_178__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_178__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_178__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_178__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_178__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_178__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_178__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_178__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_178__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_178__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_178__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_178__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_178__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_178__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_178__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_178__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_178__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_178__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(w_C_32_), .Y(o_result[32]) );
INVX1 INVX1_87 ( .A(w_C_4_), .Y(_182_) );
OR2X2 OR2X2_5 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_183_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_184_) );
NAND3X1 NAND3X1_30 ( .A(_182_), .B(_184_), .C(_183_), .Y(_185_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_179_) );
AND2X2 AND2X2_21 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_180_) );
OAI21X1 OAI21X1_20 ( .A(_179_), .B(_180_), .C(w_C_4_), .Y(_181_) );
NAND2X1 NAND2X1_19 ( .A(_181_), .B(_185_), .Y(_178__4_) );
INVX1 INVX1_88 ( .A(w_C_5_), .Y(_189_) );
OR2X2 OR2X2_6 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_190_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_191_) );
NAND3X1 NAND3X1_31 ( .A(_189_), .B(_191_), .C(_190_), .Y(_192_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_186_) );
AND2X2 AND2X2_22 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_187_) );
OAI21X1 OAI21X1_21 ( .A(_186_), .B(_187_), .C(w_C_5_), .Y(_188_) );
NAND2X1 NAND2X1_21 ( .A(_188_), .B(_192_), .Y(_178__5_) );
INVX1 INVX1_89 ( .A(w_C_6_), .Y(_196_) );
OR2X2 OR2X2_7 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_197_) );
NAND2X1 NAND2X1_22 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_198_) );
NAND3X1 NAND3X1_32 ( .A(_196_), .B(_198_), .C(_197_), .Y(_199_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_193_) );
AND2X2 AND2X2_23 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_194_) );
OAI21X1 OAI21X1_22 ( .A(_193_), .B(_194_), .C(w_C_6_), .Y(_195_) );
NAND2X1 NAND2X1_23 ( .A(_195_), .B(_199_), .Y(_178__6_) );
INVX1 INVX1_90 ( .A(w_C_7_), .Y(_203_) );
OR2X2 OR2X2_8 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_204_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_205_) );
NAND3X1 NAND3X1_33 ( .A(_203_), .B(_205_), .C(_204_), .Y(_206_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_200_) );
AND2X2 AND2X2_24 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_201_) );
OAI21X1 OAI21X1_23 ( .A(_200_), .B(_201_), .C(w_C_7_), .Y(_202_) );
NAND2X1 NAND2X1_25 ( .A(_202_), .B(_206_), .Y(_178__7_) );
INVX1 INVX1_91 ( .A(w_C_8_), .Y(_210_) );
OR2X2 OR2X2_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_211_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_212_) );
NAND3X1 NAND3X1_34 ( .A(_210_), .B(_212_), .C(_211_), .Y(_213_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_207_) );
AND2X2 AND2X2_25 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_208_) );
OAI21X1 OAI21X1_24 ( .A(_207_), .B(_208_), .C(w_C_8_), .Y(_209_) );
NAND2X1 NAND2X1_27 ( .A(_209_), .B(_213_), .Y(_178__8_) );
INVX1 INVX1_92 ( .A(w_C_9_), .Y(_217_) );
OR2X2 OR2X2_10 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_218_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_219_) );
NAND3X1 NAND3X1_35 ( .A(_217_), .B(_219_), .C(_218_), .Y(_220_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_214_) );
AND2X2 AND2X2_26 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_215_) );
OAI21X1 OAI21X1_25 ( .A(_214_), .B(_215_), .C(w_C_9_), .Y(_216_) );
NAND2X1 NAND2X1_29 ( .A(_216_), .B(_220_), .Y(_178__9_) );
INVX1 INVX1_93 ( .A(w_C_10_), .Y(_224_) );
OR2X2 OR2X2_11 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_225_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_226_) );
NAND3X1 NAND3X1_36 ( .A(_224_), .B(_226_), .C(_225_), .Y(_227_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_221_) );
AND2X2 AND2X2_27 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_222_) );
OAI21X1 OAI21X1_26 ( .A(_221_), .B(_222_), .C(w_C_10_), .Y(_223_) );
NAND2X1 NAND2X1_31 ( .A(_223_), .B(_227_), .Y(_178__10_) );
INVX1 INVX1_94 ( .A(w_C_11_), .Y(_231_) );
OR2X2 OR2X2_12 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_232_) );
NAND2X1 NAND2X1_32 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_233_) );
NAND3X1 NAND3X1_37 ( .A(_231_), .B(_233_), .C(_232_), .Y(_234_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_228_) );
AND2X2 AND2X2_28 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_229_) );
OAI21X1 OAI21X1_27 ( .A(_228_), .B(_229_), .C(w_C_11_), .Y(_230_) );
NAND2X1 NAND2X1_33 ( .A(_230_), .B(_234_), .Y(_178__11_) );
INVX1 INVX1_95 ( .A(w_C_12_), .Y(_238_) );
OR2X2 OR2X2_13 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_239_) );
NAND2X1 NAND2X1_34 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_240_) );
NAND3X1 NAND3X1_38 ( .A(_238_), .B(_240_), .C(_239_), .Y(_241_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_235_) );
AND2X2 AND2X2_29 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_236_) );
OAI21X1 OAI21X1_28 ( .A(_235_), .B(_236_), .C(w_C_12_), .Y(_237_) );
NAND2X1 NAND2X1_35 ( .A(_237_), .B(_241_), .Y(_178__12_) );
INVX1 INVX1_96 ( .A(w_C_13_), .Y(_245_) );
OR2X2 OR2X2_14 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_246_) );
NAND2X1 NAND2X1_36 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_247_) );
NAND3X1 NAND3X1_39 ( .A(_245_), .B(_247_), .C(_246_), .Y(_248_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_242_) );
AND2X2 AND2X2_30 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_243_) );
OAI21X1 OAI21X1_29 ( .A(_242_), .B(_243_), .C(w_C_13_), .Y(_244_) );
NAND2X1 NAND2X1_37 ( .A(_244_), .B(_248_), .Y(_178__13_) );
INVX1 INVX1_97 ( .A(w_C_14_), .Y(_252_) );
OR2X2 OR2X2_15 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_253_) );
NAND2X1 NAND2X1_38 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_254_) );
NAND3X1 NAND3X1_40 ( .A(_252_), .B(_254_), .C(_253_), .Y(_255_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_249_) );
AND2X2 AND2X2_31 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_250_) );
OAI21X1 OAI21X1_30 ( .A(_249_), .B(_250_), .C(w_C_14_), .Y(_251_) );
NAND2X1 NAND2X1_39 ( .A(_251_), .B(_255_), .Y(_178__14_) );
INVX1 INVX1_98 ( .A(w_C_15_), .Y(_259_) );
OR2X2 OR2X2_16 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_260_) );
NAND2X1 NAND2X1_40 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_261_) );
NAND3X1 NAND3X1_41 ( .A(_259_), .B(_261_), .C(_260_), .Y(_262_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_256_) );
AND2X2 AND2X2_32 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_257_) );
OAI21X1 OAI21X1_31 ( .A(_256_), .B(_257_), .C(w_C_15_), .Y(_258_) );
NAND2X1 NAND2X1_41 ( .A(_258_), .B(_262_), .Y(_178__15_) );
INVX1 INVX1_99 ( .A(w_C_16_), .Y(_266_) );
OR2X2 OR2X2_17 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_267_) );
NAND2X1 NAND2X1_42 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_268_) );
NAND3X1 NAND3X1_42 ( .A(_266_), .B(_268_), .C(_267_), .Y(_269_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_263_) );
AND2X2 AND2X2_33 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_264_) );
OAI21X1 OAI21X1_32 ( .A(_263_), .B(_264_), .C(w_C_16_), .Y(_265_) );
NAND2X1 NAND2X1_43 ( .A(_265_), .B(_269_), .Y(_178__16_) );
INVX1 INVX1_100 ( .A(w_C_17_), .Y(_273_) );
OR2X2 OR2X2_18 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_274_) );
NAND2X1 NAND2X1_44 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_275_) );
NAND3X1 NAND3X1_43 ( .A(_273_), .B(_275_), .C(_274_), .Y(_276_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_270_) );
AND2X2 AND2X2_34 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_271_) );
OAI21X1 OAI21X1_33 ( .A(_270_), .B(_271_), .C(w_C_17_), .Y(_272_) );
NAND2X1 NAND2X1_45 ( .A(_272_), .B(_276_), .Y(_178__17_) );
INVX1 INVX1_101 ( .A(w_C_18_), .Y(_280_) );
OR2X2 OR2X2_19 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_281_) );
NAND2X1 NAND2X1_46 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_282_) );
NAND3X1 NAND3X1_44 ( .A(_280_), .B(_282_), .C(_281_), .Y(_283_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_277_) );
AND2X2 AND2X2_35 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_278_) );
OAI21X1 OAI21X1_34 ( .A(_277_), .B(_278_), .C(w_C_18_), .Y(_279_) );
NAND2X1 NAND2X1_47 ( .A(_279_), .B(_283_), .Y(_178__18_) );
INVX1 INVX1_102 ( .A(w_C_19_), .Y(_287_) );
OR2X2 OR2X2_20 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_288_) );
NAND2X1 NAND2X1_48 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_289_) );
NAND3X1 NAND3X1_45 ( .A(_287_), .B(_289_), .C(_288_), .Y(_290_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_284_) );
AND2X2 AND2X2_36 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_285_) );
OAI21X1 OAI21X1_35 ( .A(_284_), .B(_285_), .C(w_C_19_), .Y(_286_) );
NAND2X1 NAND2X1_49 ( .A(_286_), .B(_290_), .Y(_178__19_) );
INVX1 INVX1_103 ( .A(w_C_20_), .Y(_294_) );
OR2X2 OR2X2_21 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_295_) );
NAND2X1 NAND2X1_50 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_296_) );
NAND3X1 NAND3X1_46 ( .A(_294_), .B(_296_), .C(_295_), .Y(_297_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_291_) );
AND2X2 AND2X2_37 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_292_) );
OAI21X1 OAI21X1_36 ( .A(_291_), .B(_292_), .C(w_C_20_), .Y(_293_) );
NAND2X1 NAND2X1_51 ( .A(_293_), .B(_297_), .Y(_178__20_) );
INVX1 INVX1_104 ( .A(w_C_21_), .Y(_301_) );
OR2X2 OR2X2_22 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_302_) );
NAND2X1 NAND2X1_52 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_303_) );
NAND3X1 NAND3X1_47 ( .A(_301_), .B(_303_), .C(_302_), .Y(_304_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_298_) );
AND2X2 AND2X2_38 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_299_) );
OAI21X1 OAI21X1_37 ( .A(_298_), .B(_299_), .C(w_C_21_), .Y(_300_) );
NAND2X1 NAND2X1_53 ( .A(_300_), .B(_304_), .Y(_178__21_) );
INVX1 INVX1_105 ( .A(w_C_22_), .Y(_308_) );
OR2X2 OR2X2_23 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_309_) );
NAND2X1 NAND2X1_54 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_310_) );
NAND3X1 NAND3X1_48 ( .A(_308_), .B(_310_), .C(_309_), .Y(_311_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_305_) );
AND2X2 AND2X2_39 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_306_) );
OAI21X1 OAI21X1_38 ( .A(_305_), .B(_306_), .C(w_C_22_), .Y(_307_) );
NAND2X1 NAND2X1_55 ( .A(_307_), .B(_311_), .Y(_178__22_) );
INVX1 INVX1_106 ( .A(w_C_23_), .Y(_315_) );
OR2X2 OR2X2_24 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_316_) );
NAND2X1 NAND2X1_56 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_317_) );
NAND3X1 NAND3X1_49 ( .A(_315_), .B(_317_), .C(_316_), .Y(_318_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_312_) );
AND2X2 AND2X2_40 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_313_) );
OAI21X1 OAI21X1_39 ( .A(_312_), .B(_313_), .C(w_C_23_), .Y(_314_) );
NAND2X1 NAND2X1_57 ( .A(_314_), .B(_318_), .Y(_178__23_) );
INVX1 INVX1_107 ( .A(w_C_24_), .Y(_322_) );
OR2X2 OR2X2_25 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_323_) );
NAND2X1 NAND2X1_58 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_324_) );
NAND3X1 NAND3X1_50 ( .A(_322_), .B(_324_), .C(_323_), .Y(_325_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_319_) );
AND2X2 AND2X2_41 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_320_) );
OAI21X1 OAI21X1_40 ( .A(_319_), .B(_320_), .C(w_C_24_), .Y(_321_) );
NAND2X1 NAND2X1_59 ( .A(_321_), .B(_325_), .Y(_178__24_) );
INVX1 INVX1_108 ( .A(w_C_25_), .Y(_329_) );
OR2X2 OR2X2_26 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_330_) );
NAND2X1 NAND2X1_60 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_331_) );
NAND3X1 NAND3X1_51 ( .A(_329_), .B(_331_), .C(_330_), .Y(_332_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_326_) );
AND2X2 AND2X2_42 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_327_) );
OAI21X1 OAI21X1_41 ( .A(_326_), .B(_327_), .C(w_C_25_), .Y(_328_) );
NAND2X1 NAND2X1_61 ( .A(_328_), .B(_332_), .Y(_178__25_) );
INVX1 INVX1_109 ( .A(w_C_26_), .Y(_336_) );
OR2X2 OR2X2_27 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_337_) );
NAND2X1 NAND2X1_62 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_338_) );
NAND3X1 NAND3X1_52 ( .A(_336_), .B(_338_), .C(_337_), .Y(_339_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_333_) );
AND2X2 AND2X2_43 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_334_) );
OAI21X1 OAI21X1_42 ( .A(_333_), .B(_334_), .C(w_C_26_), .Y(_335_) );
NAND2X1 NAND2X1_63 ( .A(_335_), .B(_339_), .Y(_178__26_) );
INVX1 INVX1_110 ( .A(w_C_27_), .Y(_343_) );
OR2X2 OR2X2_28 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_344_) );
NAND2X1 NAND2X1_64 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_345_) );
NAND3X1 NAND3X1_53 ( .A(_343_), .B(_345_), .C(_344_), .Y(_346_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_340_) );
AND2X2 AND2X2_44 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_341_) );
OAI21X1 OAI21X1_43 ( .A(_340_), .B(_341_), .C(w_C_27_), .Y(_342_) );
NAND2X1 NAND2X1_65 ( .A(_342_), .B(_346_), .Y(_178__27_) );
INVX1 INVX1_111 ( .A(w_C_28_), .Y(_350_) );
OR2X2 OR2X2_29 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_351_) );
NAND2X1 NAND2X1_66 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_352_) );
NAND3X1 NAND3X1_54 ( .A(_350_), .B(_352_), .C(_351_), .Y(_353_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_347_) );
AND2X2 AND2X2_45 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_348_) );
OAI21X1 OAI21X1_44 ( .A(_347_), .B(_348_), .C(w_C_28_), .Y(_349_) );
NAND2X1 NAND2X1_67 ( .A(_349_), .B(_353_), .Y(_178__28_) );
INVX1 INVX1_112 ( .A(w_C_29_), .Y(_357_) );
OR2X2 OR2X2_30 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_358_) );
NAND2X1 NAND2X1_68 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_359_) );
NAND3X1 NAND3X1_55 ( .A(_357_), .B(_359_), .C(_358_), .Y(_360_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_354_) );
AND2X2 AND2X2_46 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_355_) );
OAI21X1 OAI21X1_45 ( .A(_354_), .B(_355_), .C(w_C_29_), .Y(_356_) );
NAND2X1 NAND2X1_69 ( .A(_356_), .B(_360_), .Y(_178__29_) );
INVX1 INVX1_113 ( .A(w_C_30_), .Y(_364_) );
OR2X2 OR2X2_31 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_365_) );
NAND2X1 NAND2X1_70 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_366_) );
NAND3X1 NAND3X1_56 ( .A(_364_), .B(_366_), .C(_365_), .Y(_367_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_361_) );
AND2X2 AND2X2_47 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_362_) );
OAI21X1 OAI21X1_46 ( .A(_361_), .B(_362_), .C(w_C_30_), .Y(_363_) );
NAND2X1 NAND2X1_71 ( .A(_363_), .B(_367_), .Y(_178__30_) );
INVX1 INVX1_114 ( .A(w_C_31_), .Y(_371_) );
OR2X2 OR2X2_32 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_372_) );
NAND2X1 NAND2X1_72 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_373_) );
NAND3X1 NAND3X1_57 ( .A(_371_), .B(_373_), .C(_372_), .Y(_374_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_368_) );
AND2X2 AND2X2_48 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_369_) );
OAI21X1 OAI21X1_47 ( .A(_368_), .B(_369_), .C(w_C_31_), .Y(_370_) );
NAND2X1 NAND2X1_73 ( .A(_370_), .B(_374_), .Y(_178__31_) );
INVX1 INVX1_115 ( .A(gnd), .Y(_378_) );
OR2X2 OR2X2_33 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_379_) );
NAND2X1 NAND2X1_74 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_380_) );
NAND3X1 NAND3X1_58 ( .A(_378_), .B(_380_), .C(_379_), .Y(_381_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_375_) );
AND2X2 AND2X2_49 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_376_) );
OAI21X1 OAI21X1_48 ( .A(_375_), .B(_376_), .C(gnd), .Y(_377_) );
NAND2X1 NAND2X1_75 ( .A(_377_), .B(_381_), .Y(_178__0_) );
INVX1 INVX1_116 ( .A(w_C_1_), .Y(_385_) );
OR2X2 OR2X2_34 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_386_) );
NAND2X1 NAND2X1_76 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_387_) );
NAND3X1 NAND3X1_59 ( .A(_385_), .B(_387_), .C(_386_), .Y(_388_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_382_) );
AND2X2 AND2X2_50 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_383_) );
OAI21X1 OAI21X1_49 ( .A(_382_), .B(_383_), .C(w_C_1_), .Y(_384_) );
NAND2X1 NAND2X1_77 ( .A(_384_), .B(_388_), .Y(_178__1_) );
INVX1 INVX1_117 ( .A(w_C_2_), .Y(_392_) );
OR2X2 OR2X2_35 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_393_) );
NAND2X1 NAND2X1_78 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_394_) );
NAND3X1 NAND3X1_60 ( .A(_392_), .B(_394_), .C(_393_), .Y(_395_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_389_) );
AND2X2 AND2X2_51 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_390_) );
OAI21X1 OAI21X1_50 ( .A(_389_), .B(_390_), .C(w_C_2_), .Y(_391_) );
NAND2X1 NAND2X1_79 ( .A(_391_), .B(_395_), .Y(_178__2_) );
INVX1 INVX1_118 ( .A(w_C_3_), .Y(_399_) );
OR2X2 OR2X2_36 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_400_) );
NAND2X1 NAND2X1_80 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_401_) );
NAND3X1 NAND3X1_61 ( .A(_399_), .B(_401_), .C(_400_), .Y(_402_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_396_) );
AND2X2 AND2X2_52 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_397_) );
OAI21X1 OAI21X1_51 ( .A(_396_), .B(_397_), .C(w_C_3_), .Y(_398_) );
NAND2X1 NAND2X1_81 ( .A(_398_), .B(_402_), .Y(_178__3_) );
BUFX2 BUFX2_34 ( .A(w_C_32_), .Y(_178__32_) );
BUFX2 BUFX2_35 ( .A(gnd), .Y(w_C_0_) );
endmodule
