module CSkipA_45bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [44:0] i_add_term1;
input [44:0] i_add_term2;
output [44:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

NAND2X1 NAND2X1_1 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_383_) );
NAND3X1 NAND3X1_1 ( .A(_381_), .B(_383_), .C(_382_), .Y(_384_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_378_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_379_) );
OAI21X1 OAI21X1_1 ( .A(_378_), .B(_379_), .C(w_cout_6_), .Y(_380_) );
NAND2X1 NAND2X1_2 ( .A(_380_), .B(_384_), .Y(_0__24_) );
OAI21X1 OAI21X1_2 ( .A(_381_), .B(_378_), .C(_383_), .Y(_20__1_) );
INVX1 INVX1_1 ( .A(_20__1_), .Y(_388_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_389_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_390_) );
NAND3X1 NAND3X1_2 ( .A(_388_), .B(_390_), .C(_389_), .Y(_391_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_385_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_386_) );
OAI21X1 OAI21X1_3 ( .A(_385_), .B(_386_), .C(_20__1_), .Y(_387_) );
NAND2X1 NAND2X1_4 ( .A(_387_), .B(_391_), .Y(_0__25_) );
OAI21X1 OAI21X1_4 ( .A(_388_), .B(_385_), .C(_390_), .Y(_20__2_) );
INVX1 INVX1_2 ( .A(_20__2_), .Y(_395_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_396_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_397_) );
NAND3X1 NAND3X1_3 ( .A(_395_), .B(_397_), .C(_396_), .Y(_398_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_392_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_393_) );
OAI21X1 OAI21X1_5 ( .A(_392_), .B(_393_), .C(_20__2_), .Y(_394_) );
NAND2X1 NAND2X1_6 ( .A(_394_), .B(_398_), .Y(_0__26_) );
OAI21X1 OAI21X1_6 ( .A(_395_), .B(_392_), .C(_397_), .Y(_20__3_) );
INVX1 INVX1_3 ( .A(_20__3_), .Y(_402_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_403_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_404_) );
NAND3X1 NAND3X1_4 ( .A(_402_), .B(_404_), .C(_403_), .Y(_405_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_399_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_400_) );
OAI21X1 OAI21X1_7 ( .A(_399_), .B(_400_), .C(_20__3_), .Y(_401_) );
NAND2X1 NAND2X1_8 ( .A(_401_), .B(_405_), .Y(_0__27_) );
OAI21X1 OAI21X1_8 ( .A(_402_), .B(_399_), .C(_404_), .Y(_19_) );
INVX1 INVX1_4 ( .A(w_cout_7_), .Y(_409_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_410_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_411_) );
NAND3X1 NAND3X1_5 ( .A(_409_), .B(_411_), .C(_410_), .Y(_412_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_406_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_407_) );
OAI21X1 OAI21X1_9 ( .A(_406_), .B(_407_), .C(w_cout_7_), .Y(_408_) );
NAND2X1 NAND2X1_10 ( .A(_408_), .B(_412_), .Y(_0__28_) );
OAI21X1 OAI21X1_10 ( .A(_409_), .B(_406_), .C(_411_), .Y(_23__1_) );
INVX1 INVX1_5 ( .A(_23__1_), .Y(_416_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_417_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_418_) );
NAND3X1 NAND3X1_6 ( .A(_416_), .B(_418_), .C(_417_), .Y(_419_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_413_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_414_) );
OAI21X1 OAI21X1_11 ( .A(_413_), .B(_414_), .C(_23__1_), .Y(_415_) );
NAND2X1 NAND2X1_12 ( .A(_415_), .B(_419_), .Y(_0__29_) );
OAI21X1 OAI21X1_12 ( .A(_416_), .B(_413_), .C(_418_), .Y(_23__2_) );
INVX1 INVX1_6 ( .A(_23__2_), .Y(_423_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_424_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_425_) );
NAND3X1 NAND3X1_7 ( .A(_423_), .B(_425_), .C(_424_), .Y(_426_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_420_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_421_) );
OAI21X1 OAI21X1_13 ( .A(_420_), .B(_421_), .C(_23__2_), .Y(_422_) );
NAND2X1 NAND2X1_14 ( .A(_422_), .B(_426_), .Y(_0__30_) );
OAI21X1 OAI21X1_14 ( .A(_423_), .B(_420_), .C(_425_), .Y(_23__3_) );
INVX1 INVX1_7 ( .A(_23__3_), .Y(_430_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_431_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_432_) );
NAND3X1 NAND3X1_8 ( .A(_430_), .B(_432_), .C(_431_), .Y(_433_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_427_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_428_) );
OAI21X1 OAI21X1_15 ( .A(_427_), .B(_428_), .C(_23__3_), .Y(_429_) );
NAND2X1 NAND2X1_16 ( .A(_429_), .B(_433_), .Y(_0__31_) );
OAI21X1 OAI21X1_16 ( .A(_430_), .B(_427_), .C(_432_), .Y(_22_) );
INVX1 INVX1_8 ( .A(w_cout_8_), .Y(_437_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_438_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_439_) );
NAND3X1 NAND3X1_9 ( .A(_437_), .B(_439_), .C(_438_), .Y(_440_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_434_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_435_) );
OAI21X1 OAI21X1_17 ( .A(_434_), .B(_435_), .C(w_cout_8_), .Y(_436_) );
NAND2X1 NAND2X1_18 ( .A(_436_), .B(_440_), .Y(_0__32_) );
OAI21X1 OAI21X1_18 ( .A(_437_), .B(_434_), .C(_439_), .Y(_26__1_) );
INVX1 INVX1_9 ( .A(_26__1_), .Y(_444_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_445_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_446_) );
NAND3X1 NAND3X1_10 ( .A(_444_), .B(_446_), .C(_445_), .Y(_447_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_441_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_442_) );
OAI21X1 OAI21X1_19 ( .A(_441_), .B(_442_), .C(_26__1_), .Y(_443_) );
NAND2X1 NAND2X1_20 ( .A(_443_), .B(_447_), .Y(_0__33_) );
OAI21X1 OAI21X1_20 ( .A(_444_), .B(_441_), .C(_446_), .Y(_26__2_) );
INVX1 INVX1_10 ( .A(_26__2_), .Y(_451_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_452_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_453_) );
NAND3X1 NAND3X1_11 ( .A(_451_), .B(_453_), .C(_452_), .Y(_454_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_448_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_449_) );
OAI21X1 OAI21X1_21 ( .A(_448_), .B(_449_), .C(_26__2_), .Y(_450_) );
NAND2X1 NAND2X1_22 ( .A(_450_), .B(_454_), .Y(_0__34_) );
OAI21X1 OAI21X1_22 ( .A(_451_), .B(_448_), .C(_453_), .Y(_26__3_) );
INVX1 INVX1_11 ( .A(_26__3_), .Y(_458_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_459_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_460_) );
NAND3X1 NAND3X1_12 ( .A(_458_), .B(_460_), .C(_459_), .Y(_461_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_455_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_456_) );
OAI21X1 OAI21X1_23 ( .A(_455_), .B(_456_), .C(_26__3_), .Y(_457_) );
NAND2X1 NAND2X1_24 ( .A(_457_), .B(_461_), .Y(_0__35_) );
OAI21X1 OAI21X1_24 ( .A(_458_), .B(_455_), .C(_460_), .Y(_25_) );
INVX1 INVX1_12 ( .A(w_cout_9_), .Y(_465_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_466_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_467_) );
NAND3X1 NAND3X1_13 ( .A(_465_), .B(_467_), .C(_466_), .Y(_468_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_462_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_463_) );
OAI21X1 OAI21X1_25 ( .A(_462_), .B(_463_), .C(w_cout_9_), .Y(_464_) );
NAND2X1 NAND2X1_26 ( .A(_464_), .B(_468_), .Y(_0__36_) );
OAI21X1 OAI21X1_26 ( .A(_465_), .B(_462_), .C(_467_), .Y(_29__1_) );
INVX1 INVX1_13 ( .A(_29__1_), .Y(_472_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_473_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_474_) );
NAND3X1 NAND3X1_14 ( .A(_472_), .B(_474_), .C(_473_), .Y(_475_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_469_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_470_) );
OAI21X1 OAI21X1_27 ( .A(_469_), .B(_470_), .C(_29__1_), .Y(_471_) );
NAND2X1 NAND2X1_28 ( .A(_471_), .B(_475_), .Y(_0__37_) );
OAI21X1 OAI21X1_28 ( .A(_472_), .B(_469_), .C(_474_), .Y(_29__2_) );
INVX1 INVX1_14 ( .A(_29__2_), .Y(_479_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_480_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_481_) );
NAND3X1 NAND3X1_15 ( .A(_479_), .B(_481_), .C(_480_), .Y(_482_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_476_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_477_) );
OAI21X1 OAI21X1_29 ( .A(_476_), .B(_477_), .C(_29__2_), .Y(_478_) );
NAND2X1 NAND2X1_30 ( .A(_478_), .B(_482_), .Y(_0__38_) );
OAI21X1 OAI21X1_30 ( .A(_479_), .B(_476_), .C(_481_), .Y(_29__3_) );
INVX1 INVX1_15 ( .A(_29__3_), .Y(_486_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_487_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_488_) );
NAND3X1 NAND3X1_16 ( .A(_486_), .B(_488_), .C(_487_), .Y(_489_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_483_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_484_) );
OAI21X1 OAI21X1_31 ( .A(_483_), .B(_484_), .C(_29__3_), .Y(_485_) );
NAND2X1 NAND2X1_32 ( .A(_485_), .B(_489_), .Y(_0__39_) );
OAI21X1 OAI21X1_32 ( .A(_486_), .B(_483_), .C(_488_), .Y(_28_) );
INVX1 INVX1_16 ( .A(w_cout_10_), .Y(_493_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_494_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_495_) );
NAND3X1 NAND3X1_17 ( .A(_493_), .B(_495_), .C(_494_), .Y(_496_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_490_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_491_) );
OAI21X1 OAI21X1_33 ( .A(_490_), .B(_491_), .C(w_cout_10_), .Y(_492_) );
NAND2X1 NAND2X1_34 ( .A(_492_), .B(_496_), .Y(_0__40_) );
OAI21X1 OAI21X1_34 ( .A(_493_), .B(_490_), .C(_495_), .Y(_32__1_) );
INVX1 INVX1_17 ( .A(_32__1_), .Y(_500_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_501_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_502_) );
NAND3X1 NAND3X1_18 ( .A(_500_), .B(_502_), .C(_501_), .Y(_503_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_497_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_498_) );
OAI21X1 OAI21X1_35 ( .A(_497_), .B(_498_), .C(_32__1_), .Y(_499_) );
NAND2X1 NAND2X1_36 ( .A(_499_), .B(_503_), .Y(_0__41_) );
OAI21X1 OAI21X1_36 ( .A(_500_), .B(_497_), .C(_502_), .Y(_32__2_) );
INVX1 INVX1_18 ( .A(_32__2_), .Y(_507_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_508_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_509_) );
NAND3X1 NAND3X1_19 ( .A(_507_), .B(_509_), .C(_508_), .Y(_510_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_504_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_505_) );
OAI21X1 OAI21X1_37 ( .A(_504_), .B(_505_), .C(_32__2_), .Y(_506_) );
NAND2X1 NAND2X1_38 ( .A(_506_), .B(_510_), .Y(_0__42_) );
OAI21X1 OAI21X1_38 ( .A(_507_), .B(_504_), .C(_509_), .Y(_32__3_) );
INVX1 INVX1_19 ( .A(_32__3_), .Y(_514_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_515_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_516_) );
NAND3X1 NAND3X1_20 ( .A(_514_), .B(_516_), .C(_515_), .Y(_517_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_511_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_512_) );
OAI21X1 OAI21X1_39 ( .A(_511_), .B(_512_), .C(_32__3_), .Y(_513_) );
NAND2X1 NAND2X1_40 ( .A(_513_), .B(_517_), .Y(_0__43_) );
OAI21X1 OAI21X1_40 ( .A(_514_), .B(_511_), .C(_516_), .Y(_31_) );
INVX1 INVX1_20 ( .A(cskip1_inst_cin), .Y(_521_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_522_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_523_) );
NAND3X1 NAND3X1_21 ( .A(_521_), .B(_523_), .C(_522_), .Y(_524_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_518_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_519_) );
OAI21X1 OAI21X1_41 ( .A(_518_), .B(_519_), .C(cskip1_inst_cin), .Y(_520_) );
NAND2X1 NAND2X1_42 ( .A(_520_), .B(_524_), .Y(cskip1_inst_sum) );
OAI21X1 OAI21X1_42 ( .A(_521_), .B(_518_), .C(_523_), .Y(cskip1_inst_rca0_w_CARRY_1_) );
INVX1 INVX1_21 ( .A(cskip1_inst_rca0_w_CARRY_1_), .Y(_526_) );
NAND2X1 NAND2X1_43 ( .A(gnd), .B(gnd), .Y(_527_) );
NOR2X1 NOR2X1_22 ( .A(gnd), .B(gnd), .Y(_525_) );
OAI21X1 OAI21X1_43 ( .A(_526_), .B(_525_), .C(_527_), .Y(cskip1_inst_rca0_w_CARRY_2_) );
INVX1 INVX1_22 ( .A(cskip1_inst_rca0_w_CARRY_2_), .Y(_529_) );
NAND2X1 NAND2X1_44 ( .A(gnd), .B(gnd), .Y(_530_) );
NOR2X1 NOR2X1_23 ( .A(gnd), .B(gnd), .Y(_528_) );
OAI21X1 OAI21X1_44 ( .A(_529_), .B(_528_), .C(_530_), .Y(cskip1_inst_rca0_w_CARRY_3_) );
INVX1 INVX1_23 ( .A(cskip1_inst_rca0_w_CARRY_3_), .Y(_532_) );
NAND2X1 NAND2X1_45 ( .A(gnd), .B(gnd), .Y(_533_) );
NOR2X1 NOR2X1_24 ( .A(gnd), .B(gnd), .Y(_531_) );
OAI21X1 OAI21X1_45 ( .A(_532_), .B(_531_), .C(_533_), .Y(cskip1_inst_cout0) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_534_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_535_) );
NOR2X1 NOR2X1_26 ( .A(_534_), .B(_535_), .Y(cskip1_inst_skip0_P) );
INVX1 INVX1_24 ( .A(cskip1_inst_cout0), .Y(_536_) );
NAND2X1 NAND2X1_46 ( .A(gnd), .B(cskip1_inst_skip0_P), .Y(_537_) );
OAI21X1 OAI21X1_46 ( .A(cskip1_inst_skip0_P), .B(_536_), .C(_537_), .Y(w_cout_12_) );
BUFX2 BUFX2_1 ( .A(w_cout_12_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(cskip1_inst_sum), .Y(sum[44]) );
INVX1 INVX1_25 ( .A(i_add_term1[0]), .Y(_34_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[0]), .B(_34_), .Y(_35_) );
INVX1 INVX1_26 ( .A(i_add_term2[0]), .Y(_36_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term1[0]), .B(_36_), .Y(_37_) );
INVX1 INVX1_27 ( .A(i_add_term1[1]), .Y(_38_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[1]), .B(_38_), .Y(_39_) );
INVX1 INVX1_28 ( .A(i_add_term2[1]), .Y(_40_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term1[1]), .B(_40_), .Y(_41_) );
OAI22X1 OAI22X1_1 ( .A(_35_), .B(_37_), .C(_39_), .D(_41_), .Y(_42_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_43_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_44_) );
NOR2X1 NOR2X1_32 ( .A(_43_), .B(_44_), .Y(_45_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_46_) );
NAND2X1 NAND2X1_47 ( .A(_45_), .B(_46_), .Y(_47_) );
NOR2X1 NOR2X1_33 ( .A(_42_), .B(_47_), .Y(_3_) );
INVX1 INVX1_29 ( .A(_1_), .Y(_48_) );
NAND2X1 NAND2X1_48 ( .A(gnd), .B(_3_), .Y(_49_) );
OAI21X1 OAI21X1_47 ( .A(_3_), .B(_48_), .C(_49_), .Y(w_cout_1_) );
INVX1 INVX1_30 ( .A(i_add_term1[4]), .Y(_50_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[4]), .B(_50_), .Y(_51_) );
INVX1 INVX1_31 ( .A(i_add_term2[4]), .Y(_52_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term1[4]), .B(_52_), .Y(_53_) );
INVX1 INVX1_32 ( .A(i_add_term1[5]), .Y(_54_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[5]), .B(_54_), .Y(_55_) );
INVX1 INVX1_33 ( .A(i_add_term2[5]), .Y(_56_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term1[5]), .B(_56_), .Y(_57_) );
OAI22X1 OAI22X1_2 ( .A(_51_), .B(_53_), .C(_55_), .D(_57_), .Y(_58_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_59_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_60_) );
NOR2X1 NOR2X1_39 ( .A(_59_), .B(_60_), .Y(_61_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_62_) );
NAND2X1 NAND2X1_49 ( .A(_61_), .B(_62_), .Y(_63_) );
NOR2X1 NOR2X1_40 ( .A(_58_), .B(_63_), .Y(_6_) );
INVX1 INVX1_34 ( .A(_4_), .Y(_64_) );
NAND2X1 NAND2X1_50 ( .A(gnd), .B(_6_), .Y(_65_) );
OAI21X1 OAI21X1_48 ( .A(_6_), .B(_64_), .C(_65_), .Y(w_cout_2_) );
INVX1 INVX1_35 ( .A(i_add_term1[8]), .Y(_66_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[8]), .B(_66_), .Y(_67_) );
INVX1 INVX1_36 ( .A(i_add_term2[8]), .Y(_68_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term1[8]), .B(_68_), .Y(_69_) );
INVX1 INVX1_37 ( .A(i_add_term1[9]), .Y(_70_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[9]), .B(_70_), .Y(_71_) );
INVX1 INVX1_38 ( .A(i_add_term2[9]), .Y(_72_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term1[9]), .B(_72_), .Y(_73_) );
OAI22X1 OAI22X1_3 ( .A(_67_), .B(_69_), .C(_71_), .D(_73_), .Y(_74_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_75_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_76_) );
NOR2X1 NOR2X1_46 ( .A(_75_), .B(_76_), .Y(_77_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_78_) );
NAND2X1 NAND2X1_51 ( .A(_77_), .B(_78_), .Y(_79_) );
NOR2X1 NOR2X1_47 ( .A(_74_), .B(_79_), .Y(_9_) );
INVX1 INVX1_39 ( .A(_7_), .Y(_80_) );
NAND2X1 NAND2X1_52 ( .A(gnd), .B(_9_), .Y(_81_) );
OAI21X1 OAI21X1_49 ( .A(_9_), .B(_80_), .C(_81_), .Y(w_cout_3_) );
INVX1 INVX1_40 ( .A(i_add_term1[12]), .Y(_82_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[12]), .B(_82_), .Y(_83_) );
INVX1 INVX1_41 ( .A(i_add_term2[12]), .Y(_84_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term1[12]), .B(_84_), .Y(_85_) );
INVX1 INVX1_42 ( .A(i_add_term1[13]), .Y(_86_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[13]), .B(_86_), .Y(_87_) );
INVX1 INVX1_43 ( .A(i_add_term2[13]), .Y(_88_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term1[13]), .B(_88_), .Y(_89_) );
OAI22X1 OAI22X1_4 ( .A(_83_), .B(_85_), .C(_87_), .D(_89_), .Y(_90_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_91_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_92_) );
NOR2X1 NOR2X1_53 ( .A(_91_), .B(_92_), .Y(_93_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_94_) );
NAND2X1 NAND2X1_53 ( .A(_93_), .B(_94_), .Y(_95_) );
NOR2X1 NOR2X1_54 ( .A(_90_), .B(_95_), .Y(_12_) );
INVX1 INVX1_44 ( .A(_10_), .Y(_96_) );
NAND2X1 NAND2X1_54 ( .A(gnd), .B(_12_), .Y(_97_) );
OAI21X1 OAI21X1_50 ( .A(_12_), .B(_96_), .C(_97_), .Y(w_cout_4_) );
INVX1 INVX1_45 ( .A(i_add_term1[16]), .Y(_98_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[16]), .B(_98_), .Y(_99_) );
INVX1 INVX1_46 ( .A(i_add_term2[16]), .Y(_100_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term1[16]), .B(_100_), .Y(_101_) );
INVX1 INVX1_47 ( .A(i_add_term1[17]), .Y(_102_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[17]), .B(_102_), .Y(_103_) );
INVX1 INVX1_48 ( .A(i_add_term2[17]), .Y(_104_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term1[17]), .B(_104_), .Y(_105_) );
OAI22X1 OAI22X1_5 ( .A(_99_), .B(_101_), .C(_103_), .D(_105_), .Y(_106_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_107_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_108_) );
NOR2X1 NOR2X1_60 ( .A(_107_), .B(_108_), .Y(_109_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_110_) );
NAND2X1 NAND2X1_55 ( .A(_109_), .B(_110_), .Y(_111_) );
NOR2X1 NOR2X1_61 ( .A(_106_), .B(_111_), .Y(_15_) );
INVX1 INVX1_49 ( .A(_13_), .Y(_112_) );
NAND2X1 NAND2X1_56 ( .A(gnd), .B(_15_), .Y(_113_) );
OAI21X1 OAI21X1_51 ( .A(_15_), .B(_112_), .C(_113_), .Y(w_cout_5_) );
INVX1 INVX1_50 ( .A(i_add_term1[20]), .Y(_114_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[20]), .B(_114_), .Y(_115_) );
INVX1 INVX1_51 ( .A(i_add_term2[20]), .Y(_116_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term1[20]), .B(_116_), .Y(_117_) );
INVX1 INVX1_52 ( .A(i_add_term1[21]), .Y(_118_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[21]), .B(_118_), .Y(_119_) );
INVX1 INVX1_53 ( .A(i_add_term2[21]), .Y(_120_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term1[21]), .B(_120_), .Y(_121_) );
OAI22X1 OAI22X1_6 ( .A(_115_), .B(_117_), .C(_119_), .D(_121_), .Y(_122_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_123_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_124_) );
NOR2X1 NOR2X1_67 ( .A(_123_), .B(_124_), .Y(_125_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_126_) );
NAND2X1 NAND2X1_57 ( .A(_125_), .B(_126_), .Y(_127_) );
NOR2X1 NOR2X1_68 ( .A(_122_), .B(_127_), .Y(_18_) );
INVX1 INVX1_54 ( .A(_16_), .Y(_128_) );
NAND2X1 NAND2X1_58 ( .A(gnd), .B(_18_), .Y(_129_) );
OAI21X1 OAI21X1_52 ( .A(_18_), .B(_128_), .C(_129_), .Y(w_cout_6_) );
INVX1 INVX1_55 ( .A(i_add_term1[24]), .Y(_130_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[24]), .B(_130_), .Y(_131_) );
INVX1 INVX1_56 ( .A(i_add_term2[24]), .Y(_132_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term1[24]), .B(_132_), .Y(_133_) );
INVX1 INVX1_57 ( .A(i_add_term1[25]), .Y(_134_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[25]), .B(_134_), .Y(_135_) );
INVX1 INVX1_58 ( .A(i_add_term2[25]), .Y(_136_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term1[25]), .B(_136_), .Y(_137_) );
OAI22X1 OAI22X1_7 ( .A(_131_), .B(_133_), .C(_135_), .D(_137_), .Y(_138_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_139_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_140_) );
NOR2X1 NOR2X1_74 ( .A(_139_), .B(_140_), .Y(_141_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_142_) );
NAND2X1 NAND2X1_59 ( .A(_141_), .B(_142_), .Y(_143_) );
NOR2X1 NOR2X1_75 ( .A(_138_), .B(_143_), .Y(_21_) );
INVX1 INVX1_59 ( .A(_19_), .Y(_144_) );
NAND2X1 NAND2X1_60 ( .A(gnd), .B(_21_), .Y(_145_) );
OAI21X1 OAI21X1_53 ( .A(_21_), .B(_144_), .C(_145_), .Y(w_cout_7_) );
INVX1 INVX1_60 ( .A(i_add_term1[28]), .Y(_146_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[28]), .B(_146_), .Y(_147_) );
INVX1 INVX1_61 ( .A(i_add_term2[28]), .Y(_148_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term1[28]), .B(_148_), .Y(_149_) );
INVX1 INVX1_62 ( .A(i_add_term1[29]), .Y(_150_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[29]), .B(_150_), .Y(_151_) );
INVX1 INVX1_63 ( .A(i_add_term2[29]), .Y(_152_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term1[29]), .B(_152_), .Y(_153_) );
OAI22X1 OAI22X1_8 ( .A(_147_), .B(_149_), .C(_151_), .D(_153_), .Y(_154_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_155_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_156_) );
NOR2X1 NOR2X1_81 ( .A(_155_), .B(_156_), .Y(_157_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_158_) );
NAND2X1 NAND2X1_61 ( .A(_157_), .B(_158_), .Y(_159_) );
NOR2X1 NOR2X1_82 ( .A(_154_), .B(_159_), .Y(_24_) );
INVX1 INVX1_64 ( .A(_22_), .Y(_160_) );
NAND2X1 NAND2X1_62 ( .A(gnd), .B(_24_), .Y(_161_) );
OAI21X1 OAI21X1_54 ( .A(_24_), .B(_160_), .C(_161_), .Y(w_cout_8_) );
INVX1 INVX1_65 ( .A(i_add_term1[32]), .Y(_162_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[32]), .B(_162_), .Y(_163_) );
INVX1 INVX1_66 ( .A(i_add_term2[32]), .Y(_164_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term1[32]), .B(_164_), .Y(_165_) );
INVX1 INVX1_67 ( .A(i_add_term1[33]), .Y(_166_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[33]), .B(_166_), .Y(_167_) );
INVX1 INVX1_68 ( .A(i_add_term2[33]), .Y(_168_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term1[33]), .B(_168_), .Y(_169_) );
OAI22X1 OAI22X1_9 ( .A(_163_), .B(_165_), .C(_167_), .D(_169_), .Y(_170_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_171_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_172_) );
NOR2X1 NOR2X1_88 ( .A(_171_), .B(_172_), .Y(_173_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_174_) );
NAND2X1 NAND2X1_63 ( .A(_173_), .B(_174_), .Y(_175_) );
NOR2X1 NOR2X1_89 ( .A(_170_), .B(_175_), .Y(_27_) );
INVX1 INVX1_69 ( .A(_25_), .Y(_176_) );
NAND2X1 NAND2X1_64 ( .A(gnd), .B(_27_), .Y(_177_) );
OAI21X1 OAI21X1_55 ( .A(_27_), .B(_176_), .C(_177_), .Y(w_cout_9_) );
INVX1 INVX1_70 ( .A(i_add_term1[36]), .Y(_178_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[36]), .B(_178_), .Y(_179_) );
INVX1 INVX1_71 ( .A(i_add_term2[36]), .Y(_180_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term1[36]), .B(_180_), .Y(_181_) );
INVX1 INVX1_72 ( .A(i_add_term1[37]), .Y(_182_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[37]), .B(_182_), .Y(_183_) );
INVX1 INVX1_73 ( .A(i_add_term2[37]), .Y(_184_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term1[37]), .B(_184_), .Y(_185_) );
OAI22X1 OAI22X1_10 ( .A(_179_), .B(_181_), .C(_183_), .D(_185_), .Y(_186_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_187_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_188_) );
NOR2X1 NOR2X1_95 ( .A(_187_), .B(_188_), .Y(_189_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_190_) );
NAND2X1 NAND2X1_65 ( .A(_189_), .B(_190_), .Y(_191_) );
NOR2X1 NOR2X1_96 ( .A(_186_), .B(_191_), .Y(_30_) );
INVX1 INVX1_74 ( .A(_28_), .Y(_192_) );
NAND2X1 NAND2X1_66 ( .A(gnd), .B(_30_), .Y(_193_) );
OAI21X1 OAI21X1_56 ( .A(_30_), .B(_192_), .C(_193_), .Y(w_cout_10_) );
INVX1 INVX1_75 ( .A(i_add_term1[40]), .Y(_194_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[40]), .B(_194_), .Y(_195_) );
INVX1 INVX1_76 ( .A(i_add_term2[40]), .Y(_196_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term1[40]), .B(_196_), .Y(_197_) );
INVX1 INVX1_77 ( .A(i_add_term1[41]), .Y(_198_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[41]), .B(_198_), .Y(_199_) );
INVX1 INVX1_78 ( .A(i_add_term2[41]), .Y(_200_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term1[41]), .B(_200_), .Y(_201_) );
OAI22X1 OAI22X1_11 ( .A(_195_), .B(_197_), .C(_199_), .D(_201_), .Y(_202_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_203_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_204_) );
NOR2X1 NOR2X1_102 ( .A(_203_), .B(_204_), .Y(_205_) );
XOR2X1 XOR2X1_11 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_206_) );
NAND2X1 NAND2X1_67 ( .A(_205_), .B(_206_), .Y(_207_) );
NOR2X1 NOR2X1_103 ( .A(_202_), .B(_207_), .Y(_33_) );
INVX1 INVX1_79 ( .A(_31_), .Y(_208_) );
NAND2X1 NAND2X1_68 ( .A(gnd), .B(_33_), .Y(_209_) );
OAI21X1 OAI21X1_57 ( .A(_33_), .B(_208_), .C(_209_), .Y(cskip1_inst_cin) );
INVX1 INVX1_80 ( .A(gnd), .Y(_213_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_214_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_215_) );
NAND3X1 NAND3X1_22 ( .A(_213_), .B(_215_), .C(_214_), .Y(_216_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_210_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_211_) );
OAI21X1 OAI21X1_58 ( .A(_210_), .B(_211_), .C(gnd), .Y(_212_) );
NAND2X1 NAND2X1_70 ( .A(_212_), .B(_216_), .Y(_0__0_) );
OAI21X1 OAI21X1_59 ( .A(_213_), .B(_210_), .C(_215_), .Y(_2__1_) );
INVX1 INVX1_81 ( .A(_2__1_), .Y(_220_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_221_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_222_) );
NAND3X1 NAND3X1_23 ( .A(_220_), .B(_222_), .C(_221_), .Y(_223_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_217_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_218_) );
OAI21X1 OAI21X1_60 ( .A(_217_), .B(_218_), .C(_2__1_), .Y(_219_) );
NAND2X1 NAND2X1_72 ( .A(_219_), .B(_223_), .Y(_0__1_) );
OAI21X1 OAI21X1_61 ( .A(_220_), .B(_217_), .C(_222_), .Y(_2__2_) );
INVX1 INVX1_82 ( .A(_2__2_), .Y(_227_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_228_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_229_) );
NAND3X1 NAND3X1_24 ( .A(_227_), .B(_229_), .C(_228_), .Y(_230_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_224_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_225_) );
OAI21X1 OAI21X1_62 ( .A(_224_), .B(_225_), .C(_2__2_), .Y(_226_) );
NAND2X1 NAND2X1_74 ( .A(_226_), .B(_230_), .Y(_0__2_) );
OAI21X1 OAI21X1_63 ( .A(_227_), .B(_224_), .C(_229_), .Y(_2__3_) );
INVX1 INVX1_83 ( .A(_2__3_), .Y(_234_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_235_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_236_) );
NAND3X1 NAND3X1_25 ( .A(_234_), .B(_236_), .C(_235_), .Y(_237_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_231_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_232_) );
OAI21X1 OAI21X1_64 ( .A(_231_), .B(_232_), .C(_2__3_), .Y(_233_) );
NAND2X1 NAND2X1_76 ( .A(_233_), .B(_237_), .Y(_0__3_) );
OAI21X1 OAI21X1_65 ( .A(_234_), .B(_231_), .C(_236_), .Y(_1_) );
INVX1 INVX1_84 ( .A(w_cout_1_), .Y(_241_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_242_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_243_) );
NAND3X1 NAND3X1_26 ( .A(_241_), .B(_243_), .C(_242_), .Y(_244_) );
NOR2X1 NOR2X1_108 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_238_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_239_) );
OAI21X1 OAI21X1_66 ( .A(_238_), .B(_239_), .C(w_cout_1_), .Y(_240_) );
NAND2X1 NAND2X1_78 ( .A(_240_), .B(_244_), .Y(_0__4_) );
OAI21X1 OAI21X1_67 ( .A(_241_), .B(_238_), .C(_243_), .Y(_5__1_) );
INVX1 INVX1_85 ( .A(_5__1_), .Y(_248_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_249_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_250_) );
NAND3X1 NAND3X1_27 ( .A(_248_), .B(_250_), .C(_249_), .Y(_251_) );
NOR2X1 NOR2X1_109 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_245_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_246_) );
OAI21X1 OAI21X1_68 ( .A(_245_), .B(_246_), .C(_5__1_), .Y(_247_) );
NAND2X1 NAND2X1_80 ( .A(_247_), .B(_251_), .Y(_0__5_) );
OAI21X1 OAI21X1_69 ( .A(_248_), .B(_245_), .C(_250_), .Y(_5__2_) );
INVX1 INVX1_86 ( .A(_5__2_), .Y(_255_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_256_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_257_) );
NAND3X1 NAND3X1_28 ( .A(_255_), .B(_257_), .C(_256_), .Y(_258_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_252_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_253_) );
OAI21X1 OAI21X1_70 ( .A(_252_), .B(_253_), .C(_5__2_), .Y(_254_) );
NAND2X1 NAND2X1_82 ( .A(_254_), .B(_258_), .Y(_0__6_) );
OAI21X1 OAI21X1_71 ( .A(_255_), .B(_252_), .C(_257_), .Y(_5__3_) );
INVX1 INVX1_87 ( .A(_5__3_), .Y(_262_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_263_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_264_) );
NAND3X1 NAND3X1_29 ( .A(_262_), .B(_264_), .C(_263_), .Y(_265_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_259_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_260_) );
OAI21X1 OAI21X1_72 ( .A(_259_), .B(_260_), .C(_5__3_), .Y(_261_) );
NAND2X1 NAND2X1_84 ( .A(_261_), .B(_265_), .Y(_0__7_) );
OAI21X1 OAI21X1_73 ( .A(_262_), .B(_259_), .C(_264_), .Y(_4_) );
INVX1 INVX1_88 ( .A(w_cout_2_), .Y(_269_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_270_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_271_) );
NAND3X1 NAND3X1_30 ( .A(_269_), .B(_271_), .C(_270_), .Y(_272_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_266_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_267_) );
OAI21X1 OAI21X1_74 ( .A(_266_), .B(_267_), .C(w_cout_2_), .Y(_268_) );
NAND2X1 NAND2X1_86 ( .A(_268_), .B(_272_), .Y(_0__8_) );
OAI21X1 OAI21X1_75 ( .A(_269_), .B(_266_), .C(_271_), .Y(_8__1_) );
INVX1 INVX1_89 ( .A(_8__1_), .Y(_276_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_277_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_278_) );
NAND3X1 NAND3X1_31 ( .A(_276_), .B(_278_), .C(_277_), .Y(_279_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_273_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_274_) );
OAI21X1 OAI21X1_76 ( .A(_273_), .B(_274_), .C(_8__1_), .Y(_275_) );
NAND2X1 NAND2X1_88 ( .A(_275_), .B(_279_), .Y(_0__9_) );
OAI21X1 OAI21X1_77 ( .A(_276_), .B(_273_), .C(_278_), .Y(_8__2_) );
INVX1 INVX1_90 ( .A(_8__2_), .Y(_283_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_284_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_285_) );
NAND3X1 NAND3X1_32 ( .A(_283_), .B(_285_), .C(_284_), .Y(_286_) );
NOR2X1 NOR2X1_114 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_280_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_281_) );
OAI21X1 OAI21X1_78 ( .A(_280_), .B(_281_), .C(_8__2_), .Y(_282_) );
NAND2X1 NAND2X1_90 ( .A(_282_), .B(_286_), .Y(_0__10_) );
OAI21X1 OAI21X1_79 ( .A(_283_), .B(_280_), .C(_285_), .Y(_8__3_) );
INVX1 INVX1_91 ( .A(_8__3_), .Y(_290_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_291_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_292_) );
NAND3X1 NAND3X1_33 ( .A(_290_), .B(_292_), .C(_291_), .Y(_293_) );
NOR2X1 NOR2X1_115 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_287_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_288_) );
OAI21X1 OAI21X1_80 ( .A(_287_), .B(_288_), .C(_8__3_), .Y(_289_) );
NAND2X1 NAND2X1_92 ( .A(_289_), .B(_293_), .Y(_0__11_) );
OAI21X1 OAI21X1_81 ( .A(_290_), .B(_287_), .C(_292_), .Y(_7_) );
INVX1 INVX1_92 ( .A(w_cout_3_), .Y(_297_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_298_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_299_) );
NAND3X1 NAND3X1_34 ( .A(_297_), .B(_299_), .C(_298_), .Y(_300_) );
NOR2X1 NOR2X1_116 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_294_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_295_) );
OAI21X1 OAI21X1_82 ( .A(_294_), .B(_295_), .C(w_cout_3_), .Y(_296_) );
NAND2X1 NAND2X1_94 ( .A(_296_), .B(_300_), .Y(_0__12_) );
OAI21X1 OAI21X1_83 ( .A(_297_), .B(_294_), .C(_299_), .Y(_11__1_) );
INVX1 INVX1_93 ( .A(_11__1_), .Y(_304_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_305_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_306_) );
NAND3X1 NAND3X1_35 ( .A(_304_), .B(_306_), .C(_305_), .Y(_307_) );
NOR2X1 NOR2X1_117 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_301_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_302_) );
OAI21X1 OAI21X1_84 ( .A(_301_), .B(_302_), .C(_11__1_), .Y(_303_) );
NAND2X1 NAND2X1_96 ( .A(_303_), .B(_307_), .Y(_0__13_) );
OAI21X1 OAI21X1_85 ( .A(_304_), .B(_301_), .C(_306_), .Y(_11__2_) );
INVX1 INVX1_94 ( .A(_11__2_), .Y(_311_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_312_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_313_) );
NAND3X1 NAND3X1_36 ( .A(_311_), .B(_313_), .C(_312_), .Y(_314_) );
NOR2X1 NOR2X1_118 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_308_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_309_) );
OAI21X1 OAI21X1_86 ( .A(_308_), .B(_309_), .C(_11__2_), .Y(_310_) );
NAND2X1 NAND2X1_98 ( .A(_310_), .B(_314_), .Y(_0__14_) );
OAI21X1 OAI21X1_87 ( .A(_311_), .B(_308_), .C(_313_), .Y(_11__3_) );
INVX1 INVX1_95 ( .A(_11__3_), .Y(_318_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_319_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_320_) );
NAND3X1 NAND3X1_37 ( .A(_318_), .B(_320_), .C(_319_), .Y(_321_) );
NOR2X1 NOR2X1_119 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_315_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_316_) );
OAI21X1 OAI21X1_88 ( .A(_315_), .B(_316_), .C(_11__3_), .Y(_317_) );
NAND2X1 NAND2X1_100 ( .A(_317_), .B(_321_), .Y(_0__15_) );
OAI21X1 OAI21X1_89 ( .A(_318_), .B(_315_), .C(_320_), .Y(_10_) );
INVX1 INVX1_96 ( .A(w_cout_4_), .Y(_325_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_326_) );
NAND2X1 NAND2X1_101 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_327_) );
NAND3X1 NAND3X1_38 ( .A(_325_), .B(_327_), .C(_326_), .Y(_328_) );
NOR2X1 NOR2X1_120 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_322_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_323_) );
OAI21X1 OAI21X1_90 ( .A(_322_), .B(_323_), .C(w_cout_4_), .Y(_324_) );
NAND2X1 NAND2X1_102 ( .A(_324_), .B(_328_), .Y(_0__16_) );
OAI21X1 OAI21X1_91 ( .A(_325_), .B(_322_), .C(_327_), .Y(_14__1_) );
INVX1 INVX1_97 ( .A(_14__1_), .Y(_332_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_333_) );
NAND2X1 NAND2X1_103 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_334_) );
NAND3X1 NAND3X1_39 ( .A(_332_), .B(_334_), .C(_333_), .Y(_335_) );
NOR2X1 NOR2X1_121 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_329_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_330_) );
OAI21X1 OAI21X1_92 ( .A(_329_), .B(_330_), .C(_14__1_), .Y(_331_) );
NAND2X1 NAND2X1_104 ( .A(_331_), .B(_335_), .Y(_0__17_) );
OAI21X1 OAI21X1_93 ( .A(_332_), .B(_329_), .C(_334_), .Y(_14__2_) );
INVX1 INVX1_98 ( .A(_14__2_), .Y(_339_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_340_) );
NAND2X1 NAND2X1_105 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_341_) );
NAND3X1 NAND3X1_40 ( .A(_339_), .B(_341_), .C(_340_), .Y(_342_) );
NOR2X1 NOR2X1_122 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_336_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_337_) );
OAI21X1 OAI21X1_94 ( .A(_336_), .B(_337_), .C(_14__2_), .Y(_338_) );
NAND2X1 NAND2X1_106 ( .A(_338_), .B(_342_), .Y(_0__18_) );
OAI21X1 OAI21X1_95 ( .A(_339_), .B(_336_), .C(_341_), .Y(_14__3_) );
INVX1 INVX1_99 ( .A(_14__3_), .Y(_346_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_347_) );
NAND2X1 NAND2X1_107 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_348_) );
NAND3X1 NAND3X1_41 ( .A(_346_), .B(_348_), .C(_347_), .Y(_349_) );
NOR2X1 NOR2X1_123 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_343_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_344_) );
OAI21X1 OAI21X1_96 ( .A(_343_), .B(_344_), .C(_14__3_), .Y(_345_) );
NAND2X1 NAND2X1_108 ( .A(_345_), .B(_349_), .Y(_0__19_) );
OAI21X1 OAI21X1_97 ( .A(_346_), .B(_343_), .C(_348_), .Y(_13_) );
INVX1 INVX1_100 ( .A(w_cout_5_), .Y(_353_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_354_) );
NAND2X1 NAND2X1_109 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_355_) );
NAND3X1 NAND3X1_42 ( .A(_353_), .B(_355_), .C(_354_), .Y(_356_) );
NOR2X1 NOR2X1_124 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_350_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_351_) );
OAI21X1 OAI21X1_98 ( .A(_350_), .B(_351_), .C(w_cout_5_), .Y(_352_) );
NAND2X1 NAND2X1_110 ( .A(_352_), .B(_356_), .Y(_0__20_) );
OAI21X1 OAI21X1_99 ( .A(_353_), .B(_350_), .C(_355_), .Y(_17__1_) );
INVX1 INVX1_101 ( .A(_17__1_), .Y(_360_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_361_) );
NAND2X1 NAND2X1_111 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_362_) );
NAND3X1 NAND3X1_43 ( .A(_360_), .B(_362_), .C(_361_), .Y(_363_) );
NOR2X1 NOR2X1_125 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_357_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_358_) );
OAI21X1 OAI21X1_100 ( .A(_357_), .B(_358_), .C(_17__1_), .Y(_359_) );
NAND2X1 NAND2X1_112 ( .A(_359_), .B(_363_), .Y(_0__21_) );
OAI21X1 OAI21X1_101 ( .A(_360_), .B(_357_), .C(_362_), .Y(_17__2_) );
INVX1 INVX1_102 ( .A(_17__2_), .Y(_367_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_368_) );
NAND2X1 NAND2X1_113 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_369_) );
NAND3X1 NAND3X1_44 ( .A(_367_), .B(_369_), .C(_368_), .Y(_370_) );
NOR2X1 NOR2X1_126 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_364_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_365_) );
OAI21X1 OAI21X1_102 ( .A(_364_), .B(_365_), .C(_17__2_), .Y(_366_) );
NAND2X1 NAND2X1_114 ( .A(_366_), .B(_370_), .Y(_0__22_) );
OAI21X1 OAI21X1_103 ( .A(_367_), .B(_364_), .C(_369_), .Y(_17__3_) );
INVX1 INVX1_103 ( .A(_17__3_), .Y(_374_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_375_) );
NAND2X1 NAND2X1_115 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_376_) );
NAND3X1 NAND3X1_45 ( .A(_374_), .B(_376_), .C(_375_), .Y(_377_) );
NOR2X1 NOR2X1_127 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_371_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_372_) );
OAI21X1 OAI21X1_104 ( .A(_371_), .B(_372_), .C(_17__3_), .Y(_373_) );
NAND2X1 NAND2X1_116 ( .A(_373_), .B(_377_), .Y(_0__23_) );
OAI21X1 OAI21X1_105 ( .A(_374_), .B(_371_), .C(_376_), .Y(_16_) );
INVX1 INVX1_104 ( .A(w_cout_6_), .Y(_381_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_382_) );
BUFX2 BUFX2_47 ( .A(cskip1_inst_sum), .Y(_0__44_) );
BUFX2 BUFX2_48 ( .A(gnd), .Y(_2__0_) );
BUFX2 BUFX2_49 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_50 ( .A(w_cout_1_), .Y(_5__0_) );
BUFX2 BUFX2_51 ( .A(_4_), .Y(_5__4_) );
BUFX2 BUFX2_52 ( .A(w_cout_2_), .Y(_8__0_) );
BUFX2 BUFX2_53 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_54 ( .A(w_cout_3_), .Y(_11__0_) );
BUFX2 BUFX2_55 ( .A(_10_), .Y(_11__4_) );
BUFX2 BUFX2_56 ( .A(w_cout_4_), .Y(_14__0_) );
BUFX2 BUFX2_57 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_58 ( .A(w_cout_5_), .Y(_17__0_) );
BUFX2 BUFX2_59 ( .A(_16_), .Y(_17__4_) );
BUFX2 BUFX2_60 ( .A(w_cout_6_), .Y(_20__0_) );
BUFX2 BUFX2_61 ( .A(_19_), .Y(_20__4_) );
BUFX2 BUFX2_62 ( .A(w_cout_7_), .Y(_23__0_) );
BUFX2 BUFX2_63 ( .A(_22_), .Y(_23__4_) );
BUFX2 BUFX2_64 ( .A(w_cout_8_), .Y(_26__0_) );
BUFX2 BUFX2_65 ( .A(_25_), .Y(_26__4_) );
BUFX2 BUFX2_66 ( .A(w_cout_9_), .Y(_29__0_) );
BUFX2 BUFX2_67 ( .A(_28_), .Y(_29__4_) );
BUFX2 BUFX2_68 ( .A(w_cout_10_), .Y(_32__0_) );
BUFX2 BUFX2_69 ( .A(_31_), .Y(_32__4_) );
BUFX2 BUFX2_70 ( .A(cskip1_inst_cin), .Y(cskip1_inst_rca0_w_CARRY_0_) );
BUFX2 BUFX2_71 ( .A(cskip1_inst_cout0), .Y(cskip1_inst_rca0_w_CARRY_4_) );
BUFX2 BUFX2_72 ( .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_73 ( .A(cskip1_inst_cin), .Y(w_cout_11_) );
endmodule
