module cla_8bit (i_add1, i_add2, o_result);

input [7:0] i_add1;
input [7:0] i_add2;
output [8:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

OAI21X1 OAI21X1_1 ( .A(i_add2[4]), .B(i_add1[4]), .C(_12_), .Y(_13_) );
INVX1 INVX1_1 ( .A(_13_), .Y(w_C_5_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_14_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_15_) );
OAI21X1 OAI21X1_2 ( .A(_15_), .B(_13_), .C(_14_), .Y(w_C_6_) );
OR2X2 OR2X2_1 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_16_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_17_) );
INVX1 INVX1_2 ( .A(_17_), .Y(_18_) );
INVX1 INVX1_3 ( .A(_15_), .Y(_19_) );
NAND3X1 NAND3X1_1 ( .A(_18_), .B(_19_), .C(_12_), .Y(_20_) );
NAND2X1 NAND2X1_2 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_21_) );
NAND3X1 NAND3X1_2 ( .A(_14_), .B(_21_), .C(_20_), .Y(_22_) );
AND2X2 AND2X2_1 ( .A(_22_), .B(_16_), .Y(w_C_7_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_23_) );
OR2X2 OR2X2_2 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_24_) );
NAND3X1 NAND3X1_3 ( .A(_16_), .B(_24_), .C(_22_), .Y(_25_) );
NAND2X1 NAND2X1_4 ( .A(_23_), .B(_25_), .Y(w_C_8_) );
BUFX2 BUFX2_1 ( .A(_26__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_26__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_26__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_26__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_26__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_26__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_26__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_26__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(w_C_8_), .Y(o_result[8]) );
INVX1 INVX1_4 ( .A(w_C_4_), .Y(_30_) );
OR2X2 OR2X2_3 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_31_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_32_) );
NAND3X1 NAND3X1_4 ( .A(_30_), .B(_32_), .C(_31_), .Y(_33_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_27_) );
AND2X2 AND2X2_2 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_28_) );
OAI21X1 OAI21X1_3 ( .A(_27_), .B(_28_), .C(w_C_4_), .Y(_29_) );
NAND2X1 NAND2X1_6 ( .A(_29_), .B(_33_), .Y(_26__4_) );
INVX1 INVX1_5 ( .A(w_C_5_), .Y(_37_) );
OR2X2 OR2X2_4 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_38_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_39_) );
NAND3X1 NAND3X1_5 ( .A(_37_), .B(_39_), .C(_38_), .Y(_40_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_34_) );
AND2X2 AND2X2_3 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_35_) );
OAI21X1 OAI21X1_4 ( .A(_34_), .B(_35_), .C(w_C_5_), .Y(_36_) );
NAND2X1 NAND2X1_8 ( .A(_36_), .B(_40_), .Y(_26__5_) );
INVX1 INVX1_6 ( .A(w_C_6_), .Y(_44_) );
OR2X2 OR2X2_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_45_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_46_) );
NAND3X1 NAND3X1_6 ( .A(_44_), .B(_46_), .C(_45_), .Y(_47_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_41_) );
AND2X2 AND2X2_4 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_42_) );
OAI21X1 OAI21X1_5 ( .A(_41_), .B(_42_), .C(w_C_6_), .Y(_43_) );
NAND2X1 NAND2X1_10 ( .A(_43_), .B(_47_), .Y(_26__6_) );
INVX1 INVX1_7 ( .A(w_C_7_), .Y(_51_) );
OR2X2 OR2X2_6 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_52_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_53_) );
NAND3X1 NAND3X1_7 ( .A(_51_), .B(_53_), .C(_52_), .Y(_54_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_48_) );
AND2X2 AND2X2_5 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_49_) );
OAI21X1 OAI21X1_6 ( .A(_48_), .B(_49_), .C(w_C_7_), .Y(_50_) );
NAND2X1 NAND2X1_12 ( .A(_50_), .B(_54_), .Y(_26__7_) );
INVX1 INVX1_8 ( .A(gnd), .Y(_58_) );
OR2X2 OR2X2_7 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_59_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_60_) );
NAND3X1 NAND3X1_8 ( .A(_58_), .B(_60_), .C(_59_), .Y(_61_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_55_) );
AND2X2 AND2X2_6 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_56_) );
OAI21X1 OAI21X1_7 ( .A(_55_), .B(_56_), .C(gnd), .Y(_57_) );
NAND2X1 NAND2X1_14 ( .A(_57_), .B(_61_), .Y(_26__0_) );
INVX1 INVX1_9 ( .A(w_C_1_), .Y(_65_) );
OR2X2 OR2X2_8 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_66_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_67_) );
NAND3X1 NAND3X1_9 ( .A(_65_), .B(_67_), .C(_66_), .Y(_68_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_62_) );
AND2X2 AND2X2_7 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_63_) );
OAI21X1 OAI21X1_8 ( .A(_62_), .B(_63_), .C(w_C_1_), .Y(_64_) );
NAND2X1 NAND2X1_16 ( .A(_64_), .B(_68_), .Y(_26__1_) );
INVX1 INVX1_10 ( .A(w_C_2_), .Y(_72_) );
OR2X2 OR2X2_9 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_73_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_74_) );
NAND3X1 NAND3X1_10 ( .A(_72_), .B(_74_), .C(_73_), .Y(_75_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_69_) );
AND2X2 AND2X2_8 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_70_) );
OAI21X1 OAI21X1_9 ( .A(_69_), .B(_70_), .C(w_C_2_), .Y(_71_) );
NAND2X1 NAND2X1_18 ( .A(_71_), .B(_75_), .Y(_26__2_) );
INVX1 INVX1_11 ( .A(w_C_3_), .Y(_79_) );
OR2X2 OR2X2_10 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_80_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_81_) );
NAND3X1 NAND3X1_11 ( .A(_79_), .B(_81_), .C(_80_), .Y(_82_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_76_) );
AND2X2 AND2X2_9 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_77_) );
OAI21X1 OAI21X1_10 ( .A(_76_), .B(_77_), .C(w_C_3_), .Y(_78_) );
NAND2X1 NAND2X1_20 ( .A(_78_), .B(_82_), .Y(_26__3_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_12 ( .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_12 ( .A(_1_), .B(_2_), .Y(w_C_2_) );
INVX1 INVX1_13 ( .A(i_add2[2]), .Y(_3_) );
INVX1 INVX1_14 ( .A(i_add1[2]), .Y(_4_) );
NAND2X1 NAND2X1_22 ( .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
OAI21X1 OAI21X1_11 ( .A(_1_), .B(_2_), .C(_6_), .Y(_7_) );
AND2X2 AND2X2_10 ( .A(_7_), .B(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
OR2X2 OR2X2_11 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_12 ( .A(_5_), .B(_9_), .C(_7_), .Y(_10_) );
NAND2X1 NAND2X1_25 ( .A(_8_), .B(_10_), .Y(w_C_4_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
NAND3X1 NAND3X1_13 ( .A(_8_), .B(_11_), .C(_10_), .Y(_12_) );
BUFX2 BUFX2_10 ( .A(w_C_8_), .Y(_26__8_) );
BUFX2 BUFX2_11 ( .A(gnd), .Y(w_C_0_) );
endmodule
