module csa_47bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term1[45], i_add_term1[46], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], i_add_term2[45], i_add_term2[46], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], sum[45], sum[46], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term1[45];
input i_add_term1[46];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
input i_add_term2[45];
input i_add_term2[46];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output sum[45];
output sum[46];
output cout;

INVX1 INVX1_1 ( .A(_15__0_), .Y(_195_) );
NAND2X1 NAND2X1_1 ( .A(_16__0_), .B(w_cout_2_), .Y(_196_) );
OAI21X1 OAI21X1_1 ( .A(w_cout_2_), .B(_195_), .C(_196_), .Y(_0__12_) );
INVX1 INVX1_2 ( .A(_15__1_), .Y(_197_) );
NAND2X1 NAND2X1_2 ( .A(w_cout_2_), .B(_16__1_), .Y(_198_) );
OAI21X1 OAI21X1_2 ( .A(w_cout_2_), .B(_197_), .C(_198_), .Y(_0__13_) );
INVX1 INVX1_3 ( .A(_15__2_), .Y(_199_) );
NAND2X1 NAND2X1_3 ( .A(w_cout_2_), .B(_16__2_), .Y(_200_) );
OAI21X1 OAI21X1_3 ( .A(w_cout_2_), .B(_199_), .C(_200_), .Y(_0__14_) );
INVX1 INVX1_4 ( .A(_15__3_), .Y(_201_) );
NAND2X1 NAND2X1_4 ( .A(w_cout_2_), .B(_16__3_), .Y(_202_) );
OAI21X1 OAI21X1_4 ( .A(w_cout_2_), .B(_201_), .C(_202_), .Y(_0__15_) );
INVX1 INVX1_5 ( .A(1'b0), .Y(_206_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_207_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_208_) );
NAND3X1 NAND3X1_1 ( .A(_206_), .B(_208_), .C(_207_), .Y(_209_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_203_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_204_) );
OAI21X1 OAI21X1_5 ( .A(_203_), .B(_204_), .C(1'b0), .Y(_205_) );
NAND2X1 NAND2X1_6 ( .A(_205_), .B(_209_), .Y(_15__0_) );
OAI21X1 OAI21X1_6 ( .A(_206_), .B(_203_), .C(_208_), .Y(_17__1_) );
INVX1 INVX1_6 ( .A(_17__3_), .Y(_213_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_214_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_215_) );
NAND3X1 NAND3X1_2 ( .A(_213_), .B(_215_), .C(_214_), .Y(_216_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_210_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_211_) );
OAI21X1 OAI21X1_7 ( .A(_210_), .B(_211_), .C(_17__3_), .Y(_212_) );
NAND2X1 NAND2X1_8 ( .A(_212_), .B(_216_), .Y(_15__3_) );
OAI21X1 OAI21X1_8 ( .A(_213_), .B(_210_), .C(_215_), .Y(_13_) );
INVX1 INVX1_7 ( .A(_17__1_), .Y(_220_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_221_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_222_) );
NAND3X1 NAND3X1_3 ( .A(_220_), .B(_222_), .C(_221_), .Y(_223_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_217_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_218_) );
OAI21X1 OAI21X1_9 ( .A(_217_), .B(_218_), .C(_17__1_), .Y(_219_) );
NAND2X1 NAND2X1_10 ( .A(_219_), .B(_223_), .Y(_15__1_) );
OAI21X1 OAI21X1_10 ( .A(_220_), .B(_217_), .C(_222_), .Y(_17__2_) );
INVX1 INVX1_8 ( .A(_17__2_), .Y(_227_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_228_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_229_) );
NAND3X1 NAND3X1_4 ( .A(_227_), .B(_229_), .C(_228_), .Y(_230_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_224_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_225_) );
OAI21X1 OAI21X1_11 ( .A(_224_), .B(_225_), .C(_17__2_), .Y(_226_) );
NAND2X1 NAND2X1_12 ( .A(_226_), .B(_230_), .Y(_15__2_) );
OAI21X1 OAI21X1_12 ( .A(_227_), .B(_224_), .C(_229_), .Y(_17__3_) );
INVX1 INVX1_9 ( .A(1'b1), .Y(_234_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_235_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_236_) );
NAND3X1 NAND3X1_5 ( .A(_234_), .B(_236_), .C(_235_), .Y(_237_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_231_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_232_) );
OAI21X1 OAI21X1_13 ( .A(_231_), .B(_232_), .C(1'b1), .Y(_233_) );
NAND2X1 NAND2X1_14 ( .A(_233_), .B(_237_), .Y(_16__0_) );
OAI21X1 OAI21X1_14 ( .A(_234_), .B(_231_), .C(_236_), .Y(_18__1_) );
INVX1 INVX1_10 ( .A(_18__3_), .Y(_241_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_242_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_243_) );
NAND3X1 NAND3X1_6 ( .A(_241_), .B(_243_), .C(_242_), .Y(_244_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_238_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_239_) );
OAI21X1 OAI21X1_15 ( .A(_238_), .B(_239_), .C(_18__3_), .Y(_240_) );
NAND2X1 NAND2X1_16 ( .A(_240_), .B(_244_), .Y(_16__3_) );
OAI21X1 OAI21X1_16 ( .A(_241_), .B(_238_), .C(_243_), .Y(_14_) );
INVX1 INVX1_11 ( .A(_18__1_), .Y(_248_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_249_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_250_) );
NAND3X1 NAND3X1_7 ( .A(_248_), .B(_250_), .C(_249_), .Y(_251_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_245_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_246_) );
OAI21X1 OAI21X1_17 ( .A(_245_), .B(_246_), .C(_18__1_), .Y(_247_) );
NAND2X1 NAND2X1_18 ( .A(_247_), .B(_251_), .Y(_16__1_) );
OAI21X1 OAI21X1_18 ( .A(_248_), .B(_245_), .C(_250_), .Y(_18__2_) );
INVX1 INVX1_12 ( .A(_18__2_), .Y(_255_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_256_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_257_) );
NAND3X1 NAND3X1_8 ( .A(_255_), .B(_257_), .C(_256_), .Y(_258_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_252_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_253_) );
OAI21X1 OAI21X1_19 ( .A(_252_), .B(_253_), .C(_18__2_), .Y(_254_) );
NAND2X1 NAND2X1_20 ( .A(_254_), .B(_258_), .Y(_16__2_) );
OAI21X1 OAI21X1_20 ( .A(_255_), .B(_252_), .C(_257_), .Y(_18__3_) );
INVX1 INVX1_13 ( .A(_19_), .Y(_259_) );
NAND2X1 NAND2X1_21 ( .A(_20_), .B(w_cout_3_), .Y(_260_) );
OAI21X1 OAI21X1_21 ( .A(w_cout_3_), .B(_259_), .C(_260_), .Y(w_cout_4_) );
INVX1 INVX1_14 ( .A(_21__0_), .Y(_261_) );
NAND2X1 NAND2X1_22 ( .A(_22__0_), .B(w_cout_3_), .Y(_262_) );
OAI21X1 OAI21X1_22 ( .A(w_cout_3_), .B(_261_), .C(_262_), .Y(_0__16_) );
INVX1 INVX1_15 ( .A(_21__1_), .Y(_263_) );
NAND2X1 NAND2X1_23 ( .A(w_cout_3_), .B(_22__1_), .Y(_264_) );
OAI21X1 OAI21X1_23 ( .A(w_cout_3_), .B(_263_), .C(_264_), .Y(_0__17_) );
INVX1 INVX1_16 ( .A(_21__2_), .Y(_265_) );
NAND2X1 NAND2X1_24 ( .A(w_cout_3_), .B(_22__2_), .Y(_266_) );
OAI21X1 OAI21X1_24 ( .A(w_cout_3_), .B(_265_), .C(_266_), .Y(_0__18_) );
INVX1 INVX1_17 ( .A(_21__3_), .Y(_267_) );
NAND2X1 NAND2X1_25 ( .A(w_cout_3_), .B(_22__3_), .Y(_268_) );
OAI21X1 OAI21X1_25 ( .A(w_cout_3_), .B(_267_), .C(_268_), .Y(_0__19_) );
INVX1 INVX1_18 ( .A(1'b0), .Y(_272_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_273_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_274_) );
NAND3X1 NAND3X1_9 ( .A(_272_), .B(_274_), .C(_273_), .Y(_275_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_269_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_270_) );
OAI21X1 OAI21X1_26 ( .A(_269_), .B(_270_), .C(1'b0), .Y(_271_) );
NAND2X1 NAND2X1_27 ( .A(_271_), .B(_275_), .Y(_21__0_) );
OAI21X1 OAI21X1_27 ( .A(_272_), .B(_269_), .C(_274_), .Y(_23__1_) );
INVX1 INVX1_19 ( .A(_23__3_), .Y(_279_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_280_) );
NAND2X1 NAND2X1_28 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_281_) );
NAND3X1 NAND3X1_10 ( .A(_279_), .B(_281_), .C(_280_), .Y(_282_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_276_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_277_) );
OAI21X1 OAI21X1_28 ( .A(_276_), .B(_277_), .C(_23__3_), .Y(_278_) );
NAND2X1 NAND2X1_29 ( .A(_278_), .B(_282_), .Y(_21__3_) );
OAI21X1 OAI21X1_29 ( .A(_279_), .B(_276_), .C(_281_), .Y(_19_) );
INVX1 INVX1_20 ( .A(_23__1_), .Y(_286_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_287_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_288_) );
NAND3X1 NAND3X1_11 ( .A(_286_), .B(_288_), .C(_287_), .Y(_289_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_283_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_284_) );
OAI21X1 OAI21X1_30 ( .A(_283_), .B(_284_), .C(_23__1_), .Y(_285_) );
NAND2X1 NAND2X1_31 ( .A(_285_), .B(_289_), .Y(_21__1_) );
OAI21X1 OAI21X1_31 ( .A(_286_), .B(_283_), .C(_288_), .Y(_23__2_) );
INVX1 INVX1_21 ( .A(_23__2_), .Y(_293_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_294_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_295_) );
NAND3X1 NAND3X1_12 ( .A(_293_), .B(_295_), .C(_294_), .Y(_296_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_290_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_291_) );
OAI21X1 OAI21X1_32 ( .A(_290_), .B(_291_), .C(_23__2_), .Y(_292_) );
NAND2X1 NAND2X1_33 ( .A(_292_), .B(_296_), .Y(_21__2_) );
OAI21X1 OAI21X1_33 ( .A(_293_), .B(_290_), .C(_295_), .Y(_23__3_) );
INVX1 INVX1_22 ( .A(1'b1), .Y(_300_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_301_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_302_) );
NAND3X1 NAND3X1_13 ( .A(_300_), .B(_302_), .C(_301_), .Y(_303_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_297_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_298_) );
OAI21X1 OAI21X1_34 ( .A(_297_), .B(_298_), .C(1'b1), .Y(_299_) );
NAND2X1 NAND2X1_35 ( .A(_299_), .B(_303_), .Y(_22__0_) );
OAI21X1 OAI21X1_35 ( .A(_300_), .B(_297_), .C(_302_), .Y(_24__1_) );
INVX1 INVX1_23 ( .A(_24__3_), .Y(_307_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_308_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_309_) );
NAND3X1 NAND3X1_14 ( .A(_307_), .B(_309_), .C(_308_), .Y(_310_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_304_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_305_) );
OAI21X1 OAI21X1_36 ( .A(_304_), .B(_305_), .C(_24__3_), .Y(_306_) );
NAND2X1 NAND2X1_37 ( .A(_306_), .B(_310_), .Y(_22__3_) );
OAI21X1 OAI21X1_37 ( .A(_307_), .B(_304_), .C(_309_), .Y(_20_) );
INVX1 INVX1_24 ( .A(_24__1_), .Y(_314_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_315_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_316_) );
NAND3X1 NAND3X1_15 ( .A(_314_), .B(_316_), .C(_315_), .Y(_317_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_311_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_312_) );
OAI21X1 OAI21X1_38 ( .A(_311_), .B(_312_), .C(_24__1_), .Y(_313_) );
NAND2X1 NAND2X1_39 ( .A(_313_), .B(_317_), .Y(_22__1_) );
OAI21X1 OAI21X1_39 ( .A(_314_), .B(_311_), .C(_316_), .Y(_24__2_) );
INVX1 INVX1_25 ( .A(_24__2_), .Y(_321_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_322_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_323_) );
NAND3X1 NAND3X1_16 ( .A(_321_), .B(_323_), .C(_322_), .Y(_324_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_318_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_319_) );
OAI21X1 OAI21X1_40 ( .A(_318_), .B(_319_), .C(_24__2_), .Y(_320_) );
NAND2X1 NAND2X1_41 ( .A(_320_), .B(_324_), .Y(_22__2_) );
OAI21X1 OAI21X1_41 ( .A(_321_), .B(_318_), .C(_323_), .Y(_24__3_) );
INVX1 INVX1_26 ( .A(_25_), .Y(_325_) );
NAND2X1 NAND2X1_42 ( .A(_26_), .B(w_cout_4_), .Y(_326_) );
OAI21X1 OAI21X1_42 ( .A(w_cout_4_), .B(_325_), .C(_326_), .Y(w_cout_5_) );
INVX1 INVX1_27 ( .A(_27__0_), .Y(_327_) );
NAND2X1 NAND2X1_43 ( .A(_28__0_), .B(w_cout_4_), .Y(_328_) );
OAI21X1 OAI21X1_43 ( .A(w_cout_4_), .B(_327_), .C(_328_), .Y(_0__20_) );
INVX1 INVX1_28 ( .A(_27__1_), .Y(_329_) );
NAND2X1 NAND2X1_44 ( .A(w_cout_4_), .B(_28__1_), .Y(_330_) );
OAI21X1 OAI21X1_44 ( .A(w_cout_4_), .B(_329_), .C(_330_), .Y(_0__21_) );
INVX1 INVX1_29 ( .A(_27__2_), .Y(_331_) );
NAND2X1 NAND2X1_45 ( .A(w_cout_4_), .B(_28__2_), .Y(_332_) );
OAI21X1 OAI21X1_45 ( .A(w_cout_4_), .B(_331_), .C(_332_), .Y(_0__22_) );
INVX1 INVX1_30 ( .A(_27__3_), .Y(_333_) );
NAND2X1 NAND2X1_46 ( .A(w_cout_4_), .B(_28__3_), .Y(_334_) );
OAI21X1 OAI21X1_46 ( .A(w_cout_4_), .B(_333_), .C(_334_), .Y(_0__23_) );
INVX1 INVX1_31 ( .A(1'b0), .Y(_338_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_339_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_340_) );
NAND3X1 NAND3X1_17 ( .A(_338_), .B(_340_), .C(_339_), .Y(_341_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_335_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_336_) );
OAI21X1 OAI21X1_47 ( .A(_335_), .B(_336_), .C(1'b0), .Y(_337_) );
NAND2X1 NAND2X1_48 ( .A(_337_), .B(_341_), .Y(_27__0_) );
OAI21X1 OAI21X1_48 ( .A(_338_), .B(_335_), .C(_340_), .Y(_29__1_) );
INVX1 INVX1_32 ( .A(_29__3_), .Y(_345_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_346_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_347_) );
NAND3X1 NAND3X1_18 ( .A(_345_), .B(_347_), .C(_346_), .Y(_348_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_342_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_343_) );
OAI21X1 OAI21X1_49 ( .A(_342_), .B(_343_), .C(_29__3_), .Y(_344_) );
NAND2X1 NAND2X1_50 ( .A(_344_), .B(_348_), .Y(_27__3_) );
OAI21X1 OAI21X1_50 ( .A(_345_), .B(_342_), .C(_347_), .Y(_25_) );
INVX1 INVX1_33 ( .A(_29__1_), .Y(_352_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_353_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_354_) );
NAND3X1 NAND3X1_19 ( .A(_352_), .B(_354_), .C(_353_), .Y(_355_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_349_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_350_) );
OAI21X1 OAI21X1_51 ( .A(_349_), .B(_350_), .C(_29__1_), .Y(_351_) );
NAND2X1 NAND2X1_52 ( .A(_351_), .B(_355_), .Y(_27__1_) );
OAI21X1 OAI21X1_52 ( .A(_352_), .B(_349_), .C(_354_), .Y(_29__2_) );
INVX1 INVX1_34 ( .A(_29__2_), .Y(_359_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_360_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_361_) );
NAND3X1 NAND3X1_20 ( .A(_359_), .B(_361_), .C(_360_), .Y(_362_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_356_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_357_) );
OAI21X1 OAI21X1_53 ( .A(_356_), .B(_357_), .C(_29__2_), .Y(_358_) );
NAND2X1 NAND2X1_54 ( .A(_358_), .B(_362_), .Y(_27__2_) );
OAI21X1 OAI21X1_54 ( .A(_359_), .B(_356_), .C(_361_), .Y(_29__3_) );
INVX1 INVX1_35 ( .A(1'b1), .Y(_366_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_367_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_368_) );
NAND3X1 NAND3X1_21 ( .A(_366_), .B(_368_), .C(_367_), .Y(_369_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_363_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_364_) );
OAI21X1 OAI21X1_55 ( .A(_363_), .B(_364_), .C(1'b1), .Y(_365_) );
NAND2X1 NAND2X1_56 ( .A(_365_), .B(_369_), .Y(_28__0_) );
OAI21X1 OAI21X1_56 ( .A(_366_), .B(_363_), .C(_368_), .Y(_30__1_) );
INVX1 INVX1_36 ( .A(_30__3_), .Y(_373_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_374_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_375_) );
NAND3X1 NAND3X1_22 ( .A(_373_), .B(_375_), .C(_374_), .Y(_376_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_370_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_371_) );
OAI21X1 OAI21X1_57 ( .A(_370_), .B(_371_), .C(_30__3_), .Y(_372_) );
NAND2X1 NAND2X1_58 ( .A(_372_), .B(_376_), .Y(_28__3_) );
OAI21X1 OAI21X1_58 ( .A(_373_), .B(_370_), .C(_375_), .Y(_26_) );
INVX1 INVX1_37 ( .A(_30__1_), .Y(_380_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_381_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_382_) );
NAND3X1 NAND3X1_23 ( .A(_380_), .B(_382_), .C(_381_), .Y(_383_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_377_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_378_) );
OAI21X1 OAI21X1_59 ( .A(_377_), .B(_378_), .C(_30__1_), .Y(_379_) );
NAND2X1 NAND2X1_60 ( .A(_379_), .B(_383_), .Y(_28__1_) );
OAI21X1 OAI21X1_60 ( .A(_380_), .B(_377_), .C(_382_), .Y(_30__2_) );
INVX1 INVX1_38 ( .A(_30__2_), .Y(_387_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_388_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_389_) );
NAND3X1 NAND3X1_24 ( .A(_387_), .B(_389_), .C(_388_), .Y(_390_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_384_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_385_) );
OAI21X1 OAI21X1_61 ( .A(_384_), .B(_385_), .C(_30__2_), .Y(_386_) );
NAND2X1 NAND2X1_62 ( .A(_386_), .B(_390_), .Y(_28__2_) );
OAI21X1 OAI21X1_62 ( .A(_387_), .B(_384_), .C(_389_), .Y(_30__3_) );
INVX1 INVX1_39 ( .A(_31_), .Y(_391_) );
NAND2X1 NAND2X1_63 ( .A(_32_), .B(w_cout_5_), .Y(_392_) );
OAI21X1 OAI21X1_63 ( .A(w_cout_5_), .B(_391_), .C(_392_), .Y(w_cout_6_) );
INVX1 INVX1_40 ( .A(_33__0_), .Y(_393_) );
NAND2X1 NAND2X1_64 ( .A(_34__0_), .B(w_cout_5_), .Y(_394_) );
OAI21X1 OAI21X1_64 ( .A(w_cout_5_), .B(_393_), .C(_394_), .Y(_0__24_) );
INVX1 INVX1_41 ( .A(_33__1_), .Y(_395_) );
NAND2X1 NAND2X1_65 ( .A(w_cout_5_), .B(_34__1_), .Y(_396_) );
OAI21X1 OAI21X1_65 ( .A(w_cout_5_), .B(_395_), .C(_396_), .Y(_0__25_) );
INVX1 INVX1_42 ( .A(_33__2_), .Y(_397_) );
NAND2X1 NAND2X1_66 ( .A(w_cout_5_), .B(_34__2_), .Y(_398_) );
OAI21X1 OAI21X1_66 ( .A(w_cout_5_), .B(_397_), .C(_398_), .Y(_0__26_) );
INVX1 INVX1_43 ( .A(_33__3_), .Y(_399_) );
NAND2X1 NAND2X1_67 ( .A(w_cout_5_), .B(_34__3_), .Y(_400_) );
OAI21X1 OAI21X1_67 ( .A(w_cout_5_), .B(_399_), .C(_400_), .Y(_0__27_) );
INVX1 INVX1_44 ( .A(1'b0), .Y(_404_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_405_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_406_) );
NAND3X1 NAND3X1_25 ( .A(_404_), .B(_406_), .C(_405_), .Y(_407_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_401_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_402_) );
OAI21X1 OAI21X1_68 ( .A(_401_), .B(_402_), .C(1'b0), .Y(_403_) );
NAND2X1 NAND2X1_69 ( .A(_403_), .B(_407_), .Y(_33__0_) );
OAI21X1 OAI21X1_69 ( .A(_404_), .B(_401_), .C(_406_), .Y(_35__1_) );
INVX1 INVX1_45 ( .A(_35__3_), .Y(_411_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_412_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_413_) );
NAND3X1 NAND3X1_26 ( .A(_411_), .B(_413_), .C(_412_), .Y(_414_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_408_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_409_) );
OAI21X1 OAI21X1_70 ( .A(_408_), .B(_409_), .C(_35__3_), .Y(_410_) );
NAND2X1 NAND2X1_71 ( .A(_410_), .B(_414_), .Y(_33__3_) );
OAI21X1 OAI21X1_71 ( .A(_411_), .B(_408_), .C(_413_), .Y(_31_) );
INVX1 INVX1_46 ( .A(_35__1_), .Y(_418_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_419_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_420_) );
NAND3X1 NAND3X1_27 ( .A(_418_), .B(_420_), .C(_419_), .Y(_421_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_415_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_416_) );
OAI21X1 OAI21X1_72 ( .A(_415_), .B(_416_), .C(_35__1_), .Y(_417_) );
NAND2X1 NAND2X1_73 ( .A(_417_), .B(_421_), .Y(_33__1_) );
OAI21X1 OAI21X1_73 ( .A(_418_), .B(_415_), .C(_420_), .Y(_35__2_) );
INVX1 INVX1_47 ( .A(_35__2_), .Y(_425_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_426_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_427_) );
NAND3X1 NAND3X1_28 ( .A(_425_), .B(_427_), .C(_426_), .Y(_428_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_422_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_423_) );
OAI21X1 OAI21X1_74 ( .A(_422_), .B(_423_), .C(_35__2_), .Y(_424_) );
NAND2X1 NAND2X1_75 ( .A(_424_), .B(_428_), .Y(_33__2_) );
OAI21X1 OAI21X1_75 ( .A(_425_), .B(_422_), .C(_427_), .Y(_35__3_) );
INVX1 INVX1_48 ( .A(1'b1), .Y(_432_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_433_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_434_) );
NAND3X1 NAND3X1_29 ( .A(_432_), .B(_434_), .C(_433_), .Y(_435_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_429_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_430_) );
OAI21X1 OAI21X1_76 ( .A(_429_), .B(_430_), .C(1'b1), .Y(_431_) );
NAND2X1 NAND2X1_77 ( .A(_431_), .B(_435_), .Y(_34__0_) );
OAI21X1 OAI21X1_77 ( .A(_432_), .B(_429_), .C(_434_), .Y(_36__1_) );
INVX1 INVX1_49 ( .A(_36__3_), .Y(_439_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_440_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_441_) );
NAND3X1 NAND3X1_30 ( .A(_439_), .B(_441_), .C(_440_), .Y(_442_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_436_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_437_) );
OAI21X1 OAI21X1_78 ( .A(_436_), .B(_437_), .C(_36__3_), .Y(_438_) );
NAND2X1 NAND2X1_79 ( .A(_438_), .B(_442_), .Y(_34__3_) );
OAI21X1 OAI21X1_79 ( .A(_439_), .B(_436_), .C(_441_), .Y(_32_) );
INVX1 INVX1_50 ( .A(_36__1_), .Y(_446_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_447_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_448_) );
NAND3X1 NAND3X1_31 ( .A(_446_), .B(_448_), .C(_447_), .Y(_449_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_443_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_444_) );
OAI21X1 OAI21X1_80 ( .A(_443_), .B(_444_), .C(_36__1_), .Y(_445_) );
NAND2X1 NAND2X1_81 ( .A(_445_), .B(_449_), .Y(_34__1_) );
OAI21X1 OAI21X1_81 ( .A(_446_), .B(_443_), .C(_448_), .Y(_36__2_) );
INVX1 INVX1_51 ( .A(_36__2_), .Y(_453_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_454_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_455_) );
NAND3X1 NAND3X1_32 ( .A(_453_), .B(_455_), .C(_454_), .Y(_456_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_450_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_451_) );
OAI21X1 OAI21X1_82 ( .A(_450_), .B(_451_), .C(_36__2_), .Y(_452_) );
NAND2X1 NAND2X1_83 ( .A(_452_), .B(_456_), .Y(_34__2_) );
OAI21X1 OAI21X1_83 ( .A(_453_), .B(_450_), .C(_455_), .Y(_36__3_) );
INVX1 INVX1_52 ( .A(_37_), .Y(_457_) );
NAND2X1 NAND2X1_84 ( .A(_38_), .B(w_cout_6_), .Y(_458_) );
OAI21X1 OAI21X1_84 ( .A(w_cout_6_), .B(_457_), .C(_458_), .Y(w_cout_7_) );
INVX1 INVX1_53 ( .A(_39__0_), .Y(_459_) );
NAND2X1 NAND2X1_85 ( .A(_40__0_), .B(w_cout_6_), .Y(_460_) );
OAI21X1 OAI21X1_85 ( .A(w_cout_6_), .B(_459_), .C(_460_), .Y(_0__28_) );
INVX1 INVX1_54 ( .A(_39__1_), .Y(_461_) );
NAND2X1 NAND2X1_86 ( .A(w_cout_6_), .B(_40__1_), .Y(_462_) );
OAI21X1 OAI21X1_86 ( .A(w_cout_6_), .B(_461_), .C(_462_), .Y(_0__29_) );
INVX1 INVX1_55 ( .A(_39__2_), .Y(_463_) );
NAND2X1 NAND2X1_87 ( .A(w_cout_6_), .B(_40__2_), .Y(_464_) );
OAI21X1 OAI21X1_87 ( .A(w_cout_6_), .B(_463_), .C(_464_), .Y(_0__30_) );
INVX1 INVX1_56 ( .A(_39__3_), .Y(_465_) );
NAND2X1 NAND2X1_88 ( .A(w_cout_6_), .B(_40__3_), .Y(_466_) );
OAI21X1 OAI21X1_88 ( .A(w_cout_6_), .B(_465_), .C(_466_), .Y(_0__31_) );
INVX1 INVX1_57 ( .A(1'b0), .Y(_470_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_471_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_472_) );
NAND3X1 NAND3X1_33 ( .A(_470_), .B(_472_), .C(_471_), .Y(_473_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_467_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_468_) );
OAI21X1 OAI21X1_89 ( .A(_467_), .B(_468_), .C(1'b0), .Y(_469_) );
NAND2X1 NAND2X1_90 ( .A(_469_), .B(_473_), .Y(_39__0_) );
OAI21X1 OAI21X1_90 ( .A(_470_), .B(_467_), .C(_472_), .Y(_41__1_) );
INVX1 INVX1_58 ( .A(_41__3_), .Y(_477_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_478_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_479_) );
NAND3X1 NAND3X1_34 ( .A(_477_), .B(_479_), .C(_478_), .Y(_480_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_474_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_475_) );
OAI21X1 OAI21X1_91 ( .A(_474_), .B(_475_), .C(_41__3_), .Y(_476_) );
NAND2X1 NAND2X1_92 ( .A(_476_), .B(_480_), .Y(_39__3_) );
OAI21X1 OAI21X1_92 ( .A(_477_), .B(_474_), .C(_479_), .Y(_37_) );
INVX1 INVX1_59 ( .A(_41__1_), .Y(_484_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_485_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_486_) );
NAND3X1 NAND3X1_35 ( .A(_484_), .B(_486_), .C(_485_), .Y(_487_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_481_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_482_) );
OAI21X1 OAI21X1_93 ( .A(_481_), .B(_482_), .C(_41__1_), .Y(_483_) );
NAND2X1 NAND2X1_94 ( .A(_483_), .B(_487_), .Y(_39__1_) );
OAI21X1 OAI21X1_94 ( .A(_484_), .B(_481_), .C(_486_), .Y(_41__2_) );
INVX1 INVX1_60 ( .A(_41__2_), .Y(_491_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_492_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_493_) );
NAND3X1 NAND3X1_36 ( .A(_491_), .B(_493_), .C(_492_), .Y(_494_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_488_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_489_) );
OAI21X1 OAI21X1_95 ( .A(_488_), .B(_489_), .C(_41__2_), .Y(_490_) );
NAND2X1 NAND2X1_96 ( .A(_490_), .B(_494_), .Y(_39__2_) );
OAI21X1 OAI21X1_96 ( .A(_491_), .B(_488_), .C(_493_), .Y(_41__3_) );
INVX1 INVX1_61 ( .A(1'b1), .Y(_498_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_499_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_500_) );
NAND3X1 NAND3X1_37 ( .A(_498_), .B(_500_), .C(_499_), .Y(_501_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_495_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_496_) );
OAI21X1 OAI21X1_97 ( .A(_495_), .B(_496_), .C(1'b1), .Y(_497_) );
NAND2X1 NAND2X1_98 ( .A(_497_), .B(_501_), .Y(_40__0_) );
OAI21X1 OAI21X1_98 ( .A(_498_), .B(_495_), .C(_500_), .Y(_42__1_) );
INVX1 INVX1_62 ( .A(_42__3_), .Y(_505_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_506_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_507_) );
NAND3X1 NAND3X1_38 ( .A(_505_), .B(_507_), .C(_506_), .Y(_508_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_502_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_503_) );
OAI21X1 OAI21X1_99 ( .A(_502_), .B(_503_), .C(_42__3_), .Y(_504_) );
NAND2X1 NAND2X1_100 ( .A(_504_), .B(_508_), .Y(_40__3_) );
OAI21X1 OAI21X1_100 ( .A(_505_), .B(_502_), .C(_507_), .Y(_38_) );
INVX1 INVX1_63 ( .A(_42__1_), .Y(_512_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_513_) );
NAND2X1 NAND2X1_101 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_514_) );
NAND3X1 NAND3X1_39 ( .A(_512_), .B(_514_), .C(_513_), .Y(_515_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_509_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_510_) );
OAI21X1 OAI21X1_101 ( .A(_509_), .B(_510_), .C(_42__1_), .Y(_511_) );
NAND2X1 NAND2X1_102 ( .A(_511_), .B(_515_), .Y(_40__1_) );
OAI21X1 OAI21X1_102 ( .A(_512_), .B(_509_), .C(_514_), .Y(_42__2_) );
INVX1 INVX1_64 ( .A(_42__2_), .Y(_519_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_520_) );
NAND2X1 NAND2X1_103 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_521_) );
NAND3X1 NAND3X1_40 ( .A(_519_), .B(_521_), .C(_520_), .Y(_522_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_516_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_517_) );
OAI21X1 OAI21X1_103 ( .A(_516_), .B(_517_), .C(_42__2_), .Y(_518_) );
NAND2X1 NAND2X1_104 ( .A(_518_), .B(_522_), .Y(_40__2_) );
OAI21X1 OAI21X1_104 ( .A(_519_), .B(_516_), .C(_521_), .Y(_42__3_) );
INVX1 INVX1_65 ( .A(_43_), .Y(_523_) );
NAND2X1 NAND2X1_105 ( .A(_44_), .B(w_cout_7_), .Y(_524_) );
OAI21X1 OAI21X1_105 ( .A(w_cout_7_), .B(_523_), .C(_524_), .Y(w_cout_8_) );
INVX1 INVX1_66 ( .A(_45__0_), .Y(_525_) );
NAND2X1 NAND2X1_106 ( .A(_46__0_), .B(w_cout_7_), .Y(_526_) );
OAI21X1 OAI21X1_106 ( .A(w_cout_7_), .B(_525_), .C(_526_), .Y(_0__32_) );
INVX1 INVX1_67 ( .A(_45__1_), .Y(_527_) );
NAND2X1 NAND2X1_107 ( .A(w_cout_7_), .B(_46__1_), .Y(_528_) );
OAI21X1 OAI21X1_107 ( .A(w_cout_7_), .B(_527_), .C(_528_), .Y(_0__33_) );
INVX1 INVX1_68 ( .A(_45__2_), .Y(_529_) );
NAND2X1 NAND2X1_108 ( .A(w_cout_7_), .B(_46__2_), .Y(_530_) );
OAI21X1 OAI21X1_108 ( .A(w_cout_7_), .B(_529_), .C(_530_), .Y(_0__34_) );
INVX1 INVX1_69 ( .A(_45__3_), .Y(_531_) );
NAND2X1 NAND2X1_109 ( .A(w_cout_7_), .B(_46__3_), .Y(_532_) );
OAI21X1 OAI21X1_109 ( .A(w_cout_7_), .B(_531_), .C(_532_), .Y(_0__35_) );
INVX1 INVX1_70 ( .A(1'b0), .Y(_536_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_537_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_538_) );
NAND3X1 NAND3X1_41 ( .A(_536_), .B(_538_), .C(_537_), .Y(_539_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_533_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_534_) );
OAI21X1 OAI21X1_110 ( .A(_533_), .B(_534_), .C(1'b0), .Y(_535_) );
NAND2X1 NAND2X1_111 ( .A(_535_), .B(_539_), .Y(_45__0_) );
OAI21X1 OAI21X1_111 ( .A(_536_), .B(_533_), .C(_538_), .Y(_47__1_) );
INVX1 INVX1_71 ( .A(_47__3_), .Y(_543_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_544_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_545_) );
NAND3X1 NAND3X1_42 ( .A(_543_), .B(_545_), .C(_544_), .Y(_546_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_540_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_541_) );
OAI21X1 OAI21X1_112 ( .A(_540_), .B(_541_), .C(_47__3_), .Y(_542_) );
NAND2X1 NAND2X1_113 ( .A(_542_), .B(_546_), .Y(_45__3_) );
OAI21X1 OAI21X1_113 ( .A(_543_), .B(_540_), .C(_545_), .Y(_43_) );
INVX1 INVX1_72 ( .A(_47__1_), .Y(_550_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_551_) );
NAND2X1 NAND2X1_114 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_552_) );
NAND3X1 NAND3X1_43 ( .A(_550_), .B(_552_), .C(_551_), .Y(_553_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_547_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_548_) );
OAI21X1 OAI21X1_114 ( .A(_547_), .B(_548_), .C(_47__1_), .Y(_549_) );
NAND2X1 NAND2X1_115 ( .A(_549_), .B(_553_), .Y(_45__1_) );
OAI21X1 OAI21X1_115 ( .A(_550_), .B(_547_), .C(_552_), .Y(_47__2_) );
INVX1 INVX1_73 ( .A(_47__2_), .Y(_557_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_558_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_559_) );
NAND3X1 NAND3X1_44 ( .A(_557_), .B(_559_), .C(_558_), .Y(_560_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_554_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_555_) );
OAI21X1 OAI21X1_116 ( .A(_554_), .B(_555_), .C(_47__2_), .Y(_556_) );
NAND2X1 NAND2X1_117 ( .A(_556_), .B(_560_), .Y(_45__2_) );
OAI21X1 OAI21X1_117 ( .A(_557_), .B(_554_), .C(_559_), .Y(_47__3_) );
INVX1 INVX1_74 ( .A(1'b1), .Y(_564_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_565_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_566_) );
NAND3X1 NAND3X1_45 ( .A(_564_), .B(_566_), .C(_565_), .Y(_567_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_561_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_562_) );
OAI21X1 OAI21X1_118 ( .A(_561_), .B(_562_), .C(1'b1), .Y(_563_) );
NAND2X1 NAND2X1_119 ( .A(_563_), .B(_567_), .Y(_46__0_) );
OAI21X1 OAI21X1_119 ( .A(_564_), .B(_561_), .C(_566_), .Y(_48__1_) );
INVX1 INVX1_75 ( .A(_48__3_), .Y(_571_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_572_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_573_) );
NAND3X1 NAND3X1_46 ( .A(_571_), .B(_573_), .C(_572_), .Y(_574_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_568_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_569_) );
OAI21X1 OAI21X1_120 ( .A(_568_), .B(_569_), .C(_48__3_), .Y(_570_) );
NAND2X1 NAND2X1_121 ( .A(_570_), .B(_574_), .Y(_46__3_) );
OAI21X1 OAI21X1_121 ( .A(_571_), .B(_568_), .C(_573_), .Y(_44_) );
INVX1 INVX1_76 ( .A(_48__1_), .Y(_578_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_579_) );
NAND2X1 NAND2X1_122 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_580_) );
NAND3X1 NAND3X1_47 ( .A(_578_), .B(_580_), .C(_579_), .Y(_581_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_575_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_576_) );
OAI21X1 OAI21X1_122 ( .A(_575_), .B(_576_), .C(_48__1_), .Y(_577_) );
NAND2X1 NAND2X1_123 ( .A(_577_), .B(_581_), .Y(_46__1_) );
OAI21X1 OAI21X1_123 ( .A(_578_), .B(_575_), .C(_580_), .Y(_48__2_) );
INVX1 INVX1_77 ( .A(_48__2_), .Y(_585_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_586_) );
NAND2X1 NAND2X1_124 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_587_) );
NAND3X1 NAND3X1_48 ( .A(_585_), .B(_587_), .C(_586_), .Y(_588_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_582_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_583_) );
OAI21X1 OAI21X1_124 ( .A(_582_), .B(_583_), .C(_48__2_), .Y(_584_) );
NAND2X1 NAND2X1_125 ( .A(_584_), .B(_588_), .Y(_46__2_) );
OAI21X1 OAI21X1_125 ( .A(_585_), .B(_582_), .C(_587_), .Y(_48__3_) );
INVX1 INVX1_78 ( .A(_49_), .Y(_589_) );
NAND2X1 NAND2X1_126 ( .A(_50_), .B(w_cout_8_), .Y(_590_) );
OAI21X1 OAI21X1_126 ( .A(w_cout_8_), .B(_589_), .C(_590_), .Y(w_cout_9_) );
INVX1 INVX1_79 ( .A(_51__0_), .Y(_591_) );
NAND2X1 NAND2X1_127 ( .A(_52__0_), .B(w_cout_8_), .Y(_592_) );
OAI21X1 OAI21X1_127 ( .A(w_cout_8_), .B(_591_), .C(_592_), .Y(_0__36_) );
INVX1 INVX1_80 ( .A(_51__1_), .Y(_593_) );
NAND2X1 NAND2X1_128 ( .A(w_cout_8_), .B(_52__1_), .Y(_594_) );
OAI21X1 OAI21X1_128 ( .A(w_cout_8_), .B(_593_), .C(_594_), .Y(_0__37_) );
INVX1 INVX1_81 ( .A(_51__2_), .Y(_595_) );
NAND2X1 NAND2X1_129 ( .A(w_cout_8_), .B(_52__2_), .Y(_596_) );
OAI21X1 OAI21X1_129 ( .A(w_cout_8_), .B(_595_), .C(_596_), .Y(_0__38_) );
INVX1 INVX1_82 ( .A(_51__3_), .Y(_597_) );
NAND2X1 NAND2X1_130 ( .A(w_cout_8_), .B(_52__3_), .Y(_598_) );
OAI21X1 OAI21X1_130 ( .A(w_cout_8_), .B(_597_), .C(_598_), .Y(_0__39_) );
INVX1 INVX1_83 ( .A(1'b0), .Y(_602_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_603_) );
NAND2X1 NAND2X1_131 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_604_) );
NAND3X1 NAND3X1_49 ( .A(_602_), .B(_604_), .C(_603_), .Y(_605_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_599_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_600_) );
OAI21X1 OAI21X1_131 ( .A(_599_), .B(_600_), .C(1'b0), .Y(_601_) );
NAND2X1 NAND2X1_132 ( .A(_601_), .B(_605_), .Y(_51__0_) );
OAI21X1 OAI21X1_132 ( .A(_602_), .B(_599_), .C(_604_), .Y(_53__1_) );
INVX1 INVX1_84 ( .A(_53__3_), .Y(_609_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_610_) );
NAND2X1 NAND2X1_133 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_611_) );
NAND3X1 NAND3X1_50 ( .A(_609_), .B(_611_), .C(_610_), .Y(_612_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_606_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_607_) );
OAI21X1 OAI21X1_133 ( .A(_606_), .B(_607_), .C(_53__3_), .Y(_608_) );
NAND2X1 NAND2X1_134 ( .A(_608_), .B(_612_), .Y(_51__3_) );
OAI21X1 OAI21X1_134 ( .A(_609_), .B(_606_), .C(_611_), .Y(_49_) );
INVX1 INVX1_85 ( .A(_53__1_), .Y(_616_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_617_) );
NAND2X1 NAND2X1_135 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_618_) );
NAND3X1 NAND3X1_51 ( .A(_616_), .B(_618_), .C(_617_), .Y(_619_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_613_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_614_) );
OAI21X1 OAI21X1_135 ( .A(_613_), .B(_614_), .C(_53__1_), .Y(_615_) );
NAND2X1 NAND2X1_136 ( .A(_615_), .B(_619_), .Y(_51__1_) );
OAI21X1 OAI21X1_136 ( .A(_616_), .B(_613_), .C(_618_), .Y(_53__2_) );
INVX1 INVX1_86 ( .A(_53__2_), .Y(_623_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_624_) );
NAND2X1 NAND2X1_137 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_625_) );
NAND3X1 NAND3X1_52 ( .A(_623_), .B(_625_), .C(_624_), .Y(_626_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_620_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_621_) );
OAI21X1 OAI21X1_137 ( .A(_620_), .B(_621_), .C(_53__2_), .Y(_622_) );
NAND2X1 NAND2X1_138 ( .A(_622_), .B(_626_), .Y(_51__2_) );
OAI21X1 OAI21X1_138 ( .A(_623_), .B(_620_), .C(_625_), .Y(_53__3_) );
INVX1 INVX1_87 ( .A(1'b1), .Y(_630_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_631_) );
NAND2X1 NAND2X1_139 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_632_) );
NAND3X1 NAND3X1_53 ( .A(_630_), .B(_632_), .C(_631_), .Y(_633_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_627_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_628_) );
OAI21X1 OAI21X1_139 ( .A(_627_), .B(_628_), .C(1'b1), .Y(_629_) );
NAND2X1 NAND2X1_140 ( .A(_629_), .B(_633_), .Y(_52__0_) );
OAI21X1 OAI21X1_140 ( .A(_630_), .B(_627_), .C(_632_), .Y(_54__1_) );
INVX1 INVX1_88 ( .A(_54__3_), .Y(_637_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_638_) );
NAND2X1 NAND2X1_141 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_639_) );
NAND3X1 NAND3X1_54 ( .A(_637_), .B(_639_), .C(_638_), .Y(_640_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_634_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_635_) );
OAI21X1 OAI21X1_141 ( .A(_634_), .B(_635_), .C(_54__3_), .Y(_636_) );
NAND2X1 NAND2X1_142 ( .A(_636_), .B(_640_), .Y(_52__3_) );
OAI21X1 OAI21X1_142 ( .A(_637_), .B(_634_), .C(_639_), .Y(_50_) );
INVX1 INVX1_89 ( .A(_54__1_), .Y(_644_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_645_) );
NAND2X1 NAND2X1_143 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_646_) );
NAND3X1 NAND3X1_55 ( .A(_644_), .B(_646_), .C(_645_), .Y(_647_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_641_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_642_) );
OAI21X1 OAI21X1_143 ( .A(_641_), .B(_642_), .C(_54__1_), .Y(_643_) );
NAND2X1 NAND2X1_144 ( .A(_643_), .B(_647_), .Y(_52__1_) );
OAI21X1 OAI21X1_144 ( .A(_644_), .B(_641_), .C(_646_), .Y(_54__2_) );
INVX1 INVX1_90 ( .A(_54__2_), .Y(_651_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_652_) );
NAND2X1 NAND2X1_145 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_653_) );
NAND3X1 NAND3X1_56 ( .A(_651_), .B(_653_), .C(_652_), .Y(_654_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_648_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_649_) );
OAI21X1 OAI21X1_145 ( .A(_648_), .B(_649_), .C(_54__2_), .Y(_650_) );
NAND2X1 NAND2X1_146 ( .A(_650_), .B(_654_), .Y(_52__2_) );
OAI21X1 OAI21X1_146 ( .A(_651_), .B(_648_), .C(_653_), .Y(_54__3_) );
INVX1 INVX1_91 ( .A(_55_), .Y(_655_) );
NAND2X1 NAND2X1_147 ( .A(_56_), .B(w_cout_9_), .Y(_656_) );
OAI21X1 OAI21X1_147 ( .A(w_cout_9_), .B(_655_), .C(_656_), .Y(csa_inst_cin) );
INVX1 INVX1_92 ( .A(_57__0_), .Y(_657_) );
NAND2X1 NAND2X1_148 ( .A(_58__0_), .B(w_cout_9_), .Y(_658_) );
OAI21X1 OAI21X1_148 ( .A(w_cout_9_), .B(_657_), .C(_658_), .Y(_0__40_) );
INVX1 INVX1_93 ( .A(_57__1_), .Y(_659_) );
NAND2X1 NAND2X1_149 ( .A(w_cout_9_), .B(_58__1_), .Y(_660_) );
OAI21X1 OAI21X1_149 ( .A(w_cout_9_), .B(_659_), .C(_660_), .Y(_0__41_) );
INVX1 INVX1_94 ( .A(_57__2_), .Y(_661_) );
NAND2X1 NAND2X1_150 ( .A(w_cout_9_), .B(_58__2_), .Y(_662_) );
OAI21X1 OAI21X1_150 ( .A(w_cout_9_), .B(_661_), .C(_662_), .Y(_0__42_) );
INVX1 INVX1_95 ( .A(_57__3_), .Y(_663_) );
NAND2X1 NAND2X1_151 ( .A(w_cout_9_), .B(_58__3_), .Y(_664_) );
OAI21X1 OAI21X1_151 ( .A(w_cout_9_), .B(_663_), .C(_664_), .Y(_0__43_) );
INVX1 INVX1_96 ( .A(1'b0), .Y(_668_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_669_) );
NAND2X1 NAND2X1_152 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_670_) );
NAND3X1 NAND3X1_57 ( .A(_668_), .B(_670_), .C(_669_), .Y(_671_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_665_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_666_) );
OAI21X1 OAI21X1_152 ( .A(_665_), .B(_666_), .C(1'b0), .Y(_667_) );
NAND2X1 NAND2X1_153 ( .A(_667_), .B(_671_), .Y(_57__0_) );
OAI21X1 OAI21X1_153 ( .A(_668_), .B(_665_), .C(_670_), .Y(_59__1_) );
INVX1 INVX1_97 ( .A(_59__3_), .Y(_675_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_676_) );
NAND2X1 NAND2X1_154 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_677_) );
NAND3X1 NAND3X1_58 ( .A(_675_), .B(_677_), .C(_676_), .Y(_678_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_672_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_673_) );
OAI21X1 OAI21X1_154 ( .A(_672_), .B(_673_), .C(_59__3_), .Y(_674_) );
NAND2X1 NAND2X1_155 ( .A(_674_), .B(_678_), .Y(_57__3_) );
OAI21X1 OAI21X1_155 ( .A(_675_), .B(_672_), .C(_677_), .Y(_55_) );
INVX1 INVX1_98 ( .A(_59__1_), .Y(_682_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_683_) );
NAND2X1 NAND2X1_156 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_684_) );
NAND3X1 NAND3X1_59 ( .A(_682_), .B(_684_), .C(_683_), .Y(_685_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_679_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_680_) );
OAI21X1 OAI21X1_156 ( .A(_679_), .B(_680_), .C(_59__1_), .Y(_681_) );
NAND2X1 NAND2X1_157 ( .A(_681_), .B(_685_), .Y(_57__1_) );
OAI21X1 OAI21X1_157 ( .A(_682_), .B(_679_), .C(_684_), .Y(_59__2_) );
INVX1 INVX1_99 ( .A(_59__2_), .Y(_689_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_690_) );
NAND2X1 NAND2X1_158 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_691_) );
NAND3X1 NAND3X1_60 ( .A(_689_), .B(_691_), .C(_690_), .Y(_692_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_686_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_687_) );
OAI21X1 OAI21X1_158 ( .A(_686_), .B(_687_), .C(_59__2_), .Y(_688_) );
NAND2X1 NAND2X1_159 ( .A(_688_), .B(_692_), .Y(_57__2_) );
OAI21X1 OAI21X1_159 ( .A(_689_), .B(_686_), .C(_691_), .Y(_59__3_) );
INVX1 INVX1_100 ( .A(1'b1), .Y(_696_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_697_) );
NAND2X1 NAND2X1_160 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_698_) );
NAND3X1 NAND3X1_61 ( .A(_696_), .B(_698_), .C(_697_), .Y(_699_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_693_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_694_) );
OAI21X1 OAI21X1_160 ( .A(_693_), .B(_694_), .C(1'b1), .Y(_695_) );
NAND2X1 NAND2X1_161 ( .A(_695_), .B(_699_), .Y(_58__0_) );
OAI21X1 OAI21X1_161 ( .A(_696_), .B(_693_), .C(_698_), .Y(_60__1_) );
INVX1 INVX1_101 ( .A(_60__3_), .Y(_703_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_704_) );
NAND2X1 NAND2X1_162 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_705_) );
NAND3X1 NAND3X1_62 ( .A(_703_), .B(_705_), .C(_704_), .Y(_706_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_700_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_701_) );
OAI21X1 OAI21X1_162 ( .A(_700_), .B(_701_), .C(_60__3_), .Y(_702_) );
NAND2X1 NAND2X1_163 ( .A(_702_), .B(_706_), .Y(_58__3_) );
OAI21X1 OAI21X1_163 ( .A(_703_), .B(_700_), .C(_705_), .Y(_56_) );
INVX1 INVX1_102 ( .A(_60__1_), .Y(_710_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_711_) );
NAND2X1 NAND2X1_164 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_712_) );
NAND3X1 NAND3X1_63 ( .A(_710_), .B(_712_), .C(_711_), .Y(_713_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_707_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_708_) );
OAI21X1 OAI21X1_164 ( .A(_707_), .B(_708_), .C(_60__1_), .Y(_709_) );
NAND2X1 NAND2X1_165 ( .A(_709_), .B(_713_), .Y(_58__1_) );
OAI21X1 OAI21X1_165 ( .A(_710_), .B(_707_), .C(_712_), .Y(_60__2_) );
INVX1 INVX1_103 ( .A(_60__2_), .Y(_717_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_718_) );
NAND2X1 NAND2X1_166 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_719_) );
NAND3X1 NAND3X1_64 ( .A(_717_), .B(_719_), .C(_718_), .Y(_720_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_714_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_715_) );
OAI21X1 OAI21X1_166 ( .A(_714_), .B(_715_), .C(_60__2_), .Y(_716_) );
NAND2X1 NAND2X1_167 ( .A(_716_), .B(_720_), .Y(_58__2_) );
OAI21X1 OAI21X1_167 ( .A(_717_), .B(_714_), .C(_719_), .Y(_60__3_) );
INVX1 INVX1_104 ( .A(csa_inst_cout0_0), .Y(_721_) );
NAND2X1 NAND2X1_168 ( .A(csa_inst_cout0_1), .B(csa_inst_cin), .Y(_722_) );
OAI21X1 OAI21X1_168 ( .A(csa_inst_cin), .B(_721_), .C(_722_), .Y(w_cout_11_) );
INVX1 INVX1_105 ( .A(1'b0), .Y(_724_) );
NAND2X1 NAND2X1_169 ( .A(1'b0), .B(1'b0), .Y(_725_) );
NOR2X1 NOR2X1_65 ( .A(1'b0), .B(1'b0), .Y(_723_) );
OAI21X1 OAI21X1_169 ( .A(_724_), .B(_723_), .C(_725_), .Y(csa_inst_rca0_0_fa0_o_carry) );
INVX1 INVX1_106 ( .A(csa_inst_rca0_0_fa31_i_carry), .Y(_727_) );
NAND2X1 NAND2X1_170 ( .A(1'b0), .B(1'b0), .Y(_728_) );
NOR2X1 NOR2X1_66 ( .A(1'b0), .B(1'b0), .Y(_726_) );
OAI21X1 OAI21X1_170 ( .A(_727_), .B(_726_), .C(_728_), .Y(csa_inst_cout0_0) );
INVX1 INVX1_107 ( .A(csa_inst_rca0_0_fa0_o_carry), .Y(_730_) );
NAND2X1 NAND2X1_171 ( .A(1'b0), .B(1'b0), .Y(_731_) );
NOR2X1 NOR2X1_67 ( .A(1'b0), .B(1'b0), .Y(_729_) );
OAI21X1 OAI21X1_171 ( .A(_730_), .B(_729_), .C(_731_), .Y(csa_inst_rca0_0_fa_1__o_carry) );
INVX1 INVX1_108 ( .A(csa_inst_rca0_0_fa_1__o_carry), .Y(_733_) );
NAND2X1 NAND2X1_172 ( .A(1'b0), .B(1'b0), .Y(_734_) );
NOR2X1 NOR2X1_68 ( .A(1'b0), .B(1'b0), .Y(_732_) );
OAI21X1 OAI21X1_172 ( .A(_733_), .B(_732_), .C(_734_), .Y(csa_inst_rca0_0_fa31_i_carry) );
INVX1 INVX1_109 ( .A(1'b1), .Y(_736_) );
NAND2X1 NAND2X1_173 ( .A(1'b0), .B(1'b0), .Y(_737_) );
NOR2X1 NOR2X1_69 ( .A(1'b0), .B(1'b0), .Y(_735_) );
OAI21X1 OAI21X1_173 ( .A(_736_), .B(_735_), .C(_737_), .Y(csa_inst_rca0_1_fa0_o_carry) );
INVX1 INVX1_110 ( .A(csa_inst_rca0_1_fa31_i_carry), .Y(_739_) );
NAND2X1 NAND2X1_174 ( .A(1'b0), .B(1'b0), .Y(_740_) );
NOR2X1 NOR2X1_70 ( .A(1'b0), .B(1'b0), .Y(_738_) );
OAI21X1 OAI21X1_174 ( .A(_739_), .B(_738_), .C(_740_), .Y(csa_inst_cout0_1) );
INVX1 INVX1_111 ( .A(csa_inst_rca0_1_fa0_o_carry), .Y(_742_) );
NAND2X1 NAND2X1_175 ( .A(1'b0), .B(1'b0), .Y(_743_) );
NOR2X1 NOR2X1_71 ( .A(1'b0), .B(1'b0), .Y(_741_) );
OAI21X1 OAI21X1_175 ( .A(_742_), .B(_741_), .C(_743_), .Y(csa_inst_rca0_1_fa_1__o_carry) );
INVX1 INVX1_112 ( .A(csa_inst_rca0_1_fa_1__o_carry), .Y(_745_) );
NAND2X1 NAND2X1_176 ( .A(1'b0), .B(1'b0), .Y(_746_) );
NOR2X1 NOR2X1_72 ( .A(1'b0), .B(1'b0), .Y(_744_) );
OAI21X1 OAI21X1_176 ( .A(_745_), .B(_744_), .C(_746_), .Y(csa_inst_rca0_1_fa31_i_carry) );
INVX1 INVX1_113 ( .A(1'b0), .Y(_750_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_751_) );
NAND2X1 NAND2X1_177 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_752_) );
NAND3X1 NAND3X1_65 ( .A(_750_), .B(_752_), .C(_751_), .Y(_753_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_747_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_748_) );
OAI21X1 OAI21X1_177 ( .A(_747_), .B(_748_), .C(1'b0), .Y(_749_) );
NAND2X1 NAND2X1_178 ( .A(_749_), .B(_753_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_178 ( .A(_750_), .B(_747_), .C(_752_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_114 ( .A(rca_inst_fa31_i_carry), .Y(_757_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_758_) );
NAND2X1 NAND2X1_179 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_759_) );
NAND3X1 NAND3X1_66 ( .A(_757_), .B(_759_), .C(_758_), .Y(_760_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_754_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_755_) );
OAI21X1 OAI21X1_179 ( .A(_754_), .B(_755_), .C(rca_inst_fa31_i_carry), .Y(_756_) );
NAND2X1 NAND2X1_180 ( .A(_756_), .B(_760_), .Y(rca_inst_fa31_o_sum) );
OAI21X1 OAI21X1_180 ( .A(_757_), .B(_754_), .C(_759_), .Y(rca_inst_cout) );
INVX1 INVX1_115 ( .A(rca_inst_fa0_o_carry), .Y(_764_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_765_) );
NAND2X1 NAND2X1_181 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_766_) );
NAND3X1 NAND3X1_67 ( .A(_764_), .B(_766_), .C(_765_), .Y(_767_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_761_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_762_) );
OAI21X1 OAI21X1_181 ( .A(_761_), .B(_762_), .C(rca_inst_fa0_o_carry), .Y(_763_) );
NAND2X1 NAND2X1_182 ( .A(_763_), .B(_767_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_182 ( .A(_764_), .B(_761_), .C(_766_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_116 ( .A(rca_inst_fa_1__o_carry), .Y(_771_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_772_) );
NAND2X1 NAND2X1_183 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_773_) );
NAND3X1 NAND3X1_68 ( .A(_771_), .B(_773_), .C(_772_), .Y(_774_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_768_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_769_) );
OAI21X1 OAI21X1_183 ( .A(_768_), .B(_769_), .C(rca_inst_fa_1__o_carry), .Y(_770_) );
NAND2X1 NAND2X1_184 ( .A(_770_), .B(_774_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_184 ( .A(_771_), .B(_768_), .C(_773_), .Y(rca_inst_fa31_i_carry) );
BUFX2 BUFX2_1 ( .A(w_cout_11_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa31_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(1'b0), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(1'b0), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(1'b0), .Y(sum[46]) );
INVX1 INVX1_117 ( .A(_1_), .Y(_61_) );
NAND2X1 NAND2X1_185 ( .A(_2_), .B(rca_inst_cout), .Y(_62_) );
OAI21X1 OAI21X1_185 ( .A(rca_inst_cout), .B(_61_), .C(_62_), .Y(w_cout_1_) );
INVX1 INVX1_118 ( .A(_3__0_), .Y(_63_) );
NAND2X1 NAND2X1_186 ( .A(_4__0_), .B(rca_inst_cout), .Y(_64_) );
OAI21X1 OAI21X1_186 ( .A(rca_inst_cout), .B(_63_), .C(_64_), .Y(_0__4_) );
INVX1 INVX1_119 ( .A(_3__1_), .Y(_65_) );
NAND2X1 NAND2X1_187 ( .A(rca_inst_cout), .B(_4__1_), .Y(_66_) );
OAI21X1 OAI21X1_187 ( .A(rca_inst_cout), .B(_65_), .C(_66_), .Y(_0__5_) );
INVX1 INVX1_120 ( .A(_3__2_), .Y(_67_) );
NAND2X1 NAND2X1_188 ( .A(rca_inst_cout), .B(_4__2_), .Y(_68_) );
OAI21X1 OAI21X1_188 ( .A(rca_inst_cout), .B(_67_), .C(_68_), .Y(_0__6_) );
INVX1 INVX1_121 ( .A(_3__3_), .Y(_69_) );
NAND2X1 NAND2X1_189 ( .A(rca_inst_cout), .B(_4__3_), .Y(_70_) );
OAI21X1 OAI21X1_189 ( .A(rca_inst_cout), .B(_69_), .C(_70_), .Y(_0__7_) );
INVX1 INVX1_122 ( .A(1'b0), .Y(_74_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_75_) );
NAND2X1 NAND2X1_190 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_76_) );
NAND3X1 NAND3X1_69 ( .A(_74_), .B(_76_), .C(_75_), .Y(_77_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_71_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_72_) );
OAI21X1 OAI21X1_190 ( .A(_71_), .B(_72_), .C(1'b0), .Y(_73_) );
NAND2X1 NAND2X1_191 ( .A(_73_), .B(_77_), .Y(_3__0_) );
OAI21X1 OAI21X1_191 ( .A(_74_), .B(_71_), .C(_76_), .Y(_5__1_) );
INVX1 INVX1_123 ( .A(_5__3_), .Y(_81_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_82_) );
NAND2X1 NAND2X1_192 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_83_) );
NAND3X1 NAND3X1_70 ( .A(_81_), .B(_83_), .C(_82_), .Y(_84_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_78_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_79_) );
OAI21X1 OAI21X1_192 ( .A(_78_), .B(_79_), .C(_5__3_), .Y(_80_) );
NAND2X1 NAND2X1_193 ( .A(_80_), .B(_84_), .Y(_3__3_) );
OAI21X1 OAI21X1_193 ( .A(_81_), .B(_78_), .C(_83_), .Y(_1_) );
INVX1 INVX1_124 ( .A(_5__1_), .Y(_88_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_89_) );
NAND2X1 NAND2X1_194 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_90_) );
NAND3X1 NAND3X1_71 ( .A(_88_), .B(_90_), .C(_89_), .Y(_91_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_85_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_86_) );
OAI21X1 OAI21X1_194 ( .A(_85_), .B(_86_), .C(_5__1_), .Y(_87_) );
NAND2X1 NAND2X1_195 ( .A(_87_), .B(_91_), .Y(_3__1_) );
OAI21X1 OAI21X1_195 ( .A(_88_), .B(_85_), .C(_90_), .Y(_5__2_) );
INVX1 INVX1_125 ( .A(_5__2_), .Y(_95_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_96_) );
NAND2X1 NAND2X1_196 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_97_) );
NAND3X1 NAND3X1_72 ( .A(_95_), .B(_97_), .C(_96_), .Y(_98_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_92_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_93_) );
OAI21X1 OAI21X1_196 ( .A(_92_), .B(_93_), .C(_5__2_), .Y(_94_) );
NAND2X1 NAND2X1_197 ( .A(_94_), .B(_98_), .Y(_3__2_) );
OAI21X1 OAI21X1_197 ( .A(_95_), .B(_92_), .C(_97_), .Y(_5__3_) );
INVX1 INVX1_126 ( .A(1'b1), .Y(_102_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_103_) );
NAND2X1 NAND2X1_198 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_104_) );
NAND3X1 NAND3X1_73 ( .A(_102_), .B(_104_), .C(_103_), .Y(_105_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_99_) );
AND2X2 AND2X2_73 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_100_) );
OAI21X1 OAI21X1_198 ( .A(_99_), .B(_100_), .C(1'b1), .Y(_101_) );
NAND2X1 NAND2X1_199 ( .A(_101_), .B(_105_), .Y(_4__0_) );
OAI21X1 OAI21X1_199 ( .A(_102_), .B(_99_), .C(_104_), .Y(_6__1_) );
INVX1 INVX1_127 ( .A(_6__3_), .Y(_109_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_110_) );
NAND2X1 NAND2X1_200 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_111_) );
NAND3X1 NAND3X1_74 ( .A(_109_), .B(_111_), .C(_110_), .Y(_112_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_106_) );
AND2X2 AND2X2_74 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_107_) );
OAI21X1 OAI21X1_200 ( .A(_106_), .B(_107_), .C(_6__3_), .Y(_108_) );
NAND2X1 NAND2X1_201 ( .A(_108_), .B(_112_), .Y(_4__3_) );
OAI21X1 OAI21X1_201 ( .A(_109_), .B(_106_), .C(_111_), .Y(_2_) );
INVX1 INVX1_128 ( .A(_6__1_), .Y(_116_) );
OR2X2 OR2X2_75 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_117_) );
NAND2X1 NAND2X1_202 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_118_) );
NAND3X1 NAND3X1_75 ( .A(_116_), .B(_118_), .C(_117_), .Y(_119_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_113_) );
AND2X2 AND2X2_75 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_114_) );
OAI21X1 OAI21X1_202 ( .A(_113_), .B(_114_), .C(_6__1_), .Y(_115_) );
NAND2X1 NAND2X1_203 ( .A(_115_), .B(_119_), .Y(_4__1_) );
OAI21X1 OAI21X1_203 ( .A(_116_), .B(_113_), .C(_118_), .Y(_6__2_) );
INVX1 INVX1_129 ( .A(_6__2_), .Y(_123_) );
OR2X2 OR2X2_76 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_124_) );
NAND2X1 NAND2X1_204 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_125_) );
NAND3X1 NAND3X1_76 ( .A(_123_), .B(_125_), .C(_124_), .Y(_126_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_120_) );
AND2X2 AND2X2_76 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_121_) );
OAI21X1 OAI21X1_204 ( .A(_120_), .B(_121_), .C(_6__2_), .Y(_122_) );
NAND2X1 NAND2X1_205 ( .A(_122_), .B(_126_), .Y(_4__2_) );
OAI21X1 OAI21X1_205 ( .A(_123_), .B(_120_), .C(_125_), .Y(_6__3_) );
INVX1 INVX1_130 ( .A(_7_), .Y(_127_) );
NAND2X1 NAND2X1_206 ( .A(_8_), .B(w_cout_1_), .Y(_128_) );
OAI21X1 OAI21X1_206 ( .A(w_cout_1_), .B(_127_), .C(_128_), .Y(w_cout_2_) );
INVX1 INVX1_131 ( .A(_9__0_), .Y(_129_) );
NAND2X1 NAND2X1_207 ( .A(_10__0_), .B(w_cout_1_), .Y(_130_) );
OAI21X1 OAI21X1_207 ( .A(w_cout_1_), .B(_129_), .C(_130_), .Y(_0__8_) );
INVX1 INVX1_132 ( .A(_9__1_), .Y(_131_) );
NAND2X1 NAND2X1_208 ( .A(w_cout_1_), .B(_10__1_), .Y(_132_) );
OAI21X1 OAI21X1_208 ( .A(w_cout_1_), .B(_131_), .C(_132_), .Y(_0__9_) );
INVX1 INVX1_133 ( .A(_9__2_), .Y(_133_) );
NAND2X1 NAND2X1_209 ( .A(w_cout_1_), .B(_10__2_), .Y(_134_) );
OAI21X1 OAI21X1_209 ( .A(w_cout_1_), .B(_133_), .C(_134_), .Y(_0__10_) );
INVX1 INVX1_134 ( .A(_9__3_), .Y(_135_) );
NAND2X1 NAND2X1_210 ( .A(w_cout_1_), .B(_10__3_), .Y(_136_) );
OAI21X1 OAI21X1_210 ( .A(w_cout_1_), .B(_135_), .C(_136_), .Y(_0__11_) );
INVX1 INVX1_135 ( .A(1'b0), .Y(_140_) );
OR2X2 OR2X2_77 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_141_) );
NAND2X1 NAND2X1_211 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_142_) );
NAND3X1 NAND3X1_77 ( .A(_140_), .B(_142_), .C(_141_), .Y(_143_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_137_) );
AND2X2 AND2X2_77 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_138_) );
OAI21X1 OAI21X1_211 ( .A(_137_), .B(_138_), .C(1'b0), .Y(_139_) );
NAND2X1 NAND2X1_212 ( .A(_139_), .B(_143_), .Y(_9__0_) );
OAI21X1 OAI21X1_212 ( .A(_140_), .B(_137_), .C(_142_), .Y(_11__1_) );
INVX1 INVX1_136 ( .A(_11__3_), .Y(_147_) );
OR2X2 OR2X2_78 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_148_) );
NAND2X1 NAND2X1_213 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_149_) );
NAND3X1 NAND3X1_78 ( .A(_147_), .B(_149_), .C(_148_), .Y(_150_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_144_) );
AND2X2 AND2X2_78 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_145_) );
OAI21X1 OAI21X1_213 ( .A(_144_), .B(_145_), .C(_11__3_), .Y(_146_) );
NAND2X1 NAND2X1_214 ( .A(_146_), .B(_150_), .Y(_9__3_) );
OAI21X1 OAI21X1_214 ( .A(_147_), .B(_144_), .C(_149_), .Y(_7_) );
INVX1 INVX1_137 ( .A(_11__1_), .Y(_154_) );
OR2X2 OR2X2_79 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_155_) );
NAND2X1 NAND2X1_215 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_156_) );
NAND3X1 NAND3X1_79 ( .A(_154_), .B(_156_), .C(_155_), .Y(_157_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_151_) );
AND2X2 AND2X2_79 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_152_) );
OAI21X1 OAI21X1_215 ( .A(_151_), .B(_152_), .C(_11__1_), .Y(_153_) );
NAND2X1 NAND2X1_216 ( .A(_153_), .B(_157_), .Y(_9__1_) );
OAI21X1 OAI21X1_216 ( .A(_154_), .B(_151_), .C(_156_), .Y(_11__2_) );
INVX1 INVX1_138 ( .A(_11__2_), .Y(_161_) );
OR2X2 OR2X2_80 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_162_) );
NAND2X1 NAND2X1_217 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_163_) );
NAND3X1 NAND3X1_80 ( .A(_161_), .B(_163_), .C(_162_), .Y(_164_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_158_) );
AND2X2 AND2X2_80 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_159_) );
OAI21X1 OAI21X1_217 ( .A(_158_), .B(_159_), .C(_11__2_), .Y(_160_) );
NAND2X1 NAND2X1_218 ( .A(_160_), .B(_164_), .Y(_9__2_) );
OAI21X1 OAI21X1_218 ( .A(_161_), .B(_158_), .C(_163_), .Y(_11__3_) );
INVX1 INVX1_139 ( .A(1'b1), .Y(_168_) );
OR2X2 OR2X2_81 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_169_) );
NAND2X1 NAND2X1_219 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_170_) );
NAND3X1 NAND3X1_81 ( .A(_168_), .B(_170_), .C(_169_), .Y(_171_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_165_) );
AND2X2 AND2X2_81 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_166_) );
OAI21X1 OAI21X1_219 ( .A(_165_), .B(_166_), .C(1'b1), .Y(_167_) );
NAND2X1 NAND2X1_220 ( .A(_167_), .B(_171_), .Y(_10__0_) );
OAI21X1 OAI21X1_220 ( .A(_168_), .B(_165_), .C(_170_), .Y(_12__1_) );
INVX1 INVX1_140 ( .A(_12__3_), .Y(_175_) );
OR2X2 OR2X2_82 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_176_) );
NAND2X1 NAND2X1_221 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_177_) );
NAND3X1 NAND3X1_82 ( .A(_175_), .B(_177_), .C(_176_), .Y(_178_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_172_) );
AND2X2 AND2X2_82 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_173_) );
OAI21X1 OAI21X1_221 ( .A(_172_), .B(_173_), .C(_12__3_), .Y(_174_) );
NAND2X1 NAND2X1_222 ( .A(_174_), .B(_178_), .Y(_10__3_) );
OAI21X1 OAI21X1_222 ( .A(_175_), .B(_172_), .C(_177_), .Y(_8_) );
INVX1 INVX1_141 ( .A(_12__1_), .Y(_182_) );
OR2X2 OR2X2_83 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_183_) );
NAND2X1 NAND2X1_223 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_184_) );
NAND3X1 NAND3X1_83 ( .A(_182_), .B(_184_), .C(_183_), .Y(_185_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_179_) );
AND2X2 AND2X2_83 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_180_) );
OAI21X1 OAI21X1_223 ( .A(_179_), .B(_180_), .C(_12__1_), .Y(_181_) );
NAND2X1 NAND2X1_224 ( .A(_181_), .B(_185_), .Y(_10__1_) );
OAI21X1 OAI21X1_224 ( .A(_182_), .B(_179_), .C(_184_), .Y(_12__2_) );
INVX1 INVX1_142 ( .A(_12__2_), .Y(_189_) );
OR2X2 OR2X2_84 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_190_) );
NAND2X1 NAND2X1_225 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_191_) );
NAND3X1 NAND3X1_84 ( .A(_189_), .B(_191_), .C(_190_), .Y(_192_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_186_) );
AND2X2 AND2X2_84 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_187_) );
OAI21X1 OAI21X1_225 ( .A(_186_), .B(_187_), .C(_12__2_), .Y(_188_) );
NAND2X1 NAND2X1_226 ( .A(_188_), .B(_192_), .Y(_10__2_) );
OAI21X1 OAI21X1_226 ( .A(_189_), .B(_186_), .C(_191_), .Y(_12__3_) );
INVX1 INVX1_143 ( .A(_13_), .Y(_193_) );
NAND2X1 NAND2X1_227 ( .A(_14_), .B(w_cout_2_), .Y(_194_) );
OAI21X1 OAI21X1_227 ( .A(w_cout_2_), .B(_193_), .C(_194_), .Y(w_cout_3_) );
BUFX2 BUFX2_49 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_50 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_51 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_52 ( .A(rca_inst_fa31_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_53 ( .A(1'b0), .Y(_0__44_) );
BUFX2 BUFX2_54 ( .A(1'b0), .Y(_0__45_) );
BUFX2 BUFX2_55 ( .A(1'b0), .Y(_0__46_) );
BUFX2 BUFX2_56 ( .A(rca_inst_cout), .Y(w_cout_0_) );
BUFX2 BUFX2_57 ( .A(csa_inst_cin), .Y(w_cout_10_) );
endmodule
