module cla_23bit (i_add1, i_add2, o_result);

input [22:0] i_add1;
input [22:0] i_add2;
output [23:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_93_) );
INVX1 INVX1_1 ( .A(_93_), .Y(w_C_1_) );
NAND2X1 NAND2X1_2 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_94_) );
NAND2X1 NAND2X1_3 ( .A(_93_), .B(_94_), .Y(_95_) );
OAI21X1 OAI21X1_1 ( .A(i_add2[1]), .B(i_add1[1]), .C(_95_), .Y(_96_) );
INVX1 INVX1_2 ( .A(_96_), .Y(w_C_2_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_97_) );
OR2X2 OR2X2_1 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_98_) );
OR2X2 OR2X2_2 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_99_) );
NAND3X1 NAND3X1_1 ( .A(_98_), .B(_99_), .C(_95_), .Y(_100_) );
NAND2X1 NAND2X1_5 ( .A(_97_), .B(_100_), .Y(w_C_3_) );
INVX1 INVX1_3 ( .A(i_add2[3]), .Y(_101_) );
INVX1 INVX1_4 ( .A(i_add1[3]), .Y(_102_) );
NAND2X1 NAND2X1_6 ( .A(_101_), .B(_102_), .Y(_103_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_104_) );
NAND3X1 NAND3X1_2 ( .A(_97_), .B(_104_), .C(_100_), .Y(_105_) );
AND2X2 AND2X2_1 ( .A(_105_), .B(_103_), .Y(w_C_4_) );
NAND2X1 NAND2X1_8 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_106_) );
OR2X2 OR2X2_3 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_107_) );
NAND3X1 NAND3X1_3 ( .A(_103_), .B(_107_), .C(_105_), .Y(_108_) );
NAND2X1 NAND2X1_9 ( .A(_106_), .B(_108_), .Y(w_C_5_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_109_) );
INVX1 INVX1_5 ( .A(_109_), .Y(_110_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_111_) );
NAND3X1 NAND3X1_4 ( .A(_106_), .B(_111_), .C(_108_), .Y(_112_) );
AND2X2 AND2X2_2 ( .A(_112_), .B(_110_), .Y(w_C_6_) );
INVX1 INVX1_6 ( .A(i_add2[6]), .Y(_113_) );
INVX1 INVX1_7 ( .A(i_add1[6]), .Y(_114_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_115_) );
INVX1 INVX1_8 ( .A(_115_), .Y(_116_) );
NAND3X1 NAND3X1_5 ( .A(_110_), .B(_116_), .C(_112_), .Y(_0_) );
OAI21X1 OAI21X1_2 ( .A(_113_), .B(_114_), .C(_0_), .Y(w_C_7_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_1_) );
INVX1 INVX1_9 ( .A(_1_), .Y(_2_) );
NOR2X1 NOR2X1_4 ( .A(_113_), .B(_114_), .Y(_3_) );
INVX1 INVX1_10 ( .A(_3_), .Y(_4_) );
INVX1 INVX1_11 ( .A(i_add2[7]), .Y(_5_) );
INVX1 INVX1_12 ( .A(i_add1[7]), .Y(_6_) );
NOR2X1 NOR2X1_5 ( .A(_5_), .B(_6_), .Y(_7_) );
INVX1 INVX1_13 ( .A(_7_), .Y(_8_) );
NAND3X1 NAND3X1_6 ( .A(_4_), .B(_8_), .C(_0_), .Y(_9_) );
AND2X2 AND2X2_3 ( .A(_9_), .B(_2_), .Y(w_C_8_) );
INVX1 INVX1_14 ( .A(i_add2[8]), .Y(_10_) );
INVX1 INVX1_15 ( .A(i_add1[8]), .Y(_11_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_12_) );
INVX1 INVX1_16 ( .A(_12_), .Y(_13_) );
NAND3X1 NAND3X1_7 ( .A(_2_), .B(_13_), .C(_9_), .Y(_14_) );
OAI21X1 OAI21X1_3 ( .A(_10_), .B(_11_), .C(_14_), .Y(w_C_9_) );
NOR2X1 NOR2X1_7 ( .A(_10_), .B(_11_), .Y(_15_) );
INVX1 INVX1_17 ( .A(_15_), .Y(_16_) );
AND2X2 AND2X2_4 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_17_) );
INVX1 INVX1_18 ( .A(_17_), .Y(_18_) );
NAND3X1 NAND3X1_8 ( .A(_16_), .B(_18_), .C(_14_), .Y(_19_) );
OAI21X1 OAI21X1_4 ( .A(i_add2[9]), .B(i_add1[9]), .C(_19_), .Y(_20_) );
INVX1 INVX1_19 ( .A(_20_), .Y(w_C_10_) );
INVX1 INVX1_20 ( .A(i_add2[10]), .Y(_21_) );
INVX1 INVX1_21 ( .A(i_add1[10]), .Y(_22_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_23_) );
INVX1 INVX1_22 ( .A(_23_), .Y(_24_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_25_) );
INVX1 INVX1_23 ( .A(_25_), .Y(_26_) );
NAND3X1 NAND3X1_9 ( .A(_24_), .B(_26_), .C(_19_), .Y(_27_) );
OAI21X1 OAI21X1_5 ( .A(_21_), .B(_22_), .C(_27_), .Y(w_C_11_) );
NOR2X1 NOR2X1_10 ( .A(_21_), .B(_22_), .Y(_28_) );
INVX1 INVX1_24 ( .A(_28_), .Y(_29_) );
AND2X2 AND2X2_5 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_30_) );
INVX1 INVX1_25 ( .A(_30_), .Y(_31_) );
NAND3X1 NAND3X1_10 ( .A(_29_), .B(_31_), .C(_27_), .Y(_32_) );
OAI21X1 OAI21X1_6 ( .A(i_add2[11]), .B(i_add1[11]), .C(_32_), .Y(_33_) );
INVX1 INVX1_26 ( .A(_33_), .Y(w_C_12_) );
INVX1 INVX1_27 ( .A(i_add2[12]), .Y(_34_) );
INVX1 INVX1_28 ( .A(i_add1[12]), .Y(_35_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_36_) );
INVX1 INVX1_29 ( .A(_36_), .Y(_37_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_38_) );
INVX1 INVX1_30 ( .A(_38_), .Y(_39_) );
NAND3X1 NAND3X1_11 ( .A(_37_), .B(_39_), .C(_32_), .Y(_40_) );
OAI21X1 OAI21X1_7 ( .A(_34_), .B(_35_), .C(_40_), .Y(w_C_13_) );
NOR2X1 NOR2X1_13 ( .A(_34_), .B(_35_), .Y(_41_) );
INVX1 INVX1_31 ( .A(_41_), .Y(_42_) );
AND2X2 AND2X2_6 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_43_) );
INVX1 INVX1_32 ( .A(_43_), .Y(_44_) );
NAND3X1 NAND3X1_12 ( .A(_42_), .B(_44_), .C(_40_), .Y(_45_) );
OAI21X1 OAI21X1_8 ( .A(i_add2[13]), .B(i_add1[13]), .C(_45_), .Y(_46_) );
INVX1 INVX1_33 ( .A(_46_), .Y(w_C_14_) );
INVX1 INVX1_34 ( .A(i_add2[14]), .Y(_47_) );
INVX1 INVX1_35 ( .A(i_add1[14]), .Y(_48_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_49_) );
INVX1 INVX1_36 ( .A(_49_), .Y(_50_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_51_) );
INVX1 INVX1_37 ( .A(_51_), .Y(_52_) );
NAND3X1 NAND3X1_13 ( .A(_50_), .B(_52_), .C(_45_), .Y(_53_) );
OAI21X1 OAI21X1_9 ( .A(_47_), .B(_48_), .C(_53_), .Y(w_C_15_) );
NOR2X1 NOR2X1_16 ( .A(_47_), .B(_48_), .Y(_54_) );
INVX1 INVX1_38 ( .A(_54_), .Y(_55_) );
AND2X2 AND2X2_7 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_56_) );
INVX1 INVX1_39 ( .A(_56_), .Y(_57_) );
NAND3X1 NAND3X1_14 ( .A(_55_), .B(_57_), .C(_53_), .Y(_58_) );
OAI21X1 OAI21X1_10 ( .A(i_add2[15]), .B(i_add1[15]), .C(_58_), .Y(_59_) );
INVX1 INVX1_40 ( .A(_59_), .Y(w_C_16_) );
INVX1 INVX1_41 ( .A(i_add2[16]), .Y(_60_) );
INVX1 INVX1_42 ( .A(i_add1[16]), .Y(_61_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_62_) );
INVX1 INVX1_43 ( .A(_62_), .Y(_63_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_64_) );
INVX1 INVX1_44 ( .A(_64_), .Y(_65_) );
NAND3X1 NAND3X1_15 ( .A(_63_), .B(_65_), .C(_58_), .Y(_66_) );
OAI21X1 OAI21X1_11 ( .A(_60_), .B(_61_), .C(_66_), .Y(w_C_17_) );
NOR2X1 NOR2X1_19 ( .A(_60_), .B(_61_), .Y(_67_) );
INVX1 INVX1_45 ( .A(_67_), .Y(_68_) );
AND2X2 AND2X2_8 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_69_) );
INVX1 INVX1_46 ( .A(_69_), .Y(_70_) );
NAND3X1 NAND3X1_16 ( .A(_68_), .B(_70_), .C(_66_), .Y(_71_) );
OAI21X1 OAI21X1_12 ( .A(i_add2[17]), .B(i_add1[17]), .C(_71_), .Y(_72_) );
INVX1 INVX1_47 ( .A(_72_), .Y(w_C_18_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_73_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_74_) );
OAI21X1 OAI21X1_13 ( .A(_74_), .B(_72_), .C(_73_), .Y(w_C_19_) );
OR2X2 OR2X2_4 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_75_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_76_) );
INVX1 INVX1_48 ( .A(_76_), .Y(_77_) );
INVX1 INVX1_49 ( .A(_74_), .Y(_78_) );
NAND3X1 NAND3X1_17 ( .A(_77_), .B(_78_), .C(_71_), .Y(_79_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_80_) );
NAND3X1 NAND3X1_18 ( .A(_73_), .B(_80_), .C(_79_), .Y(_81_) );
AND2X2 AND2X2_9 ( .A(_81_), .B(_75_), .Y(w_C_20_) );
INVX1 INVX1_50 ( .A(i_add2[20]), .Y(_82_) );
INVX1 INVX1_51 ( .A(i_add1[20]), .Y(_83_) );
NAND2X1 NAND2X1_13 ( .A(_82_), .B(_83_), .Y(_84_) );
NAND3X1 NAND3X1_19 ( .A(_75_), .B(_84_), .C(_81_), .Y(_85_) );
OAI21X1 OAI21X1_14 ( .A(_82_), .B(_83_), .C(_85_), .Y(w_C_21_) );
OR2X2 OR2X2_5 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_86_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_87_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_88_) );
NAND3X1 NAND3X1_20 ( .A(_87_), .B(_88_), .C(_85_), .Y(_89_) );
AND2X2 AND2X2_10 ( .A(_89_), .B(_86_), .Y(w_C_22_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_90_) );
OR2X2 OR2X2_6 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_91_) );
NAND3X1 NAND3X1_21 ( .A(_86_), .B(_91_), .C(_89_), .Y(_92_) );
NAND2X1 NAND2X1_17 ( .A(_90_), .B(_92_), .Y(w_C_23_) );
BUFX2 BUFX2_1 ( .A(_117__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_117__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_117__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_117__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_117__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_117__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_117__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_117__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_117__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_117__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_117__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_117__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_117__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_117__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_117__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_117__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_117__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_117__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_117__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_117__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_117__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_117__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_117__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(w_C_23_), .Y(o_result[23]) );
INVX1 INVX1_52 ( .A(w_C_4_), .Y(_121_) );
OR2X2 OR2X2_7 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_122_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_123_) );
NAND3X1 NAND3X1_22 ( .A(_121_), .B(_123_), .C(_122_), .Y(_124_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_118_) );
AND2X2 AND2X2_11 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_119_) );
OAI21X1 OAI21X1_15 ( .A(_118_), .B(_119_), .C(w_C_4_), .Y(_120_) );
NAND2X1 NAND2X1_19 ( .A(_120_), .B(_124_), .Y(_117__4_) );
INVX1 INVX1_53 ( .A(w_C_5_), .Y(_128_) );
OR2X2 OR2X2_8 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_129_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_130_) );
NAND3X1 NAND3X1_23 ( .A(_128_), .B(_130_), .C(_129_), .Y(_131_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_125_) );
AND2X2 AND2X2_12 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_126_) );
OAI21X1 OAI21X1_16 ( .A(_125_), .B(_126_), .C(w_C_5_), .Y(_127_) );
NAND2X1 NAND2X1_21 ( .A(_127_), .B(_131_), .Y(_117__5_) );
INVX1 INVX1_54 ( .A(w_C_6_), .Y(_135_) );
OR2X2 OR2X2_9 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_136_) );
NAND2X1 NAND2X1_22 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_137_) );
NAND3X1 NAND3X1_24 ( .A(_135_), .B(_137_), .C(_136_), .Y(_138_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_132_) );
AND2X2 AND2X2_13 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_133_) );
OAI21X1 OAI21X1_17 ( .A(_132_), .B(_133_), .C(w_C_6_), .Y(_134_) );
NAND2X1 NAND2X1_23 ( .A(_134_), .B(_138_), .Y(_117__6_) );
INVX1 INVX1_55 ( .A(w_C_7_), .Y(_142_) );
OR2X2 OR2X2_10 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_143_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_144_) );
NAND3X1 NAND3X1_25 ( .A(_142_), .B(_144_), .C(_143_), .Y(_145_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_139_) );
AND2X2 AND2X2_14 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_140_) );
OAI21X1 OAI21X1_18 ( .A(_139_), .B(_140_), .C(w_C_7_), .Y(_141_) );
NAND2X1 NAND2X1_25 ( .A(_141_), .B(_145_), .Y(_117__7_) );
INVX1 INVX1_56 ( .A(w_C_8_), .Y(_149_) );
OR2X2 OR2X2_11 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_150_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_151_) );
NAND3X1 NAND3X1_26 ( .A(_149_), .B(_151_), .C(_150_), .Y(_152_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_146_) );
AND2X2 AND2X2_15 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_147_) );
OAI21X1 OAI21X1_19 ( .A(_146_), .B(_147_), .C(w_C_8_), .Y(_148_) );
NAND2X1 NAND2X1_27 ( .A(_148_), .B(_152_), .Y(_117__8_) );
INVX1 INVX1_57 ( .A(w_C_9_), .Y(_156_) );
OR2X2 OR2X2_12 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_157_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_158_) );
NAND3X1 NAND3X1_27 ( .A(_156_), .B(_158_), .C(_157_), .Y(_159_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_153_) );
AND2X2 AND2X2_16 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_154_) );
OAI21X1 OAI21X1_20 ( .A(_153_), .B(_154_), .C(w_C_9_), .Y(_155_) );
NAND2X1 NAND2X1_29 ( .A(_155_), .B(_159_), .Y(_117__9_) );
INVX1 INVX1_58 ( .A(w_C_10_), .Y(_163_) );
OR2X2 OR2X2_13 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_164_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_165_) );
NAND3X1 NAND3X1_28 ( .A(_163_), .B(_165_), .C(_164_), .Y(_166_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_160_) );
AND2X2 AND2X2_17 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_161_) );
OAI21X1 OAI21X1_21 ( .A(_160_), .B(_161_), .C(w_C_10_), .Y(_162_) );
NAND2X1 NAND2X1_31 ( .A(_162_), .B(_166_), .Y(_117__10_) );
INVX1 INVX1_59 ( .A(w_C_11_), .Y(_170_) );
OR2X2 OR2X2_14 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_171_) );
NAND2X1 NAND2X1_32 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_172_) );
NAND3X1 NAND3X1_29 ( .A(_170_), .B(_172_), .C(_171_), .Y(_173_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_167_) );
AND2X2 AND2X2_18 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_168_) );
OAI21X1 OAI21X1_22 ( .A(_167_), .B(_168_), .C(w_C_11_), .Y(_169_) );
NAND2X1 NAND2X1_33 ( .A(_169_), .B(_173_), .Y(_117__11_) );
INVX1 INVX1_60 ( .A(w_C_12_), .Y(_177_) );
OR2X2 OR2X2_15 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_178_) );
NAND2X1 NAND2X1_34 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_179_) );
NAND3X1 NAND3X1_30 ( .A(_177_), .B(_179_), .C(_178_), .Y(_180_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_174_) );
AND2X2 AND2X2_19 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_175_) );
OAI21X1 OAI21X1_23 ( .A(_174_), .B(_175_), .C(w_C_12_), .Y(_176_) );
NAND2X1 NAND2X1_35 ( .A(_176_), .B(_180_), .Y(_117__12_) );
INVX1 INVX1_61 ( .A(w_C_13_), .Y(_184_) );
OR2X2 OR2X2_16 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_185_) );
NAND2X1 NAND2X1_36 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_186_) );
NAND3X1 NAND3X1_31 ( .A(_184_), .B(_186_), .C(_185_), .Y(_187_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_181_) );
AND2X2 AND2X2_20 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_182_) );
OAI21X1 OAI21X1_24 ( .A(_181_), .B(_182_), .C(w_C_13_), .Y(_183_) );
NAND2X1 NAND2X1_37 ( .A(_183_), .B(_187_), .Y(_117__13_) );
INVX1 INVX1_62 ( .A(w_C_14_), .Y(_191_) );
OR2X2 OR2X2_17 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_192_) );
NAND2X1 NAND2X1_38 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_193_) );
NAND3X1 NAND3X1_32 ( .A(_191_), .B(_193_), .C(_192_), .Y(_194_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_188_) );
AND2X2 AND2X2_21 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_189_) );
OAI21X1 OAI21X1_25 ( .A(_188_), .B(_189_), .C(w_C_14_), .Y(_190_) );
NAND2X1 NAND2X1_39 ( .A(_190_), .B(_194_), .Y(_117__14_) );
INVX1 INVX1_63 ( .A(w_C_15_), .Y(_198_) );
OR2X2 OR2X2_18 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_199_) );
NAND2X1 NAND2X1_40 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_200_) );
NAND3X1 NAND3X1_33 ( .A(_198_), .B(_200_), .C(_199_), .Y(_201_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_195_) );
AND2X2 AND2X2_22 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_196_) );
OAI21X1 OAI21X1_26 ( .A(_195_), .B(_196_), .C(w_C_15_), .Y(_197_) );
NAND2X1 NAND2X1_41 ( .A(_197_), .B(_201_), .Y(_117__15_) );
INVX1 INVX1_64 ( .A(w_C_16_), .Y(_205_) );
OR2X2 OR2X2_19 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_206_) );
NAND2X1 NAND2X1_42 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_207_) );
NAND3X1 NAND3X1_34 ( .A(_205_), .B(_207_), .C(_206_), .Y(_208_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_202_) );
AND2X2 AND2X2_23 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_203_) );
OAI21X1 OAI21X1_27 ( .A(_202_), .B(_203_), .C(w_C_16_), .Y(_204_) );
NAND2X1 NAND2X1_43 ( .A(_204_), .B(_208_), .Y(_117__16_) );
INVX1 INVX1_65 ( .A(w_C_17_), .Y(_212_) );
OR2X2 OR2X2_20 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_213_) );
NAND2X1 NAND2X1_44 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_214_) );
NAND3X1 NAND3X1_35 ( .A(_212_), .B(_214_), .C(_213_), .Y(_215_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_209_) );
AND2X2 AND2X2_24 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_210_) );
OAI21X1 OAI21X1_28 ( .A(_209_), .B(_210_), .C(w_C_17_), .Y(_211_) );
NAND2X1 NAND2X1_45 ( .A(_211_), .B(_215_), .Y(_117__17_) );
INVX1 INVX1_66 ( .A(w_C_18_), .Y(_219_) );
OR2X2 OR2X2_21 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_220_) );
NAND2X1 NAND2X1_46 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_221_) );
NAND3X1 NAND3X1_36 ( .A(_219_), .B(_221_), .C(_220_), .Y(_222_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_216_) );
AND2X2 AND2X2_25 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_217_) );
OAI21X1 OAI21X1_29 ( .A(_216_), .B(_217_), .C(w_C_18_), .Y(_218_) );
NAND2X1 NAND2X1_47 ( .A(_218_), .B(_222_), .Y(_117__18_) );
INVX1 INVX1_67 ( .A(w_C_19_), .Y(_226_) );
OR2X2 OR2X2_22 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_227_) );
NAND2X1 NAND2X1_48 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_228_) );
NAND3X1 NAND3X1_37 ( .A(_226_), .B(_228_), .C(_227_), .Y(_229_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_223_) );
AND2X2 AND2X2_26 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_224_) );
OAI21X1 OAI21X1_30 ( .A(_223_), .B(_224_), .C(w_C_19_), .Y(_225_) );
NAND2X1 NAND2X1_49 ( .A(_225_), .B(_229_), .Y(_117__19_) );
INVX1 INVX1_68 ( .A(w_C_20_), .Y(_233_) );
OR2X2 OR2X2_23 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_234_) );
NAND2X1 NAND2X1_50 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_235_) );
NAND3X1 NAND3X1_38 ( .A(_233_), .B(_235_), .C(_234_), .Y(_236_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_230_) );
AND2X2 AND2X2_27 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_231_) );
OAI21X1 OAI21X1_31 ( .A(_230_), .B(_231_), .C(w_C_20_), .Y(_232_) );
NAND2X1 NAND2X1_51 ( .A(_232_), .B(_236_), .Y(_117__20_) );
INVX1 INVX1_69 ( .A(w_C_21_), .Y(_240_) );
OR2X2 OR2X2_24 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_241_) );
NAND2X1 NAND2X1_52 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_242_) );
NAND3X1 NAND3X1_39 ( .A(_240_), .B(_242_), .C(_241_), .Y(_243_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_237_) );
AND2X2 AND2X2_28 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_238_) );
OAI21X1 OAI21X1_32 ( .A(_237_), .B(_238_), .C(w_C_21_), .Y(_239_) );
NAND2X1 NAND2X1_53 ( .A(_239_), .B(_243_), .Y(_117__21_) );
INVX1 INVX1_70 ( .A(w_C_22_), .Y(_247_) );
OR2X2 OR2X2_25 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_248_) );
NAND2X1 NAND2X1_54 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_249_) );
NAND3X1 NAND3X1_40 ( .A(_247_), .B(_249_), .C(_248_), .Y(_250_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_244_) );
AND2X2 AND2X2_29 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_245_) );
OAI21X1 OAI21X1_33 ( .A(_244_), .B(_245_), .C(w_C_22_), .Y(_246_) );
NAND2X1 NAND2X1_55 ( .A(_246_), .B(_250_), .Y(_117__22_) );
INVX1 INVX1_71 ( .A(gnd), .Y(_254_) );
OR2X2 OR2X2_26 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_255_) );
NAND2X1 NAND2X1_56 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_256_) );
NAND3X1 NAND3X1_41 ( .A(_254_), .B(_256_), .C(_255_), .Y(_257_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_251_) );
AND2X2 AND2X2_30 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_252_) );
OAI21X1 OAI21X1_34 ( .A(_251_), .B(_252_), .C(gnd), .Y(_253_) );
NAND2X1 NAND2X1_57 ( .A(_253_), .B(_257_), .Y(_117__0_) );
INVX1 INVX1_72 ( .A(w_C_1_), .Y(_261_) );
OR2X2 OR2X2_27 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_262_) );
NAND2X1 NAND2X1_58 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_263_) );
NAND3X1 NAND3X1_42 ( .A(_261_), .B(_263_), .C(_262_), .Y(_264_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_258_) );
AND2X2 AND2X2_31 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_259_) );
OAI21X1 OAI21X1_35 ( .A(_258_), .B(_259_), .C(w_C_1_), .Y(_260_) );
NAND2X1 NAND2X1_59 ( .A(_260_), .B(_264_), .Y(_117__1_) );
INVX1 INVX1_73 ( .A(w_C_2_), .Y(_268_) );
OR2X2 OR2X2_28 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_269_) );
NAND2X1 NAND2X1_60 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_270_) );
NAND3X1 NAND3X1_43 ( .A(_268_), .B(_270_), .C(_269_), .Y(_271_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_265_) );
AND2X2 AND2X2_32 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_266_) );
OAI21X1 OAI21X1_36 ( .A(_265_), .B(_266_), .C(w_C_2_), .Y(_267_) );
NAND2X1 NAND2X1_61 ( .A(_267_), .B(_271_), .Y(_117__2_) );
INVX1 INVX1_74 ( .A(w_C_3_), .Y(_275_) );
OR2X2 OR2X2_29 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_276_) );
NAND2X1 NAND2X1_62 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_277_) );
NAND3X1 NAND3X1_44 ( .A(_275_), .B(_277_), .C(_276_), .Y(_278_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_272_) );
AND2X2 AND2X2_33 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_273_) );
OAI21X1 OAI21X1_37 ( .A(_272_), .B(_273_), .C(w_C_3_), .Y(_274_) );
NAND2X1 NAND2X1_63 ( .A(_274_), .B(_278_), .Y(_117__3_) );
BUFX2 BUFX2_25 ( .A(w_C_23_), .Y(_117__23_) );
BUFX2 BUFX2_26 ( .A(gnd), .Y(w_C_0_) );
endmodule
