module csa_61bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term1[45], i_add_term1[46], i_add_term1[47], i_add_term1[48], i_add_term1[49], i_add_term1[50], i_add_term1[51], i_add_term1[52], i_add_term1[53], i_add_term1[54], i_add_term1[55], i_add_term1[56], i_add_term1[57], i_add_term1[58], i_add_term1[59], i_add_term1[60], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], i_add_term2[45], i_add_term2[46], i_add_term2[47], i_add_term2[48], i_add_term2[49], i_add_term2[50], i_add_term2[51], i_add_term2[52], i_add_term2[53], i_add_term2[54], i_add_term2[55], i_add_term2[56], i_add_term2[57], i_add_term2[58], i_add_term2[59], i_add_term2[60], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], sum[45], sum[46], sum[47], sum[48], sum[49], sum[50], sum[51], sum[52], sum[53], sum[54], sum[55], sum[56], sum[57], sum[58], sum[59], sum[60], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term1[45];
input i_add_term1[46];
input i_add_term1[47];
input i_add_term1[48];
input i_add_term1[49];
input i_add_term1[50];
input i_add_term1[51];
input i_add_term1[52];
input i_add_term1[53];
input i_add_term1[54];
input i_add_term1[55];
input i_add_term1[56];
input i_add_term1[57];
input i_add_term1[58];
input i_add_term1[59];
input i_add_term1[60];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
input i_add_term2[45];
input i_add_term2[46];
input i_add_term2[47];
input i_add_term2[48];
input i_add_term2[49];
input i_add_term2[50];
input i_add_term2[51];
input i_add_term2[52];
input i_add_term2[53];
input i_add_term2[54];
input i_add_term2[55];
input i_add_term2[56];
input i_add_term2[57];
input i_add_term2[58];
input i_add_term2[59];
input i_add_term2[60];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output sum[45];
output sum[46];
output sum[47];
output sum[48];
output sum[49];
output sum[50];
output sum[51];
output sum[52];
output sum[53];
output sum[54];
output sum[55];
output sum[56];
output sum[57];
output sum[58];
output sum[59];
output sum[60];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_15_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_w_SUM), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .A(_0__54_), .Y(sum[54]) );
BUFX2 BUFX2_57 ( .A(_0__55_), .Y(sum[55]) );
BUFX2 BUFX2_58 ( .A(_0__56_), .Y(sum[56]) );
BUFX2 BUFX2_59 ( .A(_0__57_), .Y(sum[57]) );
BUFX2 BUFX2_60 ( .A(_0__58_), .Y(sum[58]) );
BUFX2 BUFX2_61 ( .A(_0__59_), .Y(sum[59]) );
BUFX2 BUFX2_62 ( .A(_0__60_), .Y(sum[60]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_91_) );
NAND2X1 NAND2X1_1 ( .A(_2_), .B(1'b0), .Y(_92_) );
OAI21X1 OAI21X1_1 ( .A(1'b0), .B(_91_), .C(_92_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3__0_), .Y(_93_) );
NAND2X1 NAND2X1_2 ( .A(_4__0_), .B(1'b0), .Y(_94_) );
OAI21X1 OAI21X1_2 ( .A(1'b0), .B(_93_), .C(_94_), .Y(_0__1_) );
INVX1 INVX1_3 ( .A(_3__1_), .Y(_95_) );
NAND2X1 NAND2X1_3 ( .A(1'b0), .B(_4__1_), .Y(_96_) );
OAI21X1 OAI21X1_3 ( .A(1'b0), .B(_95_), .C(_96_), .Y(_0__2_) );
INVX1 INVX1_4 ( .A(_3__2_), .Y(_97_) );
NAND2X1 NAND2X1_4 ( .A(1'b0), .B(_4__2_), .Y(_98_) );
OAI21X1 OAI21X1_4 ( .A(1'b0), .B(_97_), .C(_98_), .Y(_0__3_) );
INVX1 INVX1_5 ( .A(_3__3_), .Y(_99_) );
NAND2X1 NAND2X1_5 ( .A(1'b0), .B(_4__3_), .Y(_100_) );
OAI21X1 OAI21X1_5 ( .A(1'b0), .B(_99_), .C(_100_), .Y(_0__4_) );
INVX1 INVX1_6 ( .A(_7_), .Y(_101_) );
NAND2X1 NAND2X1_6 ( .A(_8_), .B(w_cout_1_), .Y(_102_) );
OAI21X1 OAI21X1_6 ( .A(w_cout_1_), .B(_101_), .C(_102_), .Y(w_cout_2_) );
INVX1 INVX1_7 ( .A(_9__0_), .Y(_103_) );
NAND2X1 NAND2X1_7 ( .A(_10__0_), .B(w_cout_1_), .Y(_104_) );
OAI21X1 OAI21X1_7 ( .A(w_cout_1_), .B(_103_), .C(_104_), .Y(_0__5_) );
INVX1 INVX1_8 ( .A(_9__1_), .Y(_105_) );
NAND2X1 NAND2X1_8 ( .A(w_cout_1_), .B(_10__1_), .Y(_106_) );
OAI21X1 OAI21X1_8 ( .A(w_cout_1_), .B(_105_), .C(_106_), .Y(_0__6_) );
INVX1 INVX1_9 ( .A(_9__2_), .Y(_107_) );
NAND2X1 NAND2X1_9 ( .A(w_cout_1_), .B(_10__2_), .Y(_108_) );
OAI21X1 OAI21X1_9 ( .A(w_cout_1_), .B(_107_), .C(_108_), .Y(_0__7_) );
INVX1 INVX1_10 ( .A(_9__3_), .Y(_109_) );
NAND2X1 NAND2X1_10 ( .A(w_cout_1_), .B(_10__3_), .Y(_110_) );
OAI21X1 OAI21X1_10 ( .A(w_cout_1_), .B(_109_), .C(_110_), .Y(_0__8_) );
INVX1 INVX1_11 ( .A(_13_), .Y(_111_) );
NAND2X1 NAND2X1_11 ( .A(_14_), .B(w_cout_2_), .Y(_112_) );
OAI21X1 OAI21X1_11 ( .A(w_cout_2_), .B(_111_), .C(_112_), .Y(w_cout_3_) );
INVX1 INVX1_12 ( .A(_15__0_), .Y(_113_) );
NAND2X1 NAND2X1_12 ( .A(_16__0_), .B(w_cout_2_), .Y(_114_) );
OAI21X1 OAI21X1_12 ( .A(w_cout_2_), .B(_113_), .C(_114_), .Y(_0__9_) );
INVX1 INVX1_13 ( .A(_15__1_), .Y(_115_) );
NAND2X1 NAND2X1_13 ( .A(w_cout_2_), .B(_16__1_), .Y(_116_) );
OAI21X1 OAI21X1_13 ( .A(w_cout_2_), .B(_115_), .C(_116_), .Y(_0__10_) );
INVX1 INVX1_14 ( .A(_15__2_), .Y(_117_) );
NAND2X1 NAND2X1_14 ( .A(w_cout_2_), .B(_16__2_), .Y(_118_) );
OAI21X1 OAI21X1_14 ( .A(w_cout_2_), .B(_117_), .C(_118_), .Y(_0__11_) );
INVX1 INVX1_15 ( .A(_15__3_), .Y(_119_) );
NAND2X1 NAND2X1_15 ( .A(w_cout_2_), .B(_16__3_), .Y(_120_) );
OAI21X1 OAI21X1_15 ( .A(w_cout_2_), .B(_119_), .C(_120_), .Y(_0__12_) );
INVX1 INVX1_16 ( .A(_19_), .Y(_121_) );
NAND2X1 NAND2X1_16 ( .A(_20_), .B(w_cout_3_), .Y(_122_) );
OAI21X1 OAI21X1_16 ( .A(w_cout_3_), .B(_121_), .C(_122_), .Y(w_cout_4_) );
INVX1 INVX1_17 ( .A(_21__0_), .Y(_123_) );
NAND2X1 NAND2X1_17 ( .A(_22__0_), .B(w_cout_3_), .Y(_124_) );
OAI21X1 OAI21X1_17 ( .A(w_cout_3_), .B(_123_), .C(_124_), .Y(_0__13_) );
INVX1 INVX1_18 ( .A(_21__1_), .Y(_125_) );
NAND2X1 NAND2X1_18 ( .A(w_cout_3_), .B(_22__1_), .Y(_126_) );
OAI21X1 OAI21X1_18 ( .A(w_cout_3_), .B(_125_), .C(_126_), .Y(_0__14_) );
INVX1 INVX1_19 ( .A(_21__2_), .Y(_127_) );
NAND2X1 NAND2X1_19 ( .A(w_cout_3_), .B(_22__2_), .Y(_128_) );
OAI21X1 OAI21X1_19 ( .A(w_cout_3_), .B(_127_), .C(_128_), .Y(_0__15_) );
INVX1 INVX1_20 ( .A(_21__3_), .Y(_129_) );
NAND2X1 NAND2X1_20 ( .A(w_cout_3_), .B(_22__3_), .Y(_130_) );
OAI21X1 OAI21X1_20 ( .A(w_cout_3_), .B(_129_), .C(_130_), .Y(_0__16_) );
INVX1 INVX1_21 ( .A(_25_), .Y(_131_) );
NAND2X1 NAND2X1_21 ( .A(_26_), .B(w_cout_4_), .Y(_132_) );
OAI21X1 OAI21X1_21 ( .A(w_cout_4_), .B(_131_), .C(_132_), .Y(w_cout_5_) );
INVX1 INVX1_22 ( .A(_27__0_), .Y(_133_) );
NAND2X1 NAND2X1_22 ( .A(_28__0_), .B(w_cout_4_), .Y(_134_) );
OAI21X1 OAI21X1_22 ( .A(w_cout_4_), .B(_133_), .C(_134_), .Y(_0__17_) );
INVX1 INVX1_23 ( .A(_27__1_), .Y(_135_) );
NAND2X1 NAND2X1_23 ( .A(w_cout_4_), .B(_28__1_), .Y(_136_) );
OAI21X1 OAI21X1_23 ( .A(w_cout_4_), .B(_135_), .C(_136_), .Y(_0__18_) );
INVX1 INVX1_24 ( .A(_27__2_), .Y(_137_) );
NAND2X1 NAND2X1_24 ( .A(w_cout_4_), .B(_28__2_), .Y(_138_) );
OAI21X1 OAI21X1_24 ( .A(w_cout_4_), .B(_137_), .C(_138_), .Y(_0__19_) );
INVX1 INVX1_25 ( .A(_27__3_), .Y(_139_) );
NAND2X1 NAND2X1_25 ( .A(w_cout_4_), .B(_28__3_), .Y(_140_) );
OAI21X1 OAI21X1_25 ( .A(w_cout_4_), .B(_139_), .C(_140_), .Y(_0__20_) );
INVX1 INVX1_26 ( .A(_31_), .Y(_141_) );
NAND2X1 NAND2X1_26 ( .A(_32_), .B(w_cout_5_), .Y(_142_) );
OAI21X1 OAI21X1_26 ( .A(w_cout_5_), .B(_141_), .C(_142_), .Y(w_cout_6_) );
INVX1 INVX1_27 ( .A(_33__0_), .Y(_143_) );
NAND2X1 NAND2X1_27 ( .A(_34__0_), .B(w_cout_5_), .Y(_144_) );
OAI21X1 OAI21X1_27 ( .A(w_cout_5_), .B(_143_), .C(_144_), .Y(_0__21_) );
INVX1 INVX1_28 ( .A(_33__1_), .Y(_145_) );
NAND2X1 NAND2X1_28 ( .A(w_cout_5_), .B(_34__1_), .Y(_146_) );
OAI21X1 OAI21X1_28 ( .A(w_cout_5_), .B(_145_), .C(_146_), .Y(_0__22_) );
INVX1 INVX1_29 ( .A(_33__2_), .Y(_147_) );
NAND2X1 NAND2X1_29 ( .A(w_cout_5_), .B(_34__2_), .Y(_148_) );
OAI21X1 OAI21X1_29 ( .A(w_cout_5_), .B(_147_), .C(_148_), .Y(_0__23_) );
INVX1 INVX1_30 ( .A(_33__3_), .Y(_149_) );
NAND2X1 NAND2X1_30 ( .A(w_cout_5_), .B(_34__3_), .Y(_150_) );
OAI21X1 OAI21X1_30 ( .A(w_cout_5_), .B(_149_), .C(_150_), .Y(_0__24_) );
INVX1 INVX1_31 ( .A(_37_), .Y(_151_) );
NAND2X1 NAND2X1_31 ( .A(_38_), .B(w_cout_6_), .Y(_152_) );
OAI21X1 OAI21X1_31 ( .A(w_cout_6_), .B(_151_), .C(_152_), .Y(w_cout_7_) );
INVX1 INVX1_32 ( .A(_39__0_), .Y(_153_) );
NAND2X1 NAND2X1_32 ( .A(_40__0_), .B(w_cout_6_), .Y(_154_) );
OAI21X1 OAI21X1_32 ( .A(w_cout_6_), .B(_153_), .C(_154_), .Y(_0__25_) );
INVX1 INVX1_33 ( .A(_39__1_), .Y(_155_) );
NAND2X1 NAND2X1_33 ( .A(w_cout_6_), .B(_40__1_), .Y(_156_) );
OAI21X1 OAI21X1_33 ( .A(w_cout_6_), .B(_155_), .C(_156_), .Y(_0__26_) );
INVX1 INVX1_34 ( .A(_39__2_), .Y(_157_) );
NAND2X1 NAND2X1_34 ( .A(w_cout_6_), .B(_40__2_), .Y(_158_) );
OAI21X1 OAI21X1_34 ( .A(w_cout_6_), .B(_157_), .C(_158_), .Y(_0__27_) );
INVX1 INVX1_35 ( .A(_39__3_), .Y(_159_) );
NAND2X1 NAND2X1_35 ( .A(w_cout_6_), .B(_40__3_), .Y(_160_) );
OAI21X1 OAI21X1_35 ( .A(w_cout_6_), .B(_159_), .C(_160_), .Y(_0__28_) );
INVX1 INVX1_36 ( .A(_43_), .Y(_161_) );
NAND2X1 NAND2X1_36 ( .A(_44_), .B(w_cout_7_), .Y(_162_) );
OAI21X1 OAI21X1_36 ( .A(w_cout_7_), .B(_161_), .C(_162_), .Y(w_cout_8_) );
INVX1 INVX1_37 ( .A(_45__0_), .Y(_163_) );
NAND2X1 NAND2X1_37 ( .A(_46__0_), .B(w_cout_7_), .Y(_164_) );
OAI21X1 OAI21X1_37 ( .A(w_cout_7_), .B(_163_), .C(_164_), .Y(_0__29_) );
INVX1 INVX1_38 ( .A(_45__1_), .Y(_165_) );
NAND2X1 NAND2X1_38 ( .A(w_cout_7_), .B(_46__1_), .Y(_166_) );
OAI21X1 OAI21X1_38 ( .A(w_cout_7_), .B(_165_), .C(_166_), .Y(_0__30_) );
INVX1 INVX1_39 ( .A(_45__2_), .Y(_167_) );
NAND2X1 NAND2X1_39 ( .A(w_cout_7_), .B(_46__2_), .Y(_168_) );
OAI21X1 OAI21X1_39 ( .A(w_cout_7_), .B(_167_), .C(_168_), .Y(_0__31_) );
INVX1 INVX1_40 ( .A(_45__3_), .Y(_169_) );
NAND2X1 NAND2X1_40 ( .A(w_cout_7_), .B(_46__3_), .Y(_170_) );
OAI21X1 OAI21X1_40 ( .A(w_cout_7_), .B(_169_), .C(_170_), .Y(_0__32_) );
INVX1 INVX1_41 ( .A(_49_), .Y(_171_) );
NAND2X1 NAND2X1_41 ( .A(_50_), .B(w_cout_8_), .Y(_172_) );
OAI21X1 OAI21X1_41 ( .A(w_cout_8_), .B(_171_), .C(_172_), .Y(w_cout_9_) );
INVX1 INVX1_42 ( .A(_51__0_), .Y(_173_) );
NAND2X1 NAND2X1_42 ( .A(_52__0_), .B(w_cout_8_), .Y(_174_) );
OAI21X1 OAI21X1_42 ( .A(w_cout_8_), .B(_173_), .C(_174_), .Y(_0__33_) );
INVX1 INVX1_43 ( .A(_51__1_), .Y(_175_) );
NAND2X1 NAND2X1_43 ( .A(w_cout_8_), .B(_52__1_), .Y(_176_) );
OAI21X1 OAI21X1_43 ( .A(w_cout_8_), .B(_175_), .C(_176_), .Y(_0__34_) );
INVX1 INVX1_44 ( .A(_51__2_), .Y(_177_) );
NAND2X1 NAND2X1_44 ( .A(w_cout_8_), .B(_52__2_), .Y(_178_) );
OAI21X1 OAI21X1_44 ( .A(w_cout_8_), .B(_177_), .C(_178_), .Y(_0__35_) );
INVX1 INVX1_45 ( .A(_51__3_), .Y(_179_) );
NAND2X1 NAND2X1_45 ( .A(w_cout_8_), .B(_52__3_), .Y(_180_) );
OAI21X1 OAI21X1_45 ( .A(w_cout_8_), .B(_179_), .C(_180_), .Y(_0__36_) );
INVX1 INVX1_46 ( .A(_55_), .Y(_181_) );
NAND2X1 NAND2X1_46 ( .A(_56_), .B(w_cout_9_), .Y(_182_) );
OAI21X1 OAI21X1_46 ( .A(w_cout_9_), .B(_181_), .C(_182_), .Y(w_cout_10_) );
INVX1 INVX1_47 ( .A(_57__0_), .Y(_183_) );
NAND2X1 NAND2X1_47 ( .A(_58__0_), .B(w_cout_9_), .Y(_184_) );
OAI21X1 OAI21X1_47 ( .A(w_cout_9_), .B(_183_), .C(_184_), .Y(_0__37_) );
INVX1 INVX1_48 ( .A(_57__1_), .Y(_185_) );
NAND2X1 NAND2X1_48 ( .A(w_cout_9_), .B(_58__1_), .Y(_186_) );
OAI21X1 OAI21X1_48 ( .A(w_cout_9_), .B(_185_), .C(_186_), .Y(_0__38_) );
INVX1 INVX1_49 ( .A(_57__2_), .Y(_187_) );
NAND2X1 NAND2X1_49 ( .A(w_cout_9_), .B(_58__2_), .Y(_188_) );
OAI21X1 OAI21X1_49 ( .A(w_cout_9_), .B(_187_), .C(_188_), .Y(_0__39_) );
INVX1 INVX1_50 ( .A(_57__3_), .Y(_189_) );
NAND2X1 NAND2X1_50 ( .A(w_cout_9_), .B(_58__3_), .Y(_190_) );
OAI21X1 OAI21X1_50 ( .A(w_cout_9_), .B(_189_), .C(_190_), .Y(_0__40_) );
INVX1 INVX1_51 ( .A(_61_), .Y(_191_) );
NAND2X1 NAND2X1_51 ( .A(_62_), .B(w_cout_10_), .Y(_192_) );
OAI21X1 OAI21X1_51 ( .A(w_cout_10_), .B(_191_), .C(_192_), .Y(w_cout_11_) );
INVX1 INVX1_52 ( .A(_63__0_), .Y(_193_) );
NAND2X1 NAND2X1_52 ( .A(_64__0_), .B(w_cout_10_), .Y(_194_) );
OAI21X1 OAI21X1_52 ( .A(w_cout_10_), .B(_193_), .C(_194_), .Y(_0__41_) );
INVX1 INVX1_53 ( .A(_63__1_), .Y(_195_) );
NAND2X1 NAND2X1_53 ( .A(w_cout_10_), .B(_64__1_), .Y(_196_) );
OAI21X1 OAI21X1_53 ( .A(w_cout_10_), .B(_195_), .C(_196_), .Y(_0__42_) );
INVX1 INVX1_54 ( .A(_63__2_), .Y(_197_) );
NAND2X1 NAND2X1_54 ( .A(w_cout_10_), .B(_64__2_), .Y(_198_) );
OAI21X1 OAI21X1_54 ( .A(w_cout_10_), .B(_197_), .C(_198_), .Y(_0__43_) );
INVX1 INVX1_55 ( .A(_63__3_), .Y(_199_) );
NAND2X1 NAND2X1_55 ( .A(w_cout_10_), .B(_64__3_), .Y(_200_) );
OAI21X1 OAI21X1_55 ( .A(w_cout_10_), .B(_199_), .C(_200_), .Y(_0__44_) );
INVX1 INVX1_56 ( .A(_67_), .Y(_201_) );
NAND2X1 NAND2X1_56 ( .A(_68_), .B(w_cout_11_), .Y(_202_) );
OAI21X1 OAI21X1_56 ( .A(w_cout_11_), .B(_201_), .C(_202_), .Y(w_cout_12_) );
INVX1 INVX1_57 ( .A(_69__0_), .Y(_203_) );
NAND2X1 NAND2X1_57 ( .A(_70__0_), .B(w_cout_11_), .Y(_204_) );
OAI21X1 OAI21X1_57 ( .A(w_cout_11_), .B(_203_), .C(_204_), .Y(_0__45_) );
INVX1 INVX1_58 ( .A(_69__1_), .Y(_205_) );
NAND2X1 NAND2X1_58 ( .A(w_cout_11_), .B(_70__1_), .Y(_206_) );
OAI21X1 OAI21X1_58 ( .A(w_cout_11_), .B(_205_), .C(_206_), .Y(_0__46_) );
INVX1 INVX1_59 ( .A(_69__2_), .Y(_207_) );
NAND2X1 NAND2X1_59 ( .A(w_cout_11_), .B(_70__2_), .Y(_208_) );
OAI21X1 OAI21X1_59 ( .A(w_cout_11_), .B(_207_), .C(_208_), .Y(_0__47_) );
INVX1 INVX1_60 ( .A(_69__3_), .Y(_209_) );
NAND2X1 NAND2X1_60 ( .A(w_cout_11_), .B(_70__3_), .Y(_210_) );
OAI21X1 OAI21X1_60 ( .A(w_cout_11_), .B(_209_), .C(_210_), .Y(_0__48_) );
INVX1 INVX1_61 ( .A(_73_), .Y(_211_) );
NAND2X1 NAND2X1_61 ( .A(_74_), .B(w_cout_12_), .Y(_212_) );
OAI21X1 OAI21X1_61 ( .A(w_cout_12_), .B(_211_), .C(_212_), .Y(w_cout_13_) );
INVX1 INVX1_62 ( .A(_75__0_), .Y(_213_) );
NAND2X1 NAND2X1_62 ( .A(_76__0_), .B(w_cout_12_), .Y(_214_) );
OAI21X1 OAI21X1_62 ( .A(w_cout_12_), .B(_213_), .C(_214_), .Y(_0__49_) );
INVX1 INVX1_63 ( .A(_75__1_), .Y(_215_) );
NAND2X1 NAND2X1_63 ( .A(w_cout_12_), .B(_76__1_), .Y(_216_) );
OAI21X1 OAI21X1_63 ( .A(w_cout_12_), .B(_215_), .C(_216_), .Y(_0__50_) );
INVX1 INVX1_64 ( .A(_75__2_), .Y(_217_) );
NAND2X1 NAND2X1_64 ( .A(w_cout_12_), .B(_76__2_), .Y(_218_) );
OAI21X1 OAI21X1_64 ( .A(w_cout_12_), .B(_217_), .C(_218_), .Y(_0__51_) );
INVX1 INVX1_65 ( .A(_75__3_), .Y(_219_) );
NAND2X1 NAND2X1_65 ( .A(w_cout_12_), .B(_76__3_), .Y(_220_) );
OAI21X1 OAI21X1_65 ( .A(w_cout_12_), .B(_219_), .C(_220_), .Y(_0__52_) );
INVX1 INVX1_66 ( .A(_79_), .Y(_221_) );
NAND2X1 NAND2X1_66 ( .A(_80_), .B(w_cout_13_), .Y(_222_) );
OAI21X1 OAI21X1_66 ( .A(w_cout_13_), .B(_221_), .C(_222_), .Y(w_cout_14_) );
INVX1 INVX1_67 ( .A(_81__0_), .Y(_223_) );
NAND2X1 NAND2X1_67 ( .A(_82__0_), .B(w_cout_13_), .Y(_224_) );
OAI21X1 OAI21X1_67 ( .A(w_cout_13_), .B(_223_), .C(_224_), .Y(_0__53_) );
INVX1 INVX1_68 ( .A(_81__1_), .Y(_225_) );
NAND2X1 NAND2X1_68 ( .A(w_cout_13_), .B(_82__1_), .Y(_226_) );
OAI21X1 OAI21X1_68 ( .A(w_cout_13_), .B(_225_), .C(_226_), .Y(_0__54_) );
INVX1 INVX1_69 ( .A(_81__2_), .Y(_227_) );
NAND2X1 NAND2X1_69 ( .A(w_cout_13_), .B(_82__2_), .Y(_228_) );
OAI21X1 OAI21X1_69 ( .A(w_cout_13_), .B(_227_), .C(_228_), .Y(_0__55_) );
INVX1 INVX1_70 ( .A(_81__3_), .Y(_229_) );
NAND2X1 NAND2X1_70 ( .A(w_cout_13_), .B(_82__3_), .Y(_230_) );
OAI21X1 OAI21X1_70 ( .A(w_cout_13_), .B(_229_), .C(_230_), .Y(_0__56_) );
INVX1 INVX1_71 ( .A(_85_), .Y(_231_) );
NAND2X1 NAND2X1_71 ( .A(_86_), .B(w_cout_14_), .Y(_232_) );
OAI21X1 OAI21X1_71 ( .A(w_cout_14_), .B(_231_), .C(_232_), .Y(w_cout_15_) );
INVX1 INVX1_72 ( .A(_87__0_), .Y(_233_) );
NAND2X1 NAND2X1_72 ( .A(_88__0_), .B(w_cout_14_), .Y(_234_) );
OAI21X1 OAI21X1_72 ( .A(w_cout_14_), .B(_233_), .C(_234_), .Y(_0__57_) );
INVX1 INVX1_73 ( .A(_87__1_), .Y(_235_) );
NAND2X1 NAND2X1_73 ( .A(w_cout_14_), .B(_88__1_), .Y(_236_) );
OAI21X1 OAI21X1_73 ( .A(w_cout_14_), .B(_235_), .C(_236_), .Y(_0__58_) );
INVX1 INVX1_74 ( .A(_87__2_), .Y(_237_) );
NAND2X1 NAND2X1_74 ( .A(w_cout_14_), .B(_88__2_), .Y(_238_) );
OAI21X1 OAI21X1_74 ( .A(w_cout_14_), .B(_237_), .C(_238_), .Y(_0__59_) );
INVX1 INVX1_75 ( .A(_87__3_), .Y(_239_) );
NAND2X1 NAND2X1_75 ( .A(w_cout_14_), .B(_88__3_), .Y(_240_) );
OAI21X1 OAI21X1_75 ( .A(w_cout_14_), .B(_239_), .C(_240_), .Y(_0__60_) );
INVX1 INVX1_76 ( .A(1'b0), .Y(_244_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_245_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_246_) );
NAND3X1 NAND3X1_1 ( .A(_244_), .B(_246_), .C(_245_), .Y(_247_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_241_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_242_) );
OAI21X1 OAI21X1_76 ( .A(_241_), .B(_242_), .C(1'b0), .Y(_243_) );
NAND2X1 NAND2X1_77 ( .A(_243_), .B(_247_), .Y(_3__0_) );
OAI21X1 OAI21X1_77 ( .A(_244_), .B(_241_), .C(_246_), .Y(_5__1_) );
INVX1 INVX1_77 ( .A(_5__1_), .Y(_251_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_252_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_253_) );
NAND3X1 NAND3X1_2 ( .A(_251_), .B(_253_), .C(_252_), .Y(_254_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_248_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_249_) );
OAI21X1 OAI21X1_78 ( .A(_248_), .B(_249_), .C(_5__1_), .Y(_250_) );
NAND2X1 NAND2X1_79 ( .A(_250_), .B(_254_), .Y(_3__1_) );
OAI21X1 OAI21X1_79 ( .A(_251_), .B(_248_), .C(_253_), .Y(_5__2_) );
INVX1 INVX1_78 ( .A(_5__2_), .Y(_258_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_259_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_260_) );
NAND3X1 NAND3X1_3 ( .A(_258_), .B(_260_), .C(_259_), .Y(_261_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_255_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_256_) );
OAI21X1 OAI21X1_80 ( .A(_255_), .B(_256_), .C(_5__2_), .Y(_257_) );
NAND2X1 NAND2X1_81 ( .A(_257_), .B(_261_), .Y(_3__2_) );
OAI21X1 OAI21X1_81 ( .A(_258_), .B(_255_), .C(_260_), .Y(_5__3_) );
INVX1 INVX1_79 ( .A(_5__3_), .Y(_265_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_266_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_267_) );
NAND3X1 NAND3X1_4 ( .A(_265_), .B(_267_), .C(_266_), .Y(_268_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_262_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_263_) );
OAI21X1 OAI21X1_82 ( .A(_262_), .B(_263_), .C(_5__3_), .Y(_264_) );
NAND2X1 NAND2X1_83 ( .A(_264_), .B(_268_), .Y(_3__3_) );
OAI21X1 OAI21X1_83 ( .A(_265_), .B(_262_), .C(_267_), .Y(_1_) );
INVX1 INVX1_80 ( .A(1'b1), .Y(_272_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_273_) );
NAND2X1 NAND2X1_84 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_274_) );
NAND3X1 NAND3X1_5 ( .A(_272_), .B(_274_), .C(_273_), .Y(_275_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_269_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_270_) );
OAI21X1 OAI21X1_84 ( .A(_269_), .B(_270_), .C(1'b1), .Y(_271_) );
NAND2X1 NAND2X1_85 ( .A(_271_), .B(_275_), .Y(_4__0_) );
OAI21X1 OAI21X1_85 ( .A(_272_), .B(_269_), .C(_274_), .Y(_6__1_) );
INVX1 INVX1_81 ( .A(_6__1_), .Y(_279_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_280_) );
NAND2X1 NAND2X1_86 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_281_) );
NAND3X1 NAND3X1_6 ( .A(_279_), .B(_281_), .C(_280_), .Y(_282_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_276_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_277_) );
OAI21X1 OAI21X1_86 ( .A(_276_), .B(_277_), .C(_6__1_), .Y(_278_) );
NAND2X1 NAND2X1_87 ( .A(_278_), .B(_282_), .Y(_4__1_) );
OAI21X1 OAI21X1_87 ( .A(_279_), .B(_276_), .C(_281_), .Y(_6__2_) );
INVX1 INVX1_82 ( .A(_6__2_), .Y(_286_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_287_) );
NAND2X1 NAND2X1_88 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_288_) );
NAND3X1 NAND3X1_7 ( .A(_286_), .B(_288_), .C(_287_), .Y(_289_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_283_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_284_) );
OAI21X1 OAI21X1_88 ( .A(_283_), .B(_284_), .C(_6__2_), .Y(_285_) );
NAND2X1 NAND2X1_89 ( .A(_285_), .B(_289_), .Y(_4__2_) );
OAI21X1 OAI21X1_89 ( .A(_286_), .B(_283_), .C(_288_), .Y(_6__3_) );
INVX1 INVX1_83 ( .A(_6__3_), .Y(_293_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_294_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_295_) );
NAND3X1 NAND3X1_8 ( .A(_293_), .B(_295_), .C(_294_), .Y(_296_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_290_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_291_) );
OAI21X1 OAI21X1_90 ( .A(_290_), .B(_291_), .C(_6__3_), .Y(_292_) );
NAND2X1 NAND2X1_91 ( .A(_292_), .B(_296_), .Y(_4__3_) );
OAI21X1 OAI21X1_91 ( .A(_293_), .B(_290_), .C(_295_), .Y(_2_) );
INVX1 INVX1_84 ( .A(1'b0), .Y(_300_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_301_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_302_) );
NAND3X1 NAND3X1_9 ( .A(_300_), .B(_302_), .C(_301_), .Y(_303_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_297_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_298_) );
OAI21X1 OAI21X1_92 ( .A(_297_), .B(_298_), .C(1'b0), .Y(_299_) );
NAND2X1 NAND2X1_93 ( .A(_299_), .B(_303_), .Y(_9__0_) );
OAI21X1 OAI21X1_93 ( .A(_300_), .B(_297_), .C(_302_), .Y(_11__1_) );
INVX1 INVX1_85 ( .A(_11__1_), .Y(_307_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_308_) );
NAND2X1 NAND2X1_94 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_309_) );
NAND3X1 NAND3X1_10 ( .A(_307_), .B(_309_), .C(_308_), .Y(_310_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_304_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_305_) );
OAI21X1 OAI21X1_94 ( .A(_304_), .B(_305_), .C(_11__1_), .Y(_306_) );
NAND2X1 NAND2X1_95 ( .A(_306_), .B(_310_), .Y(_9__1_) );
OAI21X1 OAI21X1_95 ( .A(_307_), .B(_304_), .C(_309_), .Y(_11__2_) );
INVX1 INVX1_86 ( .A(_11__2_), .Y(_314_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_315_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_316_) );
NAND3X1 NAND3X1_11 ( .A(_314_), .B(_316_), .C(_315_), .Y(_317_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_311_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_312_) );
OAI21X1 OAI21X1_96 ( .A(_311_), .B(_312_), .C(_11__2_), .Y(_313_) );
NAND2X1 NAND2X1_97 ( .A(_313_), .B(_317_), .Y(_9__2_) );
OAI21X1 OAI21X1_97 ( .A(_314_), .B(_311_), .C(_316_), .Y(_11__3_) );
INVX1 INVX1_87 ( .A(_11__3_), .Y(_321_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_322_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_323_) );
NAND3X1 NAND3X1_12 ( .A(_321_), .B(_323_), .C(_322_), .Y(_324_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_318_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_319_) );
OAI21X1 OAI21X1_98 ( .A(_318_), .B(_319_), .C(_11__3_), .Y(_320_) );
NAND2X1 NAND2X1_99 ( .A(_320_), .B(_324_), .Y(_9__3_) );
OAI21X1 OAI21X1_99 ( .A(_321_), .B(_318_), .C(_323_), .Y(_7_) );
INVX1 INVX1_88 ( .A(1'b1), .Y(_328_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_329_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_330_) );
NAND3X1 NAND3X1_13 ( .A(_328_), .B(_330_), .C(_329_), .Y(_331_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_325_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_326_) );
OAI21X1 OAI21X1_100 ( .A(_325_), .B(_326_), .C(1'b1), .Y(_327_) );
NAND2X1 NAND2X1_101 ( .A(_327_), .B(_331_), .Y(_10__0_) );
OAI21X1 OAI21X1_101 ( .A(_328_), .B(_325_), .C(_330_), .Y(_12__1_) );
INVX1 INVX1_89 ( .A(_12__1_), .Y(_335_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_336_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_337_) );
NAND3X1 NAND3X1_14 ( .A(_335_), .B(_337_), .C(_336_), .Y(_338_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_332_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_333_) );
OAI21X1 OAI21X1_102 ( .A(_332_), .B(_333_), .C(_12__1_), .Y(_334_) );
NAND2X1 NAND2X1_103 ( .A(_334_), .B(_338_), .Y(_10__1_) );
OAI21X1 OAI21X1_103 ( .A(_335_), .B(_332_), .C(_337_), .Y(_12__2_) );
INVX1 INVX1_90 ( .A(_12__2_), .Y(_342_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_343_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_344_) );
NAND3X1 NAND3X1_15 ( .A(_342_), .B(_344_), .C(_343_), .Y(_345_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_339_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_340_) );
OAI21X1 OAI21X1_104 ( .A(_339_), .B(_340_), .C(_12__2_), .Y(_341_) );
NAND2X1 NAND2X1_105 ( .A(_341_), .B(_345_), .Y(_10__2_) );
OAI21X1 OAI21X1_105 ( .A(_342_), .B(_339_), .C(_344_), .Y(_12__3_) );
INVX1 INVX1_91 ( .A(_12__3_), .Y(_349_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_350_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_351_) );
NAND3X1 NAND3X1_16 ( .A(_349_), .B(_351_), .C(_350_), .Y(_352_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_346_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_347_) );
OAI21X1 OAI21X1_106 ( .A(_346_), .B(_347_), .C(_12__3_), .Y(_348_) );
NAND2X1 NAND2X1_107 ( .A(_348_), .B(_352_), .Y(_10__3_) );
OAI21X1 OAI21X1_107 ( .A(_349_), .B(_346_), .C(_351_), .Y(_8_) );
INVX1 INVX1_92 ( .A(1'b0), .Y(_356_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_357_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_358_) );
NAND3X1 NAND3X1_17 ( .A(_356_), .B(_358_), .C(_357_), .Y(_359_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_353_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_354_) );
OAI21X1 OAI21X1_108 ( .A(_353_), .B(_354_), .C(1'b0), .Y(_355_) );
NAND2X1 NAND2X1_109 ( .A(_355_), .B(_359_), .Y(_15__0_) );
OAI21X1 OAI21X1_109 ( .A(_356_), .B(_353_), .C(_358_), .Y(_17__1_) );
INVX1 INVX1_93 ( .A(_17__1_), .Y(_363_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_364_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_365_) );
NAND3X1 NAND3X1_18 ( .A(_363_), .B(_365_), .C(_364_), .Y(_366_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_360_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_361_) );
OAI21X1 OAI21X1_110 ( .A(_360_), .B(_361_), .C(_17__1_), .Y(_362_) );
NAND2X1 NAND2X1_111 ( .A(_362_), .B(_366_), .Y(_15__1_) );
OAI21X1 OAI21X1_111 ( .A(_363_), .B(_360_), .C(_365_), .Y(_17__2_) );
INVX1 INVX1_94 ( .A(_17__2_), .Y(_370_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_371_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_372_) );
NAND3X1 NAND3X1_19 ( .A(_370_), .B(_372_), .C(_371_), .Y(_373_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_367_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_368_) );
OAI21X1 OAI21X1_112 ( .A(_367_), .B(_368_), .C(_17__2_), .Y(_369_) );
NAND2X1 NAND2X1_113 ( .A(_369_), .B(_373_), .Y(_15__2_) );
OAI21X1 OAI21X1_113 ( .A(_370_), .B(_367_), .C(_372_), .Y(_17__3_) );
INVX1 INVX1_95 ( .A(_17__3_), .Y(_377_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_378_) );
NAND2X1 NAND2X1_114 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_379_) );
NAND3X1 NAND3X1_20 ( .A(_377_), .B(_379_), .C(_378_), .Y(_380_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_374_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_375_) );
OAI21X1 OAI21X1_114 ( .A(_374_), .B(_375_), .C(_17__3_), .Y(_376_) );
NAND2X1 NAND2X1_115 ( .A(_376_), .B(_380_), .Y(_15__3_) );
OAI21X1 OAI21X1_115 ( .A(_377_), .B(_374_), .C(_379_), .Y(_13_) );
INVX1 INVX1_96 ( .A(1'b1), .Y(_384_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_385_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_386_) );
NAND3X1 NAND3X1_21 ( .A(_384_), .B(_386_), .C(_385_), .Y(_387_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_381_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_382_) );
OAI21X1 OAI21X1_116 ( .A(_381_), .B(_382_), .C(1'b1), .Y(_383_) );
NAND2X1 NAND2X1_117 ( .A(_383_), .B(_387_), .Y(_16__0_) );
OAI21X1 OAI21X1_117 ( .A(_384_), .B(_381_), .C(_386_), .Y(_18__1_) );
INVX1 INVX1_97 ( .A(_18__1_), .Y(_391_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_392_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_393_) );
NAND3X1 NAND3X1_22 ( .A(_391_), .B(_393_), .C(_392_), .Y(_394_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_388_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_389_) );
OAI21X1 OAI21X1_118 ( .A(_388_), .B(_389_), .C(_18__1_), .Y(_390_) );
NAND2X1 NAND2X1_119 ( .A(_390_), .B(_394_), .Y(_16__1_) );
OAI21X1 OAI21X1_119 ( .A(_391_), .B(_388_), .C(_393_), .Y(_18__2_) );
INVX1 INVX1_98 ( .A(_18__2_), .Y(_398_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_399_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_400_) );
NAND3X1 NAND3X1_23 ( .A(_398_), .B(_400_), .C(_399_), .Y(_401_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_395_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_396_) );
OAI21X1 OAI21X1_120 ( .A(_395_), .B(_396_), .C(_18__2_), .Y(_397_) );
NAND2X1 NAND2X1_121 ( .A(_397_), .B(_401_), .Y(_16__2_) );
OAI21X1 OAI21X1_121 ( .A(_398_), .B(_395_), .C(_400_), .Y(_18__3_) );
INVX1 INVX1_99 ( .A(_18__3_), .Y(_405_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_406_) );
NAND2X1 NAND2X1_122 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_407_) );
NAND3X1 NAND3X1_24 ( .A(_405_), .B(_407_), .C(_406_), .Y(_408_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_402_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_403_) );
OAI21X1 OAI21X1_122 ( .A(_402_), .B(_403_), .C(_18__3_), .Y(_404_) );
NAND2X1 NAND2X1_123 ( .A(_404_), .B(_408_), .Y(_16__3_) );
OAI21X1 OAI21X1_123 ( .A(_405_), .B(_402_), .C(_407_), .Y(_14_) );
INVX1 INVX1_100 ( .A(1'b0), .Y(_412_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_413_) );
NAND2X1 NAND2X1_124 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_414_) );
NAND3X1 NAND3X1_25 ( .A(_412_), .B(_414_), .C(_413_), .Y(_415_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_409_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_410_) );
OAI21X1 OAI21X1_124 ( .A(_409_), .B(_410_), .C(1'b0), .Y(_411_) );
NAND2X1 NAND2X1_125 ( .A(_411_), .B(_415_), .Y(_21__0_) );
OAI21X1 OAI21X1_125 ( .A(_412_), .B(_409_), .C(_414_), .Y(_23__1_) );
INVX1 INVX1_101 ( .A(_23__1_), .Y(_419_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_420_) );
NAND2X1 NAND2X1_126 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_421_) );
NAND3X1 NAND3X1_26 ( .A(_419_), .B(_421_), .C(_420_), .Y(_422_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_416_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_417_) );
OAI21X1 OAI21X1_126 ( .A(_416_), .B(_417_), .C(_23__1_), .Y(_418_) );
NAND2X1 NAND2X1_127 ( .A(_418_), .B(_422_), .Y(_21__1_) );
OAI21X1 OAI21X1_127 ( .A(_419_), .B(_416_), .C(_421_), .Y(_23__2_) );
INVX1 INVX1_102 ( .A(_23__2_), .Y(_426_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_427_) );
NAND2X1 NAND2X1_128 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_428_) );
NAND3X1 NAND3X1_27 ( .A(_426_), .B(_428_), .C(_427_), .Y(_429_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_423_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_424_) );
OAI21X1 OAI21X1_128 ( .A(_423_), .B(_424_), .C(_23__2_), .Y(_425_) );
NAND2X1 NAND2X1_129 ( .A(_425_), .B(_429_), .Y(_21__2_) );
OAI21X1 OAI21X1_129 ( .A(_426_), .B(_423_), .C(_428_), .Y(_23__3_) );
INVX1 INVX1_103 ( .A(_23__3_), .Y(_433_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_434_) );
NAND2X1 NAND2X1_130 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_435_) );
NAND3X1 NAND3X1_28 ( .A(_433_), .B(_435_), .C(_434_), .Y(_436_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_430_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_431_) );
OAI21X1 OAI21X1_130 ( .A(_430_), .B(_431_), .C(_23__3_), .Y(_432_) );
NAND2X1 NAND2X1_131 ( .A(_432_), .B(_436_), .Y(_21__3_) );
OAI21X1 OAI21X1_131 ( .A(_433_), .B(_430_), .C(_435_), .Y(_19_) );
INVX1 INVX1_104 ( .A(1'b1), .Y(_440_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_441_) );
NAND2X1 NAND2X1_132 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_442_) );
NAND3X1 NAND3X1_29 ( .A(_440_), .B(_442_), .C(_441_), .Y(_443_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_437_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_438_) );
OAI21X1 OAI21X1_132 ( .A(_437_), .B(_438_), .C(1'b1), .Y(_439_) );
NAND2X1 NAND2X1_133 ( .A(_439_), .B(_443_), .Y(_22__0_) );
OAI21X1 OAI21X1_133 ( .A(_440_), .B(_437_), .C(_442_), .Y(_24__1_) );
INVX1 INVX1_105 ( .A(_24__1_), .Y(_447_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_448_) );
NAND2X1 NAND2X1_134 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_449_) );
NAND3X1 NAND3X1_30 ( .A(_447_), .B(_449_), .C(_448_), .Y(_450_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_444_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_445_) );
OAI21X1 OAI21X1_134 ( .A(_444_), .B(_445_), .C(_24__1_), .Y(_446_) );
NAND2X1 NAND2X1_135 ( .A(_446_), .B(_450_), .Y(_22__1_) );
OAI21X1 OAI21X1_135 ( .A(_447_), .B(_444_), .C(_449_), .Y(_24__2_) );
INVX1 INVX1_106 ( .A(_24__2_), .Y(_454_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_455_) );
NAND2X1 NAND2X1_136 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_456_) );
NAND3X1 NAND3X1_31 ( .A(_454_), .B(_456_), .C(_455_), .Y(_457_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_451_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_452_) );
OAI21X1 OAI21X1_136 ( .A(_451_), .B(_452_), .C(_24__2_), .Y(_453_) );
NAND2X1 NAND2X1_137 ( .A(_453_), .B(_457_), .Y(_22__2_) );
OAI21X1 OAI21X1_137 ( .A(_454_), .B(_451_), .C(_456_), .Y(_24__3_) );
INVX1 INVX1_107 ( .A(_24__3_), .Y(_461_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_462_) );
NAND2X1 NAND2X1_138 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_463_) );
NAND3X1 NAND3X1_32 ( .A(_461_), .B(_463_), .C(_462_), .Y(_464_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_458_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_459_) );
OAI21X1 OAI21X1_138 ( .A(_458_), .B(_459_), .C(_24__3_), .Y(_460_) );
NAND2X1 NAND2X1_139 ( .A(_460_), .B(_464_), .Y(_22__3_) );
OAI21X1 OAI21X1_139 ( .A(_461_), .B(_458_), .C(_463_), .Y(_20_) );
INVX1 INVX1_108 ( .A(1'b0), .Y(_468_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_469_) );
NAND2X1 NAND2X1_140 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_470_) );
NAND3X1 NAND3X1_33 ( .A(_468_), .B(_470_), .C(_469_), .Y(_471_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_465_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_466_) );
OAI21X1 OAI21X1_140 ( .A(_465_), .B(_466_), .C(1'b0), .Y(_467_) );
NAND2X1 NAND2X1_141 ( .A(_467_), .B(_471_), .Y(_27__0_) );
OAI21X1 OAI21X1_141 ( .A(_468_), .B(_465_), .C(_470_), .Y(_29__1_) );
INVX1 INVX1_109 ( .A(_29__1_), .Y(_475_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_476_) );
NAND2X1 NAND2X1_142 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_477_) );
NAND3X1 NAND3X1_34 ( .A(_475_), .B(_477_), .C(_476_), .Y(_478_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_472_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_473_) );
OAI21X1 OAI21X1_142 ( .A(_472_), .B(_473_), .C(_29__1_), .Y(_474_) );
NAND2X1 NAND2X1_143 ( .A(_474_), .B(_478_), .Y(_27__1_) );
OAI21X1 OAI21X1_143 ( .A(_475_), .B(_472_), .C(_477_), .Y(_29__2_) );
INVX1 INVX1_110 ( .A(_29__2_), .Y(_482_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_483_) );
NAND2X1 NAND2X1_144 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_484_) );
NAND3X1 NAND3X1_35 ( .A(_482_), .B(_484_), .C(_483_), .Y(_485_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_479_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_480_) );
OAI21X1 OAI21X1_144 ( .A(_479_), .B(_480_), .C(_29__2_), .Y(_481_) );
NAND2X1 NAND2X1_145 ( .A(_481_), .B(_485_), .Y(_27__2_) );
OAI21X1 OAI21X1_145 ( .A(_482_), .B(_479_), .C(_484_), .Y(_29__3_) );
INVX1 INVX1_111 ( .A(_29__3_), .Y(_489_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_490_) );
NAND2X1 NAND2X1_146 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_491_) );
NAND3X1 NAND3X1_36 ( .A(_489_), .B(_491_), .C(_490_), .Y(_492_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_486_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_487_) );
OAI21X1 OAI21X1_146 ( .A(_486_), .B(_487_), .C(_29__3_), .Y(_488_) );
NAND2X1 NAND2X1_147 ( .A(_488_), .B(_492_), .Y(_27__3_) );
OAI21X1 OAI21X1_147 ( .A(_489_), .B(_486_), .C(_491_), .Y(_25_) );
INVX1 INVX1_112 ( .A(1'b1), .Y(_496_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_497_) );
NAND2X1 NAND2X1_148 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_498_) );
NAND3X1 NAND3X1_37 ( .A(_496_), .B(_498_), .C(_497_), .Y(_499_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_493_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_494_) );
OAI21X1 OAI21X1_148 ( .A(_493_), .B(_494_), .C(1'b1), .Y(_495_) );
NAND2X1 NAND2X1_149 ( .A(_495_), .B(_499_), .Y(_28__0_) );
OAI21X1 OAI21X1_149 ( .A(_496_), .B(_493_), .C(_498_), .Y(_30__1_) );
INVX1 INVX1_113 ( .A(_30__1_), .Y(_503_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_504_) );
NAND2X1 NAND2X1_150 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_505_) );
NAND3X1 NAND3X1_38 ( .A(_503_), .B(_505_), .C(_504_), .Y(_506_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_500_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_501_) );
OAI21X1 OAI21X1_150 ( .A(_500_), .B(_501_), .C(_30__1_), .Y(_502_) );
NAND2X1 NAND2X1_151 ( .A(_502_), .B(_506_), .Y(_28__1_) );
OAI21X1 OAI21X1_151 ( .A(_503_), .B(_500_), .C(_505_), .Y(_30__2_) );
INVX1 INVX1_114 ( .A(_30__2_), .Y(_510_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_511_) );
NAND2X1 NAND2X1_152 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_512_) );
NAND3X1 NAND3X1_39 ( .A(_510_), .B(_512_), .C(_511_), .Y(_513_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_507_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_508_) );
OAI21X1 OAI21X1_152 ( .A(_507_), .B(_508_), .C(_30__2_), .Y(_509_) );
NAND2X1 NAND2X1_153 ( .A(_509_), .B(_513_), .Y(_28__2_) );
OAI21X1 OAI21X1_153 ( .A(_510_), .B(_507_), .C(_512_), .Y(_30__3_) );
INVX1 INVX1_115 ( .A(_30__3_), .Y(_517_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_518_) );
NAND2X1 NAND2X1_154 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_519_) );
NAND3X1 NAND3X1_40 ( .A(_517_), .B(_519_), .C(_518_), .Y(_520_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_514_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_515_) );
OAI21X1 OAI21X1_154 ( .A(_514_), .B(_515_), .C(_30__3_), .Y(_516_) );
NAND2X1 NAND2X1_155 ( .A(_516_), .B(_520_), .Y(_28__3_) );
OAI21X1 OAI21X1_155 ( .A(_517_), .B(_514_), .C(_519_), .Y(_26_) );
INVX1 INVX1_116 ( .A(1'b0), .Y(_524_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_525_) );
NAND2X1 NAND2X1_156 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_526_) );
NAND3X1 NAND3X1_41 ( .A(_524_), .B(_526_), .C(_525_), .Y(_527_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_521_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_522_) );
OAI21X1 OAI21X1_156 ( .A(_521_), .B(_522_), .C(1'b0), .Y(_523_) );
NAND2X1 NAND2X1_157 ( .A(_523_), .B(_527_), .Y(_33__0_) );
OAI21X1 OAI21X1_157 ( .A(_524_), .B(_521_), .C(_526_), .Y(_35__1_) );
INVX1 INVX1_117 ( .A(_35__1_), .Y(_531_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_532_) );
NAND2X1 NAND2X1_158 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_533_) );
NAND3X1 NAND3X1_42 ( .A(_531_), .B(_533_), .C(_532_), .Y(_534_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_528_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_529_) );
OAI21X1 OAI21X1_158 ( .A(_528_), .B(_529_), .C(_35__1_), .Y(_530_) );
NAND2X1 NAND2X1_159 ( .A(_530_), .B(_534_), .Y(_33__1_) );
OAI21X1 OAI21X1_159 ( .A(_531_), .B(_528_), .C(_533_), .Y(_35__2_) );
INVX1 INVX1_118 ( .A(_35__2_), .Y(_538_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_539_) );
NAND2X1 NAND2X1_160 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_540_) );
NAND3X1 NAND3X1_43 ( .A(_538_), .B(_540_), .C(_539_), .Y(_541_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_535_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_536_) );
OAI21X1 OAI21X1_160 ( .A(_535_), .B(_536_), .C(_35__2_), .Y(_537_) );
NAND2X1 NAND2X1_161 ( .A(_537_), .B(_541_), .Y(_33__2_) );
OAI21X1 OAI21X1_161 ( .A(_538_), .B(_535_), .C(_540_), .Y(_35__3_) );
INVX1 INVX1_119 ( .A(_35__3_), .Y(_545_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_546_) );
NAND2X1 NAND2X1_162 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_547_) );
NAND3X1 NAND3X1_44 ( .A(_545_), .B(_547_), .C(_546_), .Y(_548_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_542_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_543_) );
OAI21X1 OAI21X1_162 ( .A(_542_), .B(_543_), .C(_35__3_), .Y(_544_) );
NAND2X1 NAND2X1_163 ( .A(_544_), .B(_548_), .Y(_33__3_) );
OAI21X1 OAI21X1_163 ( .A(_545_), .B(_542_), .C(_547_), .Y(_31_) );
INVX1 INVX1_120 ( .A(1'b1), .Y(_552_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_553_) );
NAND2X1 NAND2X1_164 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_554_) );
NAND3X1 NAND3X1_45 ( .A(_552_), .B(_554_), .C(_553_), .Y(_555_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_549_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_550_) );
OAI21X1 OAI21X1_164 ( .A(_549_), .B(_550_), .C(1'b1), .Y(_551_) );
NAND2X1 NAND2X1_165 ( .A(_551_), .B(_555_), .Y(_34__0_) );
OAI21X1 OAI21X1_165 ( .A(_552_), .B(_549_), .C(_554_), .Y(_36__1_) );
INVX1 INVX1_121 ( .A(_36__1_), .Y(_559_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_560_) );
NAND2X1 NAND2X1_166 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_561_) );
NAND3X1 NAND3X1_46 ( .A(_559_), .B(_561_), .C(_560_), .Y(_562_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_556_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_557_) );
OAI21X1 OAI21X1_166 ( .A(_556_), .B(_557_), .C(_36__1_), .Y(_558_) );
NAND2X1 NAND2X1_167 ( .A(_558_), .B(_562_), .Y(_34__1_) );
OAI21X1 OAI21X1_167 ( .A(_559_), .B(_556_), .C(_561_), .Y(_36__2_) );
INVX1 INVX1_122 ( .A(_36__2_), .Y(_566_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_567_) );
NAND2X1 NAND2X1_168 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_568_) );
NAND3X1 NAND3X1_47 ( .A(_566_), .B(_568_), .C(_567_), .Y(_569_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_563_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_564_) );
OAI21X1 OAI21X1_168 ( .A(_563_), .B(_564_), .C(_36__2_), .Y(_565_) );
NAND2X1 NAND2X1_169 ( .A(_565_), .B(_569_), .Y(_34__2_) );
OAI21X1 OAI21X1_169 ( .A(_566_), .B(_563_), .C(_568_), .Y(_36__3_) );
INVX1 INVX1_123 ( .A(_36__3_), .Y(_573_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_574_) );
NAND2X1 NAND2X1_170 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_575_) );
NAND3X1 NAND3X1_48 ( .A(_573_), .B(_575_), .C(_574_), .Y(_576_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_570_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_571_) );
OAI21X1 OAI21X1_170 ( .A(_570_), .B(_571_), .C(_36__3_), .Y(_572_) );
NAND2X1 NAND2X1_171 ( .A(_572_), .B(_576_), .Y(_34__3_) );
OAI21X1 OAI21X1_171 ( .A(_573_), .B(_570_), .C(_575_), .Y(_32_) );
INVX1 INVX1_124 ( .A(1'b0), .Y(_580_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_581_) );
NAND2X1 NAND2X1_172 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_582_) );
NAND3X1 NAND3X1_49 ( .A(_580_), .B(_582_), .C(_581_), .Y(_583_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_577_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_578_) );
OAI21X1 OAI21X1_172 ( .A(_577_), .B(_578_), .C(1'b0), .Y(_579_) );
NAND2X1 NAND2X1_173 ( .A(_579_), .B(_583_), .Y(_39__0_) );
OAI21X1 OAI21X1_173 ( .A(_580_), .B(_577_), .C(_582_), .Y(_41__1_) );
INVX1 INVX1_125 ( .A(_41__1_), .Y(_587_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_588_) );
NAND2X1 NAND2X1_174 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_589_) );
NAND3X1 NAND3X1_50 ( .A(_587_), .B(_589_), .C(_588_), .Y(_590_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_584_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_585_) );
OAI21X1 OAI21X1_174 ( .A(_584_), .B(_585_), .C(_41__1_), .Y(_586_) );
NAND2X1 NAND2X1_175 ( .A(_586_), .B(_590_), .Y(_39__1_) );
OAI21X1 OAI21X1_175 ( .A(_587_), .B(_584_), .C(_589_), .Y(_41__2_) );
INVX1 INVX1_126 ( .A(_41__2_), .Y(_594_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_595_) );
NAND2X1 NAND2X1_176 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_596_) );
NAND3X1 NAND3X1_51 ( .A(_594_), .B(_596_), .C(_595_), .Y(_597_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_591_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_592_) );
OAI21X1 OAI21X1_176 ( .A(_591_), .B(_592_), .C(_41__2_), .Y(_593_) );
NAND2X1 NAND2X1_177 ( .A(_593_), .B(_597_), .Y(_39__2_) );
OAI21X1 OAI21X1_177 ( .A(_594_), .B(_591_), .C(_596_), .Y(_41__3_) );
INVX1 INVX1_127 ( .A(_41__3_), .Y(_601_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_602_) );
NAND2X1 NAND2X1_178 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_603_) );
NAND3X1 NAND3X1_52 ( .A(_601_), .B(_603_), .C(_602_), .Y(_604_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_598_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_599_) );
OAI21X1 OAI21X1_178 ( .A(_598_), .B(_599_), .C(_41__3_), .Y(_600_) );
NAND2X1 NAND2X1_179 ( .A(_600_), .B(_604_), .Y(_39__3_) );
OAI21X1 OAI21X1_179 ( .A(_601_), .B(_598_), .C(_603_), .Y(_37_) );
INVX1 INVX1_128 ( .A(1'b1), .Y(_608_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_609_) );
NAND2X1 NAND2X1_180 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_610_) );
NAND3X1 NAND3X1_53 ( .A(_608_), .B(_610_), .C(_609_), .Y(_611_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_605_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_606_) );
OAI21X1 OAI21X1_180 ( .A(_605_), .B(_606_), .C(1'b1), .Y(_607_) );
NAND2X1 NAND2X1_181 ( .A(_607_), .B(_611_), .Y(_40__0_) );
OAI21X1 OAI21X1_181 ( .A(_608_), .B(_605_), .C(_610_), .Y(_42__1_) );
INVX1 INVX1_129 ( .A(_42__1_), .Y(_615_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_616_) );
NAND2X1 NAND2X1_182 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_617_) );
NAND3X1 NAND3X1_54 ( .A(_615_), .B(_617_), .C(_616_), .Y(_618_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_612_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_613_) );
OAI21X1 OAI21X1_182 ( .A(_612_), .B(_613_), .C(_42__1_), .Y(_614_) );
NAND2X1 NAND2X1_183 ( .A(_614_), .B(_618_), .Y(_40__1_) );
OAI21X1 OAI21X1_183 ( .A(_615_), .B(_612_), .C(_617_), .Y(_42__2_) );
INVX1 INVX1_130 ( .A(_42__2_), .Y(_622_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_623_) );
NAND2X1 NAND2X1_184 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_624_) );
NAND3X1 NAND3X1_55 ( .A(_622_), .B(_624_), .C(_623_), .Y(_625_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_619_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_620_) );
OAI21X1 OAI21X1_184 ( .A(_619_), .B(_620_), .C(_42__2_), .Y(_621_) );
NAND2X1 NAND2X1_185 ( .A(_621_), .B(_625_), .Y(_40__2_) );
OAI21X1 OAI21X1_185 ( .A(_622_), .B(_619_), .C(_624_), .Y(_42__3_) );
INVX1 INVX1_131 ( .A(_42__3_), .Y(_629_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_630_) );
NAND2X1 NAND2X1_186 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_631_) );
NAND3X1 NAND3X1_56 ( .A(_629_), .B(_631_), .C(_630_), .Y(_632_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_626_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_627_) );
OAI21X1 OAI21X1_186 ( .A(_626_), .B(_627_), .C(_42__3_), .Y(_628_) );
NAND2X1 NAND2X1_187 ( .A(_628_), .B(_632_), .Y(_40__3_) );
OAI21X1 OAI21X1_187 ( .A(_629_), .B(_626_), .C(_631_), .Y(_38_) );
INVX1 INVX1_132 ( .A(1'b0), .Y(_636_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_637_) );
NAND2X1 NAND2X1_188 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_638_) );
NAND3X1 NAND3X1_57 ( .A(_636_), .B(_638_), .C(_637_), .Y(_639_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_633_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_634_) );
OAI21X1 OAI21X1_188 ( .A(_633_), .B(_634_), .C(1'b0), .Y(_635_) );
NAND2X1 NAND2X1_189 ( .A(_635_), .B(_639_), .Y(_45__0_) );
OAI21X1 OAI21X1_189 ( .A(_636_), .B(_633_), .C(_638_), .Y(_47__1_) );
INVX1 INVX1_133 ( .A(_47__1_), .Y(_643_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_644_) );
NAND2X1 NAND2X1_190 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_645_) );
NAND3X1 NAND3X1_58 ( .A(_643_), .B(_645_), .C(_644_), .Y(_646_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_640_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_641_) );
OAI21X1 OAI21X1_190 ( .A(_640_), .B(_641_), .C(_47__1_), .Y(_642_) );
NAND2X1 NAND2X1_191 ( .A(_642_), .B(_646_), .Y(_45__1_) );
OAI21X1 OAI21X1_191 ( .A(_643_), .B(_640_), .C(_645_), .Y(_47__2_) );
INVX1 INVX1_134 ( .A(_47__2_), .Y(_650_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_651_) );
NAND2X1 NAND2X1_192 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_652_) );
NAND3X1 NAND3X1_59 ( .A(_650_), .B(_652_), .C(_651_), .Y(_653_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_647_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_648_) );
OAI21X1 OAI21X1_192 ( .A(_647_), .B(_648_), .C(_47__2_), .Y(_649_) );
NAND2X1 NAND2X1_193 ( .A(_649_), .B(_653_), .Y(_45__2_) );
OAI21X1 OAI21X1_193 ( .A(_650_), .B(_647_), .C(_652_), .Y(_47__3_) );
INVX1 INVX1_135 ( .A(_47__3_), .Y(_657_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_658_) );
NAND2X1 NAND2X1_194 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_659_) );
NAND3X1 NAND3X1_60 ( .A(_657_), .B(_659_), .C(_658_), .Y(_660_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_654_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_655_) );
OAI21X1 OAI21X1_194 ( .A(_654_), .B(_655_), .C(_47__3_), .Y(_656_) );
NAND2X1 NAND2X1_195 ( .A(_656_), .B(_660_), .Y(_45__3_) );
OAI21X1 OAI21X1_195 ( .A(_657_), .B(_654_), .C(_659_), .Y(_43_) );
INVX1 INVX1_136 ( .A(1'b1), .Y(_664_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_665_) );
NAND2X1 NAND2X1_196 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_666_) );
NAND3X1 NAND3X1_61 ( .A(_664_), .B(_666_), .C(_665_), .Y(_667_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_661_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_662_) );
OAI21X1 OAI21X1_196 ( .A(_661_), .B(_662_), .C(1'b1), .Y(_663_) );
NAND2X1 NAND2X1_197 ( .A(_663_), .B(_667_), .Y(_46__0_) );
OAI21X1 OAI21X1_197 ( .A(_664_), .B(_661_), .C(_666_), .Y(_48__1_) );
INVX1 INVX1_137 ( .A(_48__1_), .Y(_671_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_672_) );
NAND2X1 NAND2X1_198 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_673_) );
NAND3X1 NAND3X1_62 ( .A(_671_), .B(_673_), .C(_672_), .Y(_674_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_668_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_669_) );
OAI21X1 OAI21X1_198 ( .A(_668_), .B(_669_), .C(_48__1_), .Y(_670_) );
NAND2X1 NAND2X1_199 ( .A(_670_), .B(_674_), .Y(_46__1_) );
OAI21X1 OAI21X1_199 ( .A(_671_), .B(_668_), .C(_673_), .Y(_48__2_) );
INVX1 INVX1_138 ( .A(_48__2_), .Y(_678_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_679_) );
NAND2X1 NAND2X1_200 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_680_) );
NAND3X1 NAND3X1_63 ( .A(_678_), .B(_680_), .C(_679_), .Y(_681_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_675_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_676_) );
OAI21X1 OAI21X1_200 ( .A(_675_), .B(_676_), .C(_48__2_), .Y(_677_) );
NAND2X1 NAND2X1_201 ( .A(_677_), .B(_681_), .Y(_46__2_) );
OAI21X1 OAI21X1_201 ( .A(_678_), .B(_675_), .C(_680_), .Y(_48__3_) );
INVX1 INVX1_139 ( .A(_48__3_), .Y(_685_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_686_) );
NAND2X1 NAND2X1_202 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_687_) );
NAND3X1 NAND3X1_64 ( .A(_685_), .B(_687_), .C(_686_), .Y(_688_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_682_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_683_) );
OAI21X1 OAI21X1_202 ( .A(_682_), .B(_683_), .C(_48__3_), .Y(_684_) );
NAND2X1 NAND2X1_203 ( .A(_684_), .B(_688_), .Y(_46__3_) );
OAI21X1 OAI21X1_203 ( .A(_685_), .B(_682_), .C(_687_), .Y(_44_) );
INVX1 INVX1_140 ( .A(1'b0), .Y(_692_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_693_) );
NAND2X1 NAND2X1_204 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_694_) );
NAND3X1 NAND3X1_65 ( .A(_692_), .B(_694_), .C(_693_), .Y(_695_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_689_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_690_) );
OAI21X1 OAI21X1_204 ( .A(_689_), .B(_690_), .C(1'b0), .Y(_691_) );
NAND2X1 NAND2X1_205 ( .A(_691_), .B(_695_), .Y(_51__0_) );
OAI21X1 OAI21X1_205 ( .A(_692_), .B(_689_), .C(_694_), .Y(_53__1_) );
INVX1 INVX1_141 ( .A(_53__1_), .Y(_699_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_700_) );
NAND2X1 NAND2X1_206 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_701_) );
NAND3X1 NAND3X1_66 ( .A(_699_), .B(_701_), .C(_700_), .Y(_702_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_696_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_697_) );
OAI21X1 OAI21X1_206 ( .A(_696_), .B(_697_), .C(_53__1_), .Y(_698_) );
NAND2X1 NAND2X1_207 ( .A(_698_), .B(_702_), .Y(_51__1_) );
OAI21X1 OAI21X1_207 ( .A(_699_), .B(_696_), .C(_701_), .Y(_53__2_) );
INVX1 INVX1_142 ( .A(_53__2_), .Y(_706_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_707_) );
NAND2X1 NAND2X1_208 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_708_) );
NAND3X1 NAND3X1_67 ( .A(_706_), .B(_708_), .C(_707_), .Y(_709_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_703_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_704_) );
OAI21X1 OAI21X1_208 ( .A(_703_), .B(_704_), .C(_53__2_), .Y(_705_) );
NAND2X1 NAND2X1_209 ( .A(_705_), .B(_709_), .Y(_51__2_) );
OAI21X1 OAI21X1_209 ( .A(_706_), .B(_703_), .C(_708_), .Y(_53__3_) );
INVX1 INVX1_143 ( .A(_53__3_), .Y(_713_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_714_) );
NAND2X1 NAND2X1_210 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_715_) );
NAND3X1 NAND3X1_68 ( .A(_713_), .B(_715_), .C(_714_), .Y(_716_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_710_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_711_) );
OAI21X1 OAI21X1_210 ( .A(_710_), .B(_711_), .C(_53__3_), .Y(_712_) );
NAND2X1 NAND2X1_211 ( .A(_712_), .B(_716_), .Y(_51__3_) );
OAI21X1 OAI21X1_211 ( .A(_713_), .B(_710_), .C(_715_), .Y(_49_) );
INVX1 INVX1_144 ( .A(1'b1), .Y(_720_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_721_) );
NAND2X1 NAND2X1_212 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_722_) );
NAND3X1 NAND3X1_69 ( .A(_720_), .B(_722_), .C(_721_), .Y(_723_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_717_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_718_) );
OAI21X1 OAI21X1_212 ( .A(_717_), .B(_718_), .C(1'b1), .Y(_719_) );
NAND2X1 NAND2X1_213 ( .A(_719_), .B(_723_), .Y(_52__0_) );
OAI21X1 OAI21X1_213 ( .A(_720_), .B(_717_), .C(_722_), .Y(_54__1_) );
INVX1 INVX1_145 ( .A(_54__1_), .Y(_727_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_728_) );
NAND2X1 NAND2X1_214 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_729_) );
NAND3X1 NAND3X1_70 ( .A(_727_), .B(_729_), .C(_728_), .Y(_730_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_724_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_725_) );
OAI21X1 OAI21X1_214 ( .A(_724_), .B(_725_), .C(_54__1_), .Y(_726_) );
NAND2X1 NAND2X1_215 ( .A(_726_), .B(_730_), .Y(_52__1_) );
OAI21X1 OAI21X1_215 ( .A(_727_), .B(_724_), .C(_729_), .Y(_54__2_) );
INVX1 INVX1_146 ( .A(_54__2_), .Y(_734_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_735_) );
NAND2X1 NAND2X1_216 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_736_) );
NAND3X1 NAND3X1_71 ( .A(_734_), .B(_736_), .C(_735_), .Y(_737_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_731_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_732_) );
OAI21X1 OAI21X1_216 ( .A(_731_), .B(_732_), .C(_54__2_), .Y(_733_) );
NAND2X1 NAND2X1_217 ( .A(_733_), .B(_737_), .Y(_52__2_) );
OAI21X1 OAI21X1_217 ( .A(_734_), .B(_731_), .C(_736_), .Y(_54__3_) );
INVX1 INVX1_147 ( .A(_54__3_), .Y(_741_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_742_) );
NAND2X1 NAND2X1_218 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_743_) );
NAND3X1 NAND3X1_72 ( .A(_741_), .B(_743_), .C(_742_), .Y(_744_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_738_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_739_) );
OAI21X1 OAI21X1_218 ( .A(_738_), .B(_739_), .C(_54__3_), .Y(_740_) );
NAND2X1 NAND2X1_219 ( .A(_740_), .B(_744_), .Y(_52__3_) );
OAI21X1 OAI21X1_219 ( .A(_741_), .B(_738_), .C(_743_), .Y(_50_) );
INVX1 INVX1_148 ( .A(1'b0), .Y(_748_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_749_) );
NAND2X1 NAND2X1_220 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_750_) );
NAND3X1 NAND3X1_73 ( .A(_748_), .B(_750_), .C(_749_), .Y(_751_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_745_) );
AND2X2 AND2X2_73 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_746_) );
OAI21X1 OAI21X1_220 ( .A(_745_), .B(_746_), .C(1'b0), .Y(_747_) );
NAND2X1 NAND2X1_221 ( .A(_747_), .B(_751_), .Y(_57__0_) );
OAI21X1 OAI21X1_221 ( .A(_748_), .B(_745_), .C(_750_), .Y(_59__1_) );
INVX1 INVX1_149 ( .A(_59__1_), .Y(_755_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_756_) );
NAND2X1 NAND2X1_222 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_757_) );
NAND3X1 NAND3X1_74 ( .A(_755_), .B(_757_), .C(_756_), .Y(_758_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_752_) );
AND2X2 AND2X2_74 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_753_) );
OAI21X1 OAI21X1_222 ( .A(_752_), .B(_753_), .C(_59__1_), .Y(_754_) );
NAND2X1 NAND2X1_223 ( .A(_754_), .B(_758_), .Y(_57__1_) );
OAI21X1 OAI21X1_223 ( .A(_755_), .B(_752_), .C(_757_), .Y(_59__2_) );
INVX1 INVX1_150 ( .A(_59__2_), .Y(_762_) );
OR2X2 OR2X2_75 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_763_) );
NAND2X1 NAND2X1_224 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_764_) );
NAND3X1 NAND3X1_75 ( .A(_762_), .B(_764_), .C(_763_), .Y(_765_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_759_) );
AND2X2 AND2X2_75 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_760_) );
OAI21X1 OAI21X1_224 ( .A(_759_), .B(_760_), .C(_59__2_), .Y(_761_) );
NAND2X1 NAND2X1_225 ( .A(_761_), .B(_765_), .Y(_57__2_) );
OAI21X1 OAI21X1_225 ( .A(_762_), .B(_759_), .C(_764_), .Y(_59__3_) );
INVX1 INVX1_151 ( .A(_59__3_), .Y(_769_) );
OR2X2 OR2X2_76 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_770_) );
NAND2X1 NAND2X1_226 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_771_) );
NAND3X1 NAND3X1_76 ( .A(_769_), .B(_771_), .C(_770_), .Y(_772_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_766_) );
AND2X2 AND2X2_76 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_767_) );
OAI21X1 OAI21X1_226 ( .A(_766_), .B(_767_), .C(_59__3_), .Y(_768_) );
NAND2X1 NAND2X1_227 ( .A(_768_), .B(_772_), .Y(_57__3_) );
OAI21X1 OAI21X1_227 ( .A(_769_), .B(_766_), .C(_771_), .Y(_55_) );
INVX1 INVX1_152 ( .A(1'b1), .Y(_776_) );
OR2X2 OR2X2_77 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_777_) );
NAND2X1 NAND2X1_228 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_778_) );
NAND3X1 NAND3X1_77 ( .A(_776_), .B(_778_), .C(_777_), .Y(_779_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_773_) );
AND2X2 AND2X2_77 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_774_) );
OAI21X1 OAI21X1_228 ( .A(_773_), .B(_774_), .C(1'b1), .Y(_775_) );
NAND2X1 NAND2X1_229 ( .A(_775_), .B(_779_), .Y(_58__0_) );
OAI21X1 OAI21X1_229 ( .A(_776_), .B(_773_), .C(_778_), .Y(_60__1_) );
INVX1 INVX1_153 ( .A(_60__1_), .Y(_783_) );
OR2X2 OR2X2_78 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_784_) );
NAND2X1 NAND2X1_230 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_785_) );
NAND3X1 NAND3X1_78 ( .A(_783_), .B(_785_), .C(_784_), .Y(_786_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_780_) );
AND2X2 AND2X2_78 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_781_) );
OAI21X1 OAI21X1_230 ( .A(_780_), .B(_781_), .C(_60__1_), .Y(_782_) );
NAND2X1 NAND2X1_231 ( .A(_782_), .B(_786_), .Y(_58__1_) );
OAI21X1 OAI21X1_231 ( .A(_783_), .B(_780_), .C(_785_), .Y(_60__2_) );
INVX1 INVX1_154 ( .A(_60__2_), .Y(_790_) );
OR2X2 OR2X2_79 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_791_) );
NAND2X1 NAND2X1_232 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_792_) );
NAND3X1 NAND3X1_79 ( .A(_790_), .B(_792_), .C(_791_), .Y(_793_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_787_) );
AND2X2 AND2X2_79 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_788_) );
OAI21X1 OAI21X1_232 ( .A(_787_), .B(_788_), .C(_60__2_), .Y(_789_) );
NAND2X1 NAND2X1_233 ( .A(_789_), .B(_793_), .Y(_58__2_) );
OAI21X1 OAI21X1_233 ( .A(_790_), .B(_787_), .C(_792_), .Y(_60__3_) );
INVX1 INVX1_155 ( .A(_60__3_), .Y(_797_) );
OR2X2 OR2X2_80 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_798_) );
NAND2X1 NAND2X1_234 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_799_) );
NAND3X1 NAND3X1_80 ( .A(_797_), .B(_799_), .C(_798_), .Y(_800_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_794_) );
AND2X2 AND2X2_80 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_795_) );
OAI21X1 OAI21X1_234 ( .A(_794_), .B(_795_), .C(_60__3_), .Y(_796_) );
NAND2X1 NAND2X1_235 ( .A(_796_), .B(_800_), .Y(_58__3_) );
OAI21X1 OAI21X1_235 ( .A(_797_), .B(_794_), .C(_799_), .Y(_56_) );
INVX1 INVX1_156 ( .A(1'b0), .Y(_804_) );
OR2X2 OR2X2_81 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_805_) );
NAND2X1 NAND2X1_236 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_806_) );
NAND3X1 NAND3X1_81 ( .A(_804_), .B(_806_), .C(_805_), .Y(_807_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_801_) );
AND2X2 AND2X2_81 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_802_) );
OAI21X1 OAI21X1_236 ( .A(_801_), .B(_802_), .C(1'b0), .Y(_803_) );
NAND2X1 NAND2X1_237 ( .A(_803_), .B(_807_), .Y(_63__0_) );
OAI21X1 OAI21X1_237 ( .A(_804_), .B(_801_), .C(_806_), .Y(_65__1_) );
INVX1 INVX1_157 ( .A(_65__1_), .Y(_811_) );
OR2X2 OR2X2_82 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_812_) );
NAND2X1 NAND2X1_238 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_813_) );
NAND3X1 NAND3X1_82 ( .A(_811_), .B(_813_), .C(_812_), .Y(_814_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_808_) );
AND2X2 AND2X2_82 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_809_) );
OAI21X1 OAI21X1_238 ( .A(_808_), .B(_809_), .C(_65__1_), .Y(_810_) );
NAND2X1 NAND2X1_239 ( .A(_810_), .B(_814_), .Y(_63__1_) );
OAI21X1 OAI21X1_239 ( .A(_811_), .B(_808_), .C(_813_), .Y(_65__2_) );
INVX1 INVX1_158 ( .A(_65__2_), .Y(_818_) );
OR2X2 OR2X2_83 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_819_) );
NAND2X1 NAND2X1_240 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_820_) );
NAND3X1 NAND3X1_83 ( .A(_818_), .B(_820_), .C(_819_), .Y(_821_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_815_) );
AND2X2 AND2X2_83 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_816_) );
OAI21X1 OAI21X1_240 ( .A(_815_), .B(_816_), .C(_65__2_), .Y(_817_) );
NAND2X1 NAND2X1_241 ( .A(_817_), .B(_821_), .Y(_63__2_) );
OAI21X1 OAI21X1_241 ( .A(_818_), .B(_815_), .C(_820_), .Y(_65__3_) );
INVX1 INVX1_159 ( .A(_65__3_), .Y(_825_) );
OR2X2 OR2X2_84 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_826_) );
NAND2X1 NAND2X1_242 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_827_) );
NAND3X1 NAND3X1_84 ( .A(_825_), .B(_827_), .C(_826_), .Y(_828_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_822_) );
AND2X2 AND2X2_84 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_823_) );
OAI21X1 OAI21X1_242 ( .A(_822_), .B(_823_), .C(_65__3_), .Y(_824_) );
NAND2X1 NAND2X1_243 ( .A(_824_), .B(_828_), .Y(_63__3_) );
OAI21X1 OAI21X1_243 ( .A(_825_), .B(_822_), .C(_827_), .Y(_61_) );
INVX1 INVX1_160 ( .A(1'b1), .Y(_832_) );
OR2X2 OR2X2_85 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_833_) );
NAND2X1 NAND2X1_244 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_834_) );
NAND3X1 NAND3X1_85 ( .A(_832_), .B(_834_), .C(_833_), .Y(_835_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_829_) );
AND2X2 AND2X2_85 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_830_) );
OAI21X1 OAI21X1_244 ( .A(_829_), .B(_830_), .C(1'b1), .Y(_831_) );
NAND2X1 NAND2X1_245 ( .A(_831_), .B(_835_), .Y(_64__0_) );
OAI21X1 OAI21X1_245 ( .A(_832_), .B(_829_), .C(_834_), .Y(_66__1_) );
INVX1 INVX1_161 ( .A(_66__1_), .Y(_839_) );
OR2X2 OR2X2_86 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_840_) );
NAND2X1 NAND2X1_246 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_841_) );
NAND3X1 NAND3X1_86 ( .A(_839_), .B(_841_), .C(_840_), .Y(_842_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_836_) );
AND2X2 AND2X2_86 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_837_) );
OAI21X1 OAI21X1_246 ( .A(_836_), .B(_837_), .C(_66__1_), .Y(_838_) );
NAND2X1 NAND2X1_247 ( .A(_838_), .B(_842_), .Y(_64__1_) );
OAI21X1 OAI21X1_247 ( .A(_839_), .B(_836_), .C(_841_), .Y(_66__2_) );
INVX1 INVX1_162 ( .A(_66__2_), .Y(_846_) );
OR2X2 OR2X2_87 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_847_) );
NAND2X1 NAND2X1_248 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_848_) );
NAND3X1 NAND3X1_87 ( .A(_846_), .B(_848_), .C(_847_), .Y(_849_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_843_) );
AND2X2 AND2X2_87 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_844_) );
OAI21X1 OAI21X1_248 ( .A(_843_), .B(_844_), .C(_66__2_), .Y(_845_) );
NAND2X1 NAND2X1_249 ( .A(_845_), .B(_849_), .Y(_64__2_) );
OAI21X1 OAI21X1_249 ( .A(_846_), .B(_843_), .C(_848_), .Y(_66__3_) );
INVX1 INVX1_163 ( .A(_66__3_), .Y(_853_) );
OR2X2 OR2X2_88 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_854_) );
NAND2X1 NAND2X1_250 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_855_) );
NAND3X1 NAND3X1_88 ( .A(_853_), .B(_855_), .C(_854_), .Y(_856_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_850_) );
AND2X2 AND2X2_88 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_851_) );
OAI21X1 OAI21X1_250 ( .A(_850_), .B(_851_), .C(_66__3_), .Y(_852_) );
NAND2X1 NAND2X1_251 ( .A(_852_), .B(_856_), .Y(_64__3_) );
OAI21X1 OAI21X1_251 ( .A(_853_), .B(_850_), .C(_855_), .Y(_62_) );
INVX1 INVX1_164 ( .A(1'b0), .Y(_860_) );
OR2X2 OR2X2_89 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_861_) );
NAND2X1 NAND2X1_252 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_862_) );
NAND3X1 NAND3X1_89 ( .A(_860_), .B(_862_), .C(_861_), .Y(_863_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_857_) );
AND2X2 AND2X2_89 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_858_) );
OAI21X1 OAI21X1_252 ( .A(_857_), .B(_858_), .C(1'b0), .Y(_859_) );
NAND2X1 NAND2X1_253 ( .A(_859_), .B(_863_), .Y(_69__0_) );
OAI21X1 OAI21X1_253 ( .A(_860_), .B(_857_), .C(_862_), .Y(_71__1_) );
INVX1 INVX1_165 ( .A(_71__1_), .Y(_867_) );
OR2X2 OR2X2_90 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_868_) );
NAND2X1 NAND2X1_254 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_869_) );
NAND3X1 NAND3X1_90 ( .A(_867_), .B(_869_), .C(_868_), .Y(_870_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_864_) );
AND2X2 AND2X2_90 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_865_) );
OAI21X1 OAI21X1_254 ( .A(_864_), .B(_865_), .C(_71__1_), .Y(_866_) );
NAND2X1 NAND2X1_255 ( .A(_866_), .B(_870_), .Y(_69__1_) );
OAI21X1 OAI21X1_255 ( .A(_867_), .B(_864_), .C(_869_), .Y(_71__2_) );
INVX1 INVX1_166 ( .A(_71__2_), .Y(_874_) );
OR2X2 OR2X2_91 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_875_) );
NAND2X1 NAND2X1_256 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_876_) );
NAND3X1 NAND3X1_91 ( .A(_874_), .B(_876_), .C(_875_), .Y(_877_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_871_) );
AND2X2 AND2X2_91 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_872_) );
OAI21X1 OAI21X1_256 ( .A(_871_), .B(_872_), .C(_71__2_), .Y(_873_) );
NAND2X1 NAND2X1_257 ( .A(_873_), .B(_877_), .Y(_69__2_) );
OAI21X1 OAI21X1_257 ( .A(_874_), .B(_871_), .C(_876_), .Y(_71__3_) );
INVX1 INVX1_167 ( .A(_71__3_), .Y(_881_) );
OR2X2 OR2X2_92 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_882_) );
NAND2X1 NAND2X1_258 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_883_) );
NAND3X1 NAND3X1_92 ( .A(_881_), .B(_883_), .C(_882_), .Y(_884_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_878_) );
AND2X2 AND2X2_92 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_879_) );
OAI21X1 OAI21X1_258 ( .A(_878_), .B(_879_), .C(_71__3_), .Y(_880_) );
NAND2X1 NAND2X1_259 ( .A(_880_), .B(_884_), .Y(_69__3_) );
OAI21X1 OAI21X1_259 ( .A(_881_), .B(_878_), .C(_883_), .Y(_67_) );
INVX1 INVX1_168 ( .A(1'b1), .Y(_888_) );
OR2X2 OR2X2_93 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_889_) );
NAND2X1 NAND2X1_260 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_890_) );
NAND3X1 NAND3X1_93 ( .A(_888_), .B(_890_), .C(_889_), .Y(_891_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_885_) );
AND2X2 AND2X2_93 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_886_) );
OAI21X1 OAI21X1_260 ( .A(_885_), .B(_886_), .C(1'b1), .Y(_887_) );
NAND2X1 NAND2X1_261 ( .A(_887_), .B(_891_), .Y(_70__0_) );
OAI21X1 OAI21X1_261 ( .A(_888_), .B(_885_), .C(_890_), .Y(_72__1_) );
INVX1 INVX1_169 ( .A(_72__1_), .Y(_895_) );
OR2X2 OR2X2_94 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_896_) );
NAND2X1 NAND2X1_262 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_897_) );
NAND3X1 NAND3X1_94 ( .A(_895_), .B(_897_), .C(_896_), .Y(_898_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_892_) );
AND2X2 AND2X2_94 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_893_) );
OAI21X1 OAI21X1_262 ( .A(_892_), .B(_893_), .C(_72__1_), .Y(_894_) );
NAND2X1 NAND2X1_263 ( .A(_894_), .B(_898_), .Y(_70__1_) );
OAI21X1 OAI21X1_263 ( .A(_895_), .B(_892_), .C(_897_), .Y(_72__2_) );
INVX1 INVX1_170 ( .A(_72__2_), .Y(_902_) );
OR2X2 OR2X2_95 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_903_) );
NAND2X1 NAND2X1_264 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_904_) );
NAND3X1 NAND3X1_95 ( .A(_902_), .B(_904_), .C(_903_), .Y(_905_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_899_) );
AND2X2 AND2X2_95 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_900_) );
OAI21X1 OAI21X1_264 ( .A(_899_), .B(_900_), .C(_72__2_), .Y(_901_) );
NAND2X1 NAND2X1_265 ( .A(_901_), .B(_905_), .Y(_70__2_) );
OAI21X1 OAI21X1_265 ( .A(_902_), .B(_899_), .C(_904_), .Y(_72__3_) );
INVX1 INVX1_171 ( .A(_72__3_), .Y(_909_) );
OR2X2 OR2X2_96 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_910_) );
NAND2X1 NAND2X1_266 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_911_) );
NAND3X1 NAND3X1_96 ( .A(_909_), .B(_911_), .C(_910_), .Y(_912_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_906_) );
AND2X2 AND2X2_96 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_907_) );
OAI21X1 OAI21X1_266 ( .A(_906_), .B(_907_), .C(_72__3_), .Y(_908_) );
NAND2X1 NAND2X1_267 ( .A(_908_), .B(_912_), .Y(_70__3_) );
OAI21X1 OAI21X1_267 ( .A(_909_), .B(_906_), .C(_911_), .Y(_68_) );
INVX1 INVX1_172 ( .A(1'b0), .Y(_916_) );
OR2X2 OR2X2_97 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_917_) );
NAND2X1 NAND2X1_268 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_918_) );
NAND3X1 NAND3X1_97 ( .A(_916_), .B(_918_), .C(_917_), .Y(_919_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_913_) );
AND2X2 AND2X2_97 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_914_) );
OAI21X1 OAI21X1_268 ( .A(_913_), .B(_914_), .C(1'b0), .Y(_915_) );
NAND2X1 NAND2X1_269 ( .A(_915_), .B(_919_), .Y(_75__0_) );
OAI21X1 OAI21X1_269 ( .A(_916_), .B(_913_), .C(_918_), .Y(_77__1_) );
INVX1 INVX1_173 ( .A(_77__1_), .Y(_923_) );
OR2X2 OR2X2_98 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_924_) );
NAND2X1 NAND2X1_270 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_925_) );
NAND3X1 NAND3X1_98 ( .A(_923_), .B(_925_), .C(_924_), .Y(_926_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_920_) );
AND2X2 AND2X2_98 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_921_) );
OAI21X1 OAI21X1_270 ( .A(_920_), .B(_921_), .C(_77__1_), .Y(_922_) );
NAND2X1 NAND2X1_271 ( .A(_922_), .B(_926_), .Y(_75__1_) );
OAI21X1 OAI21X1_271 ( .A(_923_), .B(_920_), .C(_925_), .Y(_77__2_) );
INVX1 INVX1_174 ( .A(_77__2_), .Y(_930_) );
OR2X2 OR2X2_99 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_931_) );
NAND2X1 NAND2X1_272 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_932_) );
NAND3X1 NAND3X1_99 ( .A(_930_), .B(_932_), .C(_931_), .Y(_933_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_927_) );
AND2X2 AND2X2_99 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_928_) );
OAI21X1 OAI21X1_272 ( .A(_927_), .B(_928_), .C(_77__2_), .Y(_929_) );
NAND2X1 NAND2X1_273 ( .A(_929_), .B(_933_), .Y(_75__2_) );
OAI21X1 OAI21X1_273 ( .A(_930_), .B(_927_), .C(_932_), .Y(_77__3_) );
INVX1 INVX1_175 ( .A(_77__3_), .Y(_937_) );
OR2X2 OR2X2_100 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_938_) );
NAND2X1 NAND2X1_274 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_939_) );
NAND3X1 NAND3X1_100 ( .A(_937_), .B(_939_), .C(_938_), .Y(_940_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_934_) );
AND2X2 AND2X2_100 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_935_) );
OAI21X1 OAI21X1_274 ( .A(_934_), .B(_935_), .C(_77__3_), .Y(_936_) );
NAND2X1 NAND2X1_275 ( .A(_936_), .B(_940_), .Y(_75__3_) );
OAI21X1 OAI21X1_275 ( .A(_937_), .B(_934_), .C(_939_), .Y(_73_) );
INVX1 INVX1_176 ( .A(1'b1), .Y(_944_) );
OR2X2 OR2X2_101 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_945_) );
NAND2X1 NAND2X1_276 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_946_) );
NAND3X1 NAND3X1_101 ( .A(_944_), .B(_946_), .C(_945_), .Y(_947_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_941_) );
AND2X2 AND2X2_101 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_942_) );
OAI21X1 OAI21X1_276 ( .A(_941_), .B(_942_), .C(1'b1), .Y(_943_) );
NAND2X1 NAND2X1_277 ( .A(_943_), .B(_947_), .Y(_76__0_) );
OAI21X1 OAI21X1_277 ( .A(_944_), .B(_941_), .C(_946_), .Y(_78__1_) );
INVX1 INVX1_177 ( .A(_78__1_), .Y(_951_) );
OR2X2 OR2X2_102 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_952_) );
NAND2X1 NAND2X1_278 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_953_) );
NAND3X1 NAND3X1_102 ( .A(_951_), .B(_953_), .C(_952_), .Y(_954_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_948_) );
AND2X2 AND2X2_102 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_949_) );
OAI21X1 OAI21X1_278 ( .A(_948_), .B(_949_), .C(_78__1_), .Y(_950_) );
NAND2X1 NAND2X1_279 ( .A(_950_), .B(_954_), .Y(_76__1_) );
OAI21X1 OAI21X1_279 ( .A(_951_), .B(_948_), .C(_953_), .Y(_78__2_) );
INVX1 INVX1_178 ( .A(_78__2_), .Y(_958_) );
OR2X2 OR2X2_103 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_959_) );
NAND2X1 NAND2X1_280 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_960_) );
NAND3X1 NAND3X1_103 ( .A(_958_), .B(_960_), .C(_959_), .Y(_961_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_955_) );
AND2X2 AND2X2_103 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_956_) );
OAI21X1 OAI21X1_280 ( .A(_955_), .B(_956_), .C(_78__2_), .Y(_957_) );
NAND2X1 NAND2X1_281 ( .A(_957_), .B(_961_), .Y(_76__2_) );
OAI21X1 OAI21X1_281 ( .A(_958_), .B(_955_), .C(_960_), .Y(_78__3_) );
INVX1 INVX1_179 ( .A(_78__3_), .Y(_965_) );
OR2X2 OR2X2_104 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_966_) );
NAND2X1 NAND2X1_282 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_967_) );
NAND3X1 NAND3X1_104 ( .A(_965_), .B(_967_), .C(_966_), .Y(_968_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_962_) );
AND2X2 AND2X2_104 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_963_) );
OAI21X1 OAI21X1_282 ( .A(_962_), .B(_963_), .C(_78__3_), .Y(_964_) );
NAND2X1 NAND2X1_283 ( .A(_964_), .B(_968_), .Y(_76__3_) );
OAI21X1 OAI21X1_283 ( .A(_965_), .B(_962_), .C(_967_), .Y(_74_) );
INVX1 INVX1_180 ( .A(1'b0), .Y(_972_) );
OR2X2 OR2X2_105 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_973_) );
NAND2X1 NAND2X1_284 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_974_) );
NAND3X1 NAND3X1_105 ( .A(_972_), .B(_974_), .C(_973_), .Y(_975_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_969_) );
AND2X2 AND2X2_105 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_970_) );
OAI21X1 OAI21X1_284 ( .A(_969_), .B(_970_), .C(1'b0), .Y(_971_) );
NAND2X1 NAND2X1_285 ( .A(_971_), .B(_975_), .Y(_81__0_) );
OAI21X1 OAI21X1_285 ( .A(_972_), .B(_969_), .C(_974_), .Y(_83__1_) );
INVX1 INVX1_181 ( .A(_83__1_), .Y(_979_) );
OR2X2 OR2X2_106 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_980_) );
NAND2X1 NAND2X1_286 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_981_) );
NAND3X1 NAND3X1_106 ( .A(_979_), .B(_981_), .C(_980_), .Y(_982_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_976_) );
AND2X2 AND2X2_106 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_977_) );
OAI21X1 OAI21X1_286 ( .A(_976_), .B(_977_), .C(_83__1_), .Y(_978_) );
NAND2X1 NAND2X1_287 ( .A(_978_), .B(_982_), .Y(_81__1_) );
OAI21X1 OAI21X1_287 ( .A(_979_), .B(_976_), .C(_981_), .Y(_83__2_) );
INVX1 INVX1_182 ( .A(_83__2_), .Y(_986_) );
OR2X2 OR2X2_107 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_987_) );
NAND2X1 NAND2X1_288 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_988_) );
NAND3X1 NAND3X1_107 ( .A(_986_), .B(_988_), .C(_987_), .Y(_989_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_983_) );
AND2X2 AND2X2_107 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_984_) );
OAI21X1 OAI21X1_288 ( .A(_983_), .B(_984_), .C(_83__2_), .Y(_985_) );
NAND2X1 NAND2X1_289 ( .A(_985_), .B(_989_), .Y(_81__2_) );
OAI21X1 OAI21X1_289 ( .A(_986_), .B(_983_), .C(_988_), .Y(_83__3_) );
INVX1 INVX1_183 ( .A(_83__3_), .Y(_993_) );
OR2X2 OR2X2_108 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_994_) );
NAND2X1 NAND2X1_290 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_995_) );
NAND3X1 NAND3X1_108 ( .A(_993_), .B(_995_), .C(_994_), .Y(_996_) );
NOR2X1 NOR2X1_108 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_990_) );
AND2X2 AND2X2_108 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_991_) );
OAI21X1 OAI21X1_290 ( .A(_990_), .B(_991_), .C(_83__3_), .Y(_992_) );
NAND2X1 NAND2X1_291 ( .A(_992_), .B(_996_), .Y(_81__3_) );
OAI21X1 OAI21X1_291 ( .A(_993_), .B(_990_), .C(_995_), .Y(_79_) );
INVX1 INVX1_184 ( .A(1'b1), .Y(_1000_) );
OR2X2 OR2X2_109 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_1001_) );
NAND2X1 NAND2X1_292 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_1002_) );
NAND3X1 NAND3X1_109 ( .A(_1000_), .B(_1002_), .C(_1001_), .Y(_1003_) );
NOR2X1 NOR2X1_109 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_997_) );
AND2X2 AND2X2_109 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_998_) );
OAI21X1 OAI21X1_292 ( .A(_997_), .B(_998_), .C(1'b1), .Y(_999_) );
NAND2X1 NAND2X1_293 ( .A(_999_), .B(_1003_), .Y(_82__0_) );
OAI21X1 OAI21X1_293 ( .A(_1000_), .B(_997_), .C(_1002_), .Y(_84__1_) );
INVX1 INVX1_185 ( .A(_84__1_), .Y(_1007_) );
OR2X2 OR2X2_110 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_1008_) );
NAND2X1 NAND2X1_294 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_1009_) );
NAND3X1 NAND3X1_110 ( .A(_1007_), .B(_1009_), .C(_1008_), .Y(_1010_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_1004_) );
AND2X2 AND2X2_110 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_1005_) );
OAI21X1 OAI21X1_294 ( .A(_1004_), .B(_1005_), .C(_84__1_), .Y(_1006_) );
NAND2X1 NAND2X1_295 ( .A(_1006_), .B(_1010_), .Y(_82__1_) );
OAI21X1 OAI21X1_295 ( .A(_1007_), .B(_1004_), .C(_1009_), .Y(_84__2_) );
INVX1 INVX1_186 ( .A(_84__2_), .Y(_1014_) );
OR2X2 OR2X2_111 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_1015_) );
NAND2X1 NAND2X1_296 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_1016_) );
NAND3X1 NAND3X1_111 ( .A(_1014_), .B(_1016_), .C(_1015_), .Y(_1017_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_1011_) );
AND2X2 AND2X2_111 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_1012_) );
OAI21X1 OAI21X1_296 ( .A(_1011_), .B(_1012_), .C(_84__2_), .Y(_1013_) );
NAND2X1 NAND2X1_297 ( .A(_1013_), .B(_1017_), .Y(_82__2_) );
OAI21X1 OAI21X1_297 ( .A(_1014_), .B(_1011_), .C(_1016_), .Y(_84__3_) );
INVX1 INVX1_187 ( .A(_84__3_), .Y(_1021_) );
OR2X2 OR2X2_112 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_1022_) );
NAND2X1 NAND2X1_298 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_1023_) );
NAND3X1 NAND3X1_112 ( .A(_1021_), .B(_1023_), .C(_1022_), .Y(_1024_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_1018_) );
AND2X2 AND2X2_112 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_1019_) );
OAI21X1 OAI21X1_298 ( .A(_1018_), .B(_1019_), .C(_84__3_), .Y(_1020_) );
NAND2X1 NAND2X1_299 ( .A(_1020_), .B(_1024_), .Y(_82__3_) );
OAI21X1 OAI21X1_299 ( .A(_1021_), .B(_1018_), .C(_1023_), .Y(_80_) );
INVX1 INVX1_188 ( .A(1'b0), .Y(_1028_) );
OR2X2 OR2X2_113 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_1029_) );
NAND2X1 NAND2X1_300 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_1030_) );
NAND3X1 NAND3X1_113 ( .A(_1028_), .B(_1030_), .C(_1029_), .Y(_1031_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_1025_) );
AND2X2 AND2X2_113 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_1026_) );
OAI21X1 OAI21X1_300 ( .A(_1025_), .B(_1026_), .C(1'b0), .Y(_1027_) );
NAND2X1 NAND2X1_301 ( .A(_1027_), .B(_1031_), .Y(_87__0_) );
OAI21X1 OAI21X1_301 ( .A(_1028_), .B(_1025_), .C(_1030_), .Y(_89__1_) );
INVX1 INVX1_189 ( .A(_89__1_), .Y(_1035_) );
OR2X2 OR2X2_114 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1036_) );
NAND2X1 NAND2X1_302 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1037_) );
NAND3X1 NAND3X1_114 ( .A(_1035_), .B(_1037_), .C(_1036_), .Y(_1038_) );
NOR2X1 NOR2X1_114 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1032_) );
AND2X2 AND2X2_114 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1033_) );
OAI21X1 OAI21X1_302 ( .A(_1032_), .B(_1033_), .C(_89__1_), .Y(_1034_) );
NAND2X1 NAND2X1_303 ( .A(_1034_), .B(_1038_), .Y(_87__1_) );
OAI21X1 OAI21X1_303 ( .A(_1035_), .B(_1032_), .C(_1037_), .Y(_89__2_) );
INVX1 INVX1_190 ( .A(_89__2_), .Y(_1042_) );
OR2X2 OR2X2_115 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_1043_) );
NAND2X1 NAND2X1_304 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_1044_) );
NAND3X1 NAND3X1_115 ( .A(_1042_), .B(_1044_), .C(_1043_), .Y(_1045_) );
NOR2X1 NOR2X1_115 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_1039_) );
AND2X2 AND2X2_115 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_1040_) );
OAI21X1 OAI21X1_304 ( .A(_1039_), .B(_1040_), .C(_89__2_), .Y(_1041_) );
NAND2X1 NAND2X1_305 ( .A(_1041_), .B(_1045_), .Y(_87__2_) );
OAI21X1 OAI21X1_305 ( .A(_1042_), .B(_1039_), .C(_1044_), .Y(_89__3_) );
INVX1 INVX1_191 ( .A(_89__3_), .Y(_1049_) );
OR2X2 OR2X2_116 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1050_) );
NAND2X1 NAND2X1_306 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1051_) );
NAND3X1 NAND3X1_116 ( .A(_1049_), .B(_1051_), .C(_1050_), .Y(_1052_) );
NOR2X1 NOR2X1_116 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1046_) );
AND2X2 AND2X2_116 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1047_) );
OAI21X1 OAI21X1_306 ( .A(_1046_), .B(_1047_), .C(_89__3_), .Y(_1048_) );
NAND2X1 NAND2X1_307 ( .A(_1048_), .B(_1052_), .Y(_87__3_) );
OAI21X1 OAI21X1_307 ( .A(_1049_), .B(_1046_), .C(_1051_), .Y(_85_) );
INVX1 INVX1_192 ( .A(1'b1), .Y(_1056_) );
OR2X2 OR2X2_117 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_1057_) );
NAND2X1 NAND2X1_308 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_1058_) );
NAND3X1 NAND3X1_117 ( .A(_1056_), .B(_1058_), .C(_1057_), .Y(_1059_) );
NOR2X1 NOR2X1_117 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_1053_) );
AND2X2 AND2X2_117 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_1054_) );
OAI21X1 OAI21X1_308 ( .A(_1053_), .B(_1054_), .C(1'b1), .Y(_1055_) );
NAND2X1 NAND2X1_309 ( .A(_1055_), .B(_1059_), .Y(_88__0_) );
OAI21X1 OAI21X1_309 ( .A(_1056_), .B(_1053_), .C(_1058_), .Y(_90__1_) );
INVX1 INVX1_193 ( .A(_90__1_), .Y(_1063_) );
OR2X2 OR2X2_118 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1064_) );
NAND2X1 NAND2X1_310 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1065_) );
NAND3X1 NAND3X1_118 ( .A(_1063_), .B(_1065_), .C(_1064_), .Y(_1066_) );
NOR2X1 NOR2X1_118 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1060_) );
AND2X2 AND2X2_118 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1061_) );
OAI21X1 OAI21X1_310 ( .A(_1060_), .B(_1061_), .C(_90__1_), .Y(_1062_) );
NAND2X1 NAND2X1_311 ( .A(_1062_), .B(_1066_), .Y(_88__1_) );
OAI21X1 OAI21X1_311 ( .A(_1063_), .B(_1060_), .C(_1065_), .Y(_90__2_) );
INVX1 INVX1_194 ( .A(_90__2_), .Y(_1070_) );
OR2X2 OR2X2_119 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_1071_) );
NAND2X1 NAND2X1_312 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_1072_) );
NAND3X1 NAND3X1_119 ( .A(_1070_), .B(_1072_), .C(_1071_), .Y(_1073_) );
NOR2X1 NOR2X1_119 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_1067_) );
AND2X2 AND2X2_119 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_1068_) );
OAI21X1 OAI21X1_312 ( .A(_1067_), .B(_1068_), .C(_90__2_), .Y(_1069_) );
NAND2X1 NAND2X1_313 ( .A(_1069_), .B(_1073_), .Y(_88__2_) );
OAI21X1 OAI21X1_313 ( .A(_1070_), .B(_1067_), .C(_1072_), .Y(_90__3_) );
INVX1 INVX1_195 ( .A(_90__3_), .Y(_1077_) );
OR2X2 OR2X2_120 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1078_) );
NAND2X1 NAND2X1_314 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1079_) );
NAND3X1 NAND3X1_120 ( .A(_1077_), .B(_1079_), .C(_1078_), .Y(_1080_) );
NOR2X1 NOR2X1_120 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1074_) );
AND2X2 AND2X2_120 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1075_) );
OAI21X1 OAI21X1_314 ( .A(_1074_), .B(_1075_), .C(_90__3_), .Y(_1076_) );
NAND2X1 NAND2X1_315 ( .A(_1076_), .B(_1080_), .Y(_88__3_) );
OAI21X1 OAI21X1_315 ( .A(_1077_), .B(_1074_), .C(_1079_), .Y(_86_) );
INVX1 INVX1_196 ( .A(1'b0), .Y(_1084_) );
OR2X2 OR2X2_121 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1085_) );
NAND2X1 NAND2X1_316 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1086_) );
NAND3X1 NAND3X1_121 ( .A(_1084_), .B(_1086_), .C(_1085_), .Y(_1087_) );
NOR2X1 NOR2X1_121 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1081_) );
AND2X2 AND2X2_121 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1082_) );
OAI21X1 OAI21X1_316 ( .A(_1081_), .B(_1082_), .C(1'b0), .Y(_1083_) );
NAND2X1 NAND2X1_317 ( .A(_1083_), .B(_1087_), .Y(rca_inst_w_SUM) );
BUFX2 BUFX2_63 ( .A(rca_inst_w_SUM), .Y(_0__0_) );
BUFX2 BUFX2_64 ( .A(1'b0), .Y(_5__0_) );
BUFX2 BUFX2_65 ( .A(_1_), .Y(_5__4_) );
BUFX2 BUFX2_66 ( .A(1'b1), .Y(_6__0_) );
BUFX2 BUFX2_67 ( .A(_2_), .Y(_6__4_) );
BUFX2 BUFX2_68 ( .A(1'b0), .Y(_11__0_) );
BUFX2 BUFX2_69 ( .A(_7_), .Y(_11__4_) );
BUFX2 BUFX2_70 ( .A(1'b1), .Y(_12__0_) );
BUFX2 BUFX2_71 ( .A(_8_), .Y(_12__4_) );
BUFX2 BUFX2_72 ( .A(1'b0), .Y(_17__0_) );
BUFX2 BUFX2_73 ( .A(_13_), .Y(_17__4_) );
BUFX2 BUFX2_74 ( .A(1'b1), .Y(_18__0_) );
BUFX2 BUFX2_75 ( .A(_14_), .Y(_18__4_) );
BUFX2 BUFX2_76 ( .A(1'b0), .Y(_23__0_) );
BUFX2 BUFX2_77 ( .A(_19_), .Y(_23__4_) );
BUFX2 BUFX2_78 ( .A(1'b1), .Y(_24__0_) );
BUFX2 BUFX2_79 ( .A(_20_), .Y(_24__4_) );
BUFX2 BUFX2_80 ( .A(1'b0), .Y(_29__0_) );
BUFX2 BUFX2_81 ( .A(_25_), .Y(_29__4_) );
BUFX2 BUFX2_82 ( .A(1'b1), .Y(_30__0_) );
BUFX2 BUFX2_83 ( .A(_26_), .Y(_30__4_) );
BUFX2 BUFX2_84 ( .A(1'b0), .Y(_35__0_) );
BUFX2 BUFX2_85 ( .A(_31_), .Y(_35__4_) );
BUFX2 BUFX2_86 ( .A(1'b1), .Y(_36__0_) );
BUFX2 BUFX2_87 ( .A(_32_), .Y(_36__4_) );
BUFX2 BUFX2_88 ( .A(1'b0), .Y(_41__0_) );
BUFX2 BUFX2_89 ( .A(_37_), .Y(_41__4_) );
BUFX2 BUFX2_90 ( .A(1'b1), .Y(_42__0_) );
BUFX2 BUFX2_91 ( .A(_38_), .Y(_42__4_) );
BUFX2 BUFX2_92 ( .A(1'b0), .Y(_47__0_) );
BUFX2 BUFX2_93 ( .A(_43_), .Y(_47__4_) );
BUFX2 BUFX2_94 ( .A(1'b1), .Y(_48__0_) );
BUFX2 BUFX2_95 ( .A(_44_), .Y(_48__4_) );
BUFX2 BUFX2_96 ( .A(1'b0), .Y(_53__0_) );
BUFX2 BUFX2_97 ( .A(_49_), .Y(_53__4_) );
BUFX2 BUFX2_98 ( .A(1'b1), .Y(_54__0_) );
BUFX2 BUFX2_99 ( .A(_50_), .Y(_54__4_) );
BUFX2 BUFX2_100 ( .A(1'b0), .Y(_59__0_) );
BUFX2 BUFX2_101 ( .A(_55_), .Y(_59__4_) );
BUFX2 BUFX2_102 ( .A(1'b1), .Y(_60__0_) );
BUFX2 BUFX2_103 ( .A(_56_), .Y(_60__4_) );
BUFX2 BUFX2_104 ( .A(1'b0), .Y(_65__0_) );
BUFX2 BUFX2_105 ( .A(_61_), .Y(_65__4_) );
BUFX2 BUFX2_106 ( .A(1'b1), .Y(_66__0_) );
BUFX2 BUFX2_107 ( .A(_62_), .Y(_66__4_) );
BUFX2 BUFX2_108 ( .A(1'b0), .Y(_71__0_) );
BUFX2 BUFX2_109 ( .A(_67_), .Y(_71__4_) );
BUFX2 BUFX2_110 ( .A(1'b1), .Y(_72__0_) );
BUFX2 BUFX2_111 ( .A(_68_), .Y(_72__4_) );
BUFX2 BUFX2_112 ( .A(1'b0), .Y(_77__0_) );
BUFX2 BUFX2_113 ( .A(_73_), .Y(_77__4_) );
BUFX2 BUFX2_114 ( .A(1'b1), .Y(_78__0_) );
BUFX2 BUFX2_115 ( .A(_74_), .Y(_78__4_) );
BUFX2 BUFX2_116 ( .A(1'b0), .Y(_83__0_) );
BUFX2 BUFX2_117 ( .A(_79_), .Y(_83__4_) );
BUFX2 BUFX2_118 ( .A(1'b1), .Y(_84__0_) );
BUFX2 BUFX2_119 ( .A(_80_), .Y(_84__4_) );
BUFX2 BUFX2_120 ( .A(1'b0), .Y(_89__0_) );
BUFX2 BUFX2_121 ( .A(_85_), .Y(_89__4_) );
BUFX2 BUFX2_122 ( .A(1'b1), .Y(_90__0_) );
BUFX2 BUFX2_123 ( .A(_86_), .Y(_90__4_) );
BUFX2 BUFX2_124 ( .A(1'b0), .Y(w_cout_0_) );
endmodule
