module csa_64bit ( gnd, vdd, i_add_term1, i_add_term2, sum, cout);

input gnd, vdd;
output cout;
input [63:0] i_add_term1;
input [63:0] i_add_term2;
output [63:0] sum;

BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(w_cout_15_), .Y(cout) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_0__54_), .Y(sum[54]) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_0__55_), .Y(sum[55]) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_0__56_), .Y(sum[56]) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_0__57_), .Y(sum[57]) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(_0__58_), .Y(sum[58]) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(_0__59_), .Y(sum[59]) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(_0__60_), .Y(sum[60]) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(_0__61_), .Y(sum[61]) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(_0__62_), .Y(sum[62]) );
BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(_0__63_), .Y(sum[63]) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_91_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(rca_inst_cout), .Y(_92_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_91_), .C(_92_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_3__0_), .Y(_93_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_4__0_), .B(rca_inst_cout), .Y(_94_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_93_), .C(_94_), .Y(_0__4_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_3__1_), .Y(_95_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_4__1_), .Y(_96_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_95_), .C(_96_), .Y(_0__5_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_3__2_), .Y(_97_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_4__2_), .Y(_98_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_97_), .C(_98_), .Y(_0__6_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_3__3_), .Y(_99_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_4__3_), .Y(_100_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_99_), .C(_100_), .Y(_0__7_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_104_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_105_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_106_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_106_), .C(_105_), .Y(_107_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_101_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_102_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_102_), .C(gnd), .Y(_103_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_107_), .Y(_3__0_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_101_), .C(_106_), .Y(_5__1_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_5__3_), .Y(_111_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_112_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_113_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_113_), .C(_112_), .Y(_114_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_108_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_109_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_109_), .C(_5__3_), .Y(_110_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_114_), .Y(_3__3_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_108_), .C(_113_), .Y(_1_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_5__1_), .Y(_118_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_119_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_120_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_120_), .C(_119_), .Y(_121_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_115_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_116_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_116_), .C(_5__1_), .Y(_117_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_121_), .Y(_3__1_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_115_), .C(_120_), .Y(_5__2_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_5__2_), .Y(_125_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_126_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_127_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_127_), .C(_126_), .Y(_128_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_122_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_123_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_123_), .C(_5__2_), .Y(_124_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_128_), .Y(_3__2_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_122_), .C(_127_), .Y(_5__3_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_132_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_133_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_134_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_134_), .C(_133_), .Y(_135_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_129_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_130_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_129_), .B(_130_), .C(vdd), .Y(_131_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_135_), .Y(_4__0_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_129_), .C(_134_), .Y(_6__1_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_6__3_), .Y(_139_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_140_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_141_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_141_), .C(_140_), .Y(_142_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_136_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_137_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_137_), .C(_6__3_), .Y(_138_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_142_), .Y(_4__3_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_136_), .C(_141_), .Y(_2_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_6__1_), .Y(_146_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_147_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_148_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_148_), .C(_147_), .Y(_149_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_143_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_144_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_144_), .C(_6__1_), .Y(_145_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_149_), .Y(_4__1_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_143_), .C(_148_), .Y(_6__2_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_6__2_), .Y(_153_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_154_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_155_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_155_), .C(_154_), .Y(_156_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_150_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_151_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_151_), .C(_6__2_), .Y(_152_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_156_), .Y(_4__2_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_150_), .C(_155_), .Y(_6__3_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_157_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(w_cout_1_), .Y(_158_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_157_), .C(_158_), .Y(w_cout_2_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_9__0_), .Y(_159_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_10__0_), .B(w_cout_1_), .Y(_160_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_159_), .C(_160_), .Y(_0__8_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_9__1_), .Y(_161_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_10__1_), .Y(_162_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_161_), .C(_162_), .Y(_0__9_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_9__2_), .Y(_163_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_10__2_), .Y(_164_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_163_), .C(_164_), .Y(_0__10_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_9__3_), .Y(_165_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_10__3_), .Y(_166_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_165_), .C(_166_), .Y(_0__11_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_170_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_171_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_172_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_172_), .C(_171_), .Y(_173_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_167_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_168_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_168_), .C(gnd), .Y(_169_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_173_), .Y(_9__0_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_167_), .C(_172_), .Y(_11__1_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_11__3_), .Y(_177_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_178_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_179_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_179_), .C(_178_), .Y(_180_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_174_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_175_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_175_), .C(_11__3_), .Y(_176_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_180_), .Y(_9__3_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_174_), .C(_179_), .Y(_7_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_11__1_), .Y(_184_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_185_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_186_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_186_), .C(_185_), .Y(_187_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_181_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_182_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_182_), .C(_11__1_), .Y(_183_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_187_), .Y(_9__1_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_181_), .C(_186_), .Y(_11__2_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_11__2_), .Y(_191_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_192_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_193_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_193_), .C(_192_), .Y(_194_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_188_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_189_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_189_), .C(_11__2_), .Y(_190_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_194_), .Y(_9__2_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_188_), .C(_193_), .Y(_11__3_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_198_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_199_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_200_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_200_), .C(_199_), .Y(_201_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_195_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_196_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_196_), .C(vdd), .Y(_197_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_201_), .Y(_10__0_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_195_), .C(_200_), .Y(_12__1_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_12__3_), .Y(_205_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_206_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_207_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_207_), .C(_206_), .Y(_208_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_202_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_203_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_203_), .C(_12__3_), .Y(_204_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_208_), .Y(_10__3_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_202_), .C(_207_), .Y(_8_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_12__1_), .Y(_212_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_213_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_214_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_214_), .C(_213_), .Y(_215_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_209_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_210_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_210_), .C(_12__1_), .Y(_211_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_215_), .Y(_10__1_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_209_), .C(_214_), .Y(_12__2_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_12__2_), .Y(_219_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_220_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_221_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_221_), .C(_220_), .Y(_222_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_216_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_217_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_217_), .C(_12__2_), .Y(_218_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(_222_), .Y(_10__2_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_216_), .C(_221_), .Y(_12__3_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_223_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(w_cout_2_), .Y(_224_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_223_), .C(_224_), .Y(w_cout_3_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_15__0_), .Y(_225_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_16__0_), .B(w_cout_2_), .Y(_226_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_225_), .C(_226_), .Y(_0__12_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_15__1_), .Y(_227_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_16__1_), .Y(_228_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_227_), .C(_228_), .Y(_0__13_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_15__2_), .Y(_229_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_16__2_), .Y(_230_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_229_), .C(_230_), .Y(_0__14_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_15__3_), .Y(_231_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_16__3_), .Y(_232_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_231_), .C(_232_), .Y(_0__15_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_236_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_237_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_238_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_238_), .C(_237_), .Y(_239_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_233_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_234_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_234_), .C(gnd), .Y(_235_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_239_), .Y(_15__0_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_233_), .C(_238_), .Y(_17__1_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_17__3_), .Y(_243_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_244_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_245_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_245_), .C(_244_), .Y(_246_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_240_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_241_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_241_), .C(_17__3_), .Y(_242_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_246_), .Y(_15__3_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_240_), .C(_245_), .Y(_13_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_17__1_), .Y(_250_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_251_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_252_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_252_), .C(_251_), .Y(_253_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_247_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_248_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_248_), .C(_17__1_), .Y(_249_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_253_), .Y(_15__1_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_247_), .C(_252_), .Y(_17__2_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_17__2_), .Y(_257_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_258_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_259_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_259_), .C(_258_), .Y(_260_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_254_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_255_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_255_), .C(_17__2_), .Y(_256_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_260_), .Y(_15__2_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_254_), .C(_259_), .Y(_17__3_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_264_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_265_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_266_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_266_), .C(_265_), .Y(_267_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_261_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_262_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_262_), .C(vdd), .Y(_263_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_267_), .Y(_16__0_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_261_), .C(_266_), .Y(_18__1_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_18__3_), .Y(_271_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_272_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_273_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_273_), .C(_272_), .Y(_274_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_268_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_269_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_269_), .C(_18__3_), .Y(_270_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_274_), .Y(_16__3_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_268_), .C(_273_), .Y(_14_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_18__1_), .Y(_278_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_279_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_280_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_280_), .C(_279_), .Y(_281_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_275_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_276_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_276_), .C(_18__1_), .Y(_277_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_281_), .Y(_16__1_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_275_), .C(_280_), .Y(_18__2_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_18__2_), .Y(_285_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_286_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_287_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_287_), .C(_286_), .Y(_288_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_282_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_283_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_283_), .C(_18__2_), .Y(_284_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_288_), .Y(_16__2_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_282_), .C(_287_), .Y(_18__3_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_289_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(w_cout_3_), .Y(_290_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_289_), .C(_290_), .Y(w_cout_4_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_21__0_), .Y(_291_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_22__0_), .B(w_cout_3_), .Y(_292_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_291_), .C(_292_), .Y(_0__16_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_21__1_), .Y(_293_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_22__1_), .Y(_294_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_293_), .C(_294_), .Y(_0__17_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_21__2_), .Y(_295_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_22__2_), .Y(_296_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_295_), .C(_296_), .Y(_0__18_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_21__3_), .Y(_297_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_22__3_), .Y(_298_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_297_), .C(_298_), .Y(_0__19_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_302_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_303_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_304_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_304_), .C(_303_), .Y(_305_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_299_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_300_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_300_), .C(gnd), .Y(_301_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_305_), .Y(_21__0_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_299_), .C(_304_), .Y(_23__1_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_23__3_), .Y(_309_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_310_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_311_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_311_), .C(_310_), .Y(_312_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_306_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_307_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_307_), .C(_23__3_), .Y(_308_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_312_), .Y(_21__3_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_306_), .C(_311_), .Y(_19_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_23__1_), .Y(_316_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_317_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_318_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_316_), .B(_318_), .C(_317_), .Y(_319_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_313_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_314_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_314_), .C(_23__1_), .Y(_315_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_319_), .Y(_21__1_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_316_), .B(_313_), .C(_318_), .Y(_23__2_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_23__2_), .Y(_323_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_324_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_325_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_325_), .C(_324_), .Y(_326_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_320_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_321_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_321_), .C(_23__2_), .Y(_322_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_326_), .Y(_21__2_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_320_), .C(_325_), .Y(_23__3_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_330_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_331_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_332_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_332_), .C(_331_), .Y(_333_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_327_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_328_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_328_), .C(vdd), .Y(_329_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_333_), .Y(_22__0_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_327_), .C(_332_), .Y(_24__1_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_24__3_), .Y(_337_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_338_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_339_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_339_), .C(_338_), .Y(_340_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_334_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_335_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_335_), .C(_24__3_), .Y(_336_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_340_), .Y(_22__3_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_334_), .C(_339_), .Y(_20_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_24__1_), .Y(_344_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_345_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_346_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_346_), .C(_345_), .Y(_347_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_341_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_342_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_342_), .C(_24__1_), .Y(_343_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_347_), .Y(_22__1_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_341_), .C(_346_), .Y(_24__2_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_24__2_), .Y(_351_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_352_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_353_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_353_), .C(_352_), .Y(_354_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_348_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_349_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_349_), .C(_24__2_), .Y(_350_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_354_), .Y(_22__2_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_348_), .C(_353_), .Y(_24__3_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(_355_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(w_cout_4_), .Y(_356_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_355_), .C(_356_), .Y(w_cout_5_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_27__0_), .Y(_357_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_28__0_), .B(w_cout_4_), .Y(_358_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_357_), .C(_358_), .Y(_0__20_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_27__1_), .Y(_359_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_28__1_), .Y(_360_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_359_), .C(_360_), .Y(_0__21_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_27__2_), .Y(_361_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_28__2_), .Y(_362_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_361_), .C(_362_), .Y(_0__22_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_27__3_), .Y(_363_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_28__3_), .Y(_364_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_363_), .C(_364_), .Y(_0__23_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_368_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_369_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_370_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_370_), .C(_369_), .Y(_371_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_365_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_366_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_365_), .B(_366_), .C(gnd), .Y(_367_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_371_), .Y(_27__0_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_365_), .C(_370_), .Y(_29__1_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_29__3_), .Y(_375_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_376_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_377_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_377_), .C(_376_), .Y(_378_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_372_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_373_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_373_), .C(_29__3_), .Y(_374_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_378_), .Y(_27__3_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_372_), .C(_377_), .Y(_25_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_29__1_), .Y(_382_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_383_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_384_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_382_), .B(_384_), .C(_383_), .Y(_385_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_379_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_380_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_380_), .C(_29__1_), .Y(_381_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_385_), .Y(_27__1_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_382_), .B(_379_), .C(_384_), .Y(_29__2_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_29__2_), .Y(_389_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_390_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_391_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_391_), .C(_390_), .Y(_392_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_386_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_387_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_387_), .C(_29__2_), .Y(_388_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(_392_), .Y(_27__2_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_386_), .C(_391_), .Y(_29__3_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_396_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_397_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_398_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_398_), .C(_397_), .Y(_399_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_393_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_394_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_394_), .C(vdd), .Y(_395_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_399_), .Y(_28__0_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_393_), .C(_398_), .Y(_30__1_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_30__3_), .Y(_403_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_404_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_405_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_405_), .C(_404_), .Y(_406_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_400_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_401_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_400_), .B(_401_), .C(_30__3_), .Y(_402_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_406_), .Y(_28__3_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_400_), .C(_405_), .Y(_26_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_30__1_), .Y(_410_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_411_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_412_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(_412_), .C(_411_), .Y(_413_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_407_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_408_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_408_), .C(_30__1_), .Y(_409_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_413_), .Y(_28__1_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(_407_), .C(_412_), .Y(_30__2_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_30__2_), .Y(_417_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_418_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_419_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_419_), .C(_418_), .Y(_420_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_414_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_415_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_414_), .B(_415_), .C(_30__2_), .Y(_416_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_420_), .Y(_28__2_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_414_), .C(_419_), .Y(_30__3_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_31_), .Y(_421_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(w_cout_5_), .Y(_422_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_421_), .C(_422_), .Y(w_cout_6_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_33__0_), .Y(_423_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_34__0_), .B(w_cout_5_), .Y(_424_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_423_), .C(_424_), .Y(_0__24_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_33__1_), .Y(_425_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_34__1_), .Y(_426_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_425_), .C(_426_), .Y(_0__25_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_33__2_), .Y(_427_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_34__2_), .Y(_428_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_427_), .C(_428_), .Y(_0__26_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_33__3_), .Y(_429_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_34__3_), .Y(_430_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_429_), .C(_430_), .Y(_0__27_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_434_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_435_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_436_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_436_), .C(_435_), .Y(_437_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_431_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_432_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_432_), .C(gnd), .Y(_433_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_437_), .Y(_33__0_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_431_), .C(_436_), .Y(_35__1_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_35__3_), .Y(_441_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_442_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_443_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_443_), .C(_442_), .Y(_444_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_438_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_439_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_439_), .C(_35__3_), .Y(_440_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_444_), .Y(_33__3_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_438_), .C(_443_), .Y(_31_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(_35__1_), .Y(_448_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_449_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_450_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_448_), .B(_450_), .C(_449_), .Y(_451_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_445_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_446_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_445_), .B(_446_), .C(_35__1_), .Y(_447_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_451_), .Y(_33__1_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_448_), .B(_445_), .C(_450_), .Y(_35__2_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_35__2_), .Y(_455_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_456_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_457_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_457_), .C(_456_), .Y(_458_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_452_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_453_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_453_), .C(_35__2_), .Y(_454_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_454_), .B(_458_), .Y(_33__2_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_452_), .C(_457_), .Y(_35__3_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_462_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_463_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_464_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_462_), .B(_464_), .C(_463_), .Y(_465_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_459_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_460_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_460_), .C(vdd), .Y(_461_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_465_), .Y(_34__0_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_462_), .B(_459_), .C(_464_), .Y(_36__1_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_36__3_), .Y(_469_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_470_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_471_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_471_), .C(_470_), .Y(_472_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_466_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_467_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_466_), .B(_467_), .C(_36__3_), .Y(_468_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_468_), .B(_472_), .Y(_34__3_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_466_), .C(_471_), .Y(_32_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_36__1_), .Y(_476_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_477_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_478_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_478_), .C(_477_), .Y(_479_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_473_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_474_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_474_), .C(_36__1_), .Y(_475_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_479_), .Y(_34__1_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_473_), .C(_478_), .Y(_36__2_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_36__2_), .Y(_483_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_484_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_485_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_483_), .B(_485_), .C(_484_), .Y(_486_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_480_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_481_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_481_), .C(_36__2_), .Y(_482_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_482_), .B(_486_), .Y(_34__2_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_483_), .B(_480_), .C(_485_), .Y(_36__3_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(_37_), .Y(_487_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(w_cout_6_), .Y(_488_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_487_), .C(_488_), .Y(w_cout_7_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_39__0_), .Y(_489_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_40__0_), .B(w_cout_6_), .Y(_490_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_489_), .C(_490_), .Y(_0__28_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_39__1_), .Y(_491_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_40__1_), .Y(_492_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_491_), .C(_492_), .Y(_0__29_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_39__2_), .Y(_493_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_40__2_), .Y(_494_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_493_), .C(_494_), .Y(_0__30_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_39__3_), .Y(_495_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_40__3_), .Y(_496_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_495_), .C(_496_), .Y(_0__31_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_500_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_501_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_502_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_502_), .C(_501_), .Y(_503_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_497_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_498_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_497_), .B(_498_), .C(gnd), .Y(_499_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_503_), .Y(_39__0_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_497_), .C(_502_), .Y(_41__1_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_41__3_), .Y(_507_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_508_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_509_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_509_), .C(_508_), .Y(_510_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_504_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_505_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_504_), .B(_505_), .C(_41__3_), .Y(_506_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_510_), .Y(_39__3_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_504_), .C(_509_), .Y(_37_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_41__1_), .Y(_514_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_515_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_516_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_516_), .C(_515_), .Y(_517_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_511_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_512_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_511_), .B(_512_), .C(_41__1_), .Y(_513_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_517_), .Y(_39__1_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_511_), .C(_516_), .Y(_41__2_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(_41__2_), .Y(_521_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_522_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_523_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_523_), .C(_522_), .Y(_524_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_518_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_519_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_518_), .B(_519_), .C(_41__2_), .Y(_520_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_524_), .Y(_39__2_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_518_), .C(_523_), .Y(_41__3_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_528_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_529_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_530_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_530_), .C(_529_), .Y(_531_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_525_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_526_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_525_), .B(_526_), .C(vdd), .Y(_527_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_531_), .Y(_40__0_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_525_), .C(_530_), .Y(_42__1_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(_42__3_), .Y(_535_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_536_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_537_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_537_), .C(_536_), .Y(_538_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_532_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_533_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_532_), .B(_533_), .C(_42__3_), .Y(_534_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_538_), .Y(_40__3_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_532_), .C(_537_), .Y(_38_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_42__1_), .Y(_542_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_543_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_544_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_542_), .B(_544_), .C(_543_), .Y(_545_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_539_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_540_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_539_), .B(_540_), .C(_42__1_), .Y(_541_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_541_), .B(_545_), .Y(_40__1_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_542_), .B(_539_), .C(_544_), .Y(_42__2_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(_42__2_), .Y(_549_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_550_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_551_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(_551_), .C(_550_), .Y(_552_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_546_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_547_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_546_), .B(_547_), .C(_42__2_), .Y(_548_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_552_), .Y(_40__2_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(_546_), .C(_551_), .Y(_42__3_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(_553_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(w_cout_7_), .Y(_554_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_553_), .C(_554_), .Y(w_cout_8_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(_45__0_), .Y(_555_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_46__0_), .B(w_cout_7_), .Y(_556_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_555_), .C(_556_), .Y(_0__32_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_45__1_), .Y(_557_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_46__1_), .Y(_558_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_557_), .C(_558_), .Y(_0__33_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_45__2_), .Y(_559_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_46__2_), .Y(_560_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_559_), .C(_560_), .Y(_0__34_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(_45__3_), .Y(_561_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_46__3_), .Y(_562_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_561_), .C(_562_), .Y(_0__35_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_566_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_567_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_568_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_568_), .C(_567_), .Y(_569_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_563_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_564_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(_564_), .C(gnd), .Y(_565_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_569_), .Y(_45__0_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_563_), .C(_568_), .Y(_47__1_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(_47__3_), .Y(_573_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_574_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_575_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_575_), .C(_574_), .Y(_576_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_570_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_571_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_571_), .C(_47__3_), .Y(_572_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_576_), .Y(_45__3_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_570_), .C(_575_), .Y(_43_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(_47__1_), .Y(_580_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_581_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_582_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(_582_), .C(_581_), .Y(_583_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_577_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_578_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_578_), .C(_47__1_), .Y(_579_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_583_), .Y(_45__1_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(_577_), .C(_582_), .Y(_47__2_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(_47__2_), .Y(_587_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_588_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_589_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(_589_), .C(_588_), .Y(_590_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_584_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_585_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_585_), .C(_47__2_), .Y(_586_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_586_), .B(_590_), .Y(_45__2_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(_584_), .C(_589_), .Y(_47__3_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_594_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_595_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_596_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_594_), .B(_596_), .C(_595_), .Y(_597_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_591_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_592_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_592_), .C(vdd), .Y(_593_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_597_), .Y(_46__0_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_594_), .B(_591_), .C(_596_), .Y(_48__1_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(_48__3_), .Y(_601_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_602_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_603_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_601_), .B(_603_), .C(_602_), .Y(_604_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_598_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_599_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_598_), .B(_599_), .C(_48__3_), .Y(_600_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_604_), .Y(_46__3_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_601_), .B(_598_), .C(_603_), .Y(_44_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_48__1_), .Y(_608_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_609_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_610_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_608_), .B(_610_), .C(_609_), .Y(_611_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_605_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_606_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_606_), .C(_48__1_), .Y(_607_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_611_), .Y(_46__1_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_608_), .B(_605_), .C(_610_), .Y(_48__2_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(_48__2_), .Y(_615_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_616_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_617_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(_617_), .C(_616_), .Y(_618_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_612_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_613_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_612_), .B(_613_), .C(_48__2_), .Y(_614_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_618_), .Y(_46__2_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(_612_), .C(_617_), .Y(_48__3_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_49_), .Y(_619_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(w_cout_8_), .Y(_620_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_619_), .C(_620_), .Y(w_cout_9_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_51__0_), .Y(_621_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_52__0_), .B(w_cout_8_), .Y(_622_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_621_), .C(_622_), .Y(_0__36_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_51__1_), .Y(_623_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_52__1_), .Y(_624_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_623_), .C(_624_), .Y(_0__37_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_51__2_), .Y(_625_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_52__2_), .Y(_626_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_625_), .C(_626_), .Y(_0__38_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_51__3_), .Y(_627_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_52__3_), .Y(_628_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_627_), .C(_628_), .Y(_0__39_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_632_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_633_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_634_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_632_), .B(_634_), .C(_633_), .Y(_635_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_629_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_630_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_629_), .B(_630_), .C(gnd), .Y(_631_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_631_), .B(_635_), .Y(_51__0_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_632_), .B(_629_), .C(_634_), .Y(_53__1_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_53__3_), .Y(_639_) );
OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_640_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_641_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_641_), .C(_640_), .Y(_642_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_636_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_637_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_636_), .B(_637_), .C(_53__3_), .Y(_638_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_642_), .Y(_51__3_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_636_), .C(_641_), .Y(_49_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(_53__1_), .Y(_646_) );
OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_647_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_648_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_646_), .B(_648_), .C(_647_), .Y(_649_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_643_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_644_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_644_), .C(_53__1_), .Y(_645_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_645_), .B(_649_), .Y(_51__1_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_646_), .B(_643_), .C(_648_), .Y(_53__2_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(_53__2_), .Y(_653_) );
OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_654_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_655_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_653_), .B(_655_), .C(_654_), .Y(_656_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_650_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_651_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(_651_), .C(_53__2_), .Y(_652_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_656_), .Y(_51__2_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_653_), .B(_650_), .C(_655_), .Y(_53__3_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_660_) );
OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_661_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_662_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_660_), .B(_662_), .C(_661_), .Y(_663_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_657_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_658_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_657_), .B(_658_), .C(vdd), .Y(_659_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(_663_), .Y(_52__0_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_660_), .B(_657_), .C(_662_), .Y(_54__1_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(_54__3_), .Y(_667_) );
OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_668_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_669_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_667_), .B(_669_), .C(_668_), .Y(_670_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_664_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_665_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_665_), .C(_54__3_), .Y(_666_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_666_), .B(_670_), .Y(_52__3_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_667_), .B(_664_), .C(_669_), .Y(_50_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(_54__1_), .Y(_674_) );
OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_675_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_676_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_676_), .C(_675_), .Y(_677_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_671_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_672_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_671_), .B(_672_), .C(_54__1_), .Y(_673_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(_677_), .Y(_52__1_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_671_), .C(_676_), .Y(_54__2_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(_54__2_), .Y(_681_) );
OR2X2 OR2X2_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_682_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_683_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_681_), .B(_683_), .C(_682_), .Y(_684_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_678_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_679_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_679_), .C(_54__2_), .Y(_680_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_680_), .B(_684_), .Y(_52__2_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_681_), .B(_678_), .C(_683_), .Y(_54__3_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(_55_), .Y(_685_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(w_cout_9_), .Y(_686_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_685_), .C(_686_), .Y(w_cout_10_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(_57__0_), .Y(_687_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_58__0_), .B(w_cout_9_), .Y(_688_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_687_), .C(_688_), .Y(_0__40_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(_57__1_), .Y(_689_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_58__1_), .Y(_690_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_689_), .C(_690_), .Y(_0__41_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(_57__2_), .Y(_691_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_58__2_), .Y(_692_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_691_), .C(_692_), .Y(_0__42_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(_57__3_), .Y(_693_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_58__3_), .Y(_694_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_693_), .C(_694_), .Y(_0__43_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_698_) );
OR2X2 OR2X2_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_699_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_700_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_700_), .C(_699_), .Y(_701_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_695_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_696_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_695_), .B(_696_), .C(gnd), .Y(_697_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_697_), .B(_701_), .Y(_57__0_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_695_), .C(_700_), .Y(_59__1_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(_59__3_), .Y(_705_) );
OR2X2 OR2X2_74 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_706_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_707_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_705_), .B(_707_), .C(_706_), .Y(_708_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_702_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_703_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(_703_), .C(_59__3_), .Y(_704_) );
NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_708_), .Y(_57__3_) );
OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_705_), .B(_702_), .C(_707_), .Y(_55_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(_59__1_), .Y(_712_) );
OR2X2 OR2X2_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_713_) );
NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_714_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_712_), .B(_714_), .C(_713_), .Y(_715_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_709_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_710_) );
OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_710_), .C(_59__1_), .Y(_711_) );
NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_715_), .Y(_57__1_) );
OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_712_), .B(_709_), .C(_714_), .Y(_59__2_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(_59__2_), .Y(_719_) );
OR2X2 OR2X2_76 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_720_) );
NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_721_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(_721_), .C(_720_), .Y(_722_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_716_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_717_) );
OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_716_), .B(_717_), .C(_59__2_), .Y(_718_) );
NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_718_), .B(_722_), .Y(_57__2_) );
OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(_716_), .C(_721_), .Y(_59__3_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_726_) );
OR2X2 OR2X2_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_727_) );
NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_728_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_726_), .B(_728_), .C(_727_), .Y(_729_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_723_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_724_) );
OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_723_), .B(_724_), .C(vdd), .Y(_725_) );
NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(_729_), .Y(_58__0_) );
OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_726_), .B(_723_), .C(_728_), .Y(_60__1_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(_60__3_), .Y(_733_) );
OR2X2 OR2X2_78 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_734_) );
NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_735_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_733_), .B(_735_), .C(_734_), .Y(_736_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_730_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_731_) );
OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_730_), .B(_731_), .C(_60__3_), .Y(_732_) );
NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_736_), .Y(_58__3_) );
OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_733_), .B(_730_), .C(_735_), .Y(_56_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(_60__1_), .Y(_740_) );
OR2X2 OR2X2_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_741_) );
NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_742_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_740_), .B(_742_), .C(_741_), .Y(_743_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_737_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_738_) );
OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_737_), .B(_738_), .C(_60__1_), .Y(_739_) );
NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_739_), .B(_743_), .Y(_58__1_) );
OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_740_), .B(_737_), .C(_742_), .Y(_60__2_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(_60__2_), .Y(_747_) );
OR2X2 OR2X2_80 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_748_) );
NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_749_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_747_), .B(_749_), .C(_748_), .Y(_750_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_744_) );
AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_745_) );
OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_744_), .B(_745_), .C(_60__2_), .Y(_746_) );
NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_750_), .Y(_58__2_) );
OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_747_), .B(_744_), .C(_749_), .Y(_60__3_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(_61_), .Y(_751_) );
NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(w_cout_10_), .Y(_752_) );
OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_751_), .C(_752_), .Y(w_cout_11_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(_63__0_), .Y(_753_) );
NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_64__0_), .B(w_cout_10_), .Y(_754_) );
OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_753_), .C(_754_), .Y(_0__44_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(_63__1_), .Y(_755_) );
NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_64__1_), .Y(_756_) );
OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_755_), .C(_756_), .Y(_0__45_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(_63__2_), .Y(_757_) );
NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_64__2_), .Y(_758_) );
OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_757_), .C(_758_), .Y(_0__46_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(_63__3_), .Y(_759_) );
NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_64__3_), .Y(_760_) );
OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_759_), .C(_760_), .Y(_0__47_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_764_) );
OR2X2 OR2X2_81 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_765_) );
NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_766_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_764_), .B(_766_), .C(_765_), .Y(_767_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_761_) );
AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_762_) );
OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_761_), .B(_762_), .C(gnd), .Y(_763_) );
NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_763_), .B(_767_), .Y(_63__0_) );
OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_764_), .B(_761_), .C(_766_), .Y(_65__1_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(_65__3_), .Y(_771_) );
OR2X2 OR2X2_82 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_772_) );
NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_773_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_771_), .B(_773_), .C(_772_), .Y(_774_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_768_) );
AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_769_) );
OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_768_), .B(_769_), .C(_65__3_), .Y(_770_) );
NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_770_), .B(_774_), .Y(_63__3_) );
OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_771_), .B(_768_), .C(_773_), .Y(_61_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(_65__1_), .Y(_778_) );
OR2X2 OR2X2_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_779_) );
NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_780_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(_780_), .C(_779_), .Y(_781_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_775_) );
AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_776_) );
OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_775_), .B(_776_), .C(_65__1_), .Y(_777_) );
NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_777_), .B(_781_), .Y(_63__1_) );
OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(_775_), .C(_780_), .Y(_65__2_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(_65__2_), .Y(_785_) );
OR2X2 OR2X2_84 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_786_) );
NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_787_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_787_), .C(_786_), .Y(_788_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_782_) );
AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_783_) );
OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_782_), .B(_783_), .C(_65__2_), .Y(_784_) );
NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_784_), .B(_788_), .Y(_63__2_) );
OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_782_), .C(_787_), .Y(_65__3_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_792_) );
OR2X2 OR2X2_85 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_793_) );
NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_794_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_792_), .B(_794_), .C(_793_), .Y(_795_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_789_) );
AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_790_) );
OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_790_), .C(vdd), .Y(_791_) );
NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_791_), .B(_795_), .Y(_64__0_) );
OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_792_), .B(_789_), .C(_794_), .Y(_66__1_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(_66__3_), .Y(_799_) );
OR2X2 OR2X2_86 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_800_) );
NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_801_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_799_), .B(_801_), .C(_800_), .Y(_802_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_796_) );
AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_797_) );
OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_796_), .B(_797_), .C(_66__3_), .Y(_798_) );
NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_798_), .B(_802_), .Y(_64__3_) );
OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_799_), .B(_796_), .C(_801_), .Y(_62_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(_66__1_), .Y(_806_) );
OR2X2 OR2X2_87 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_807_) );
NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_808_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_806_), .B(_808_), .C(_807_), .Y(_809_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_803_) );
AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_804_) );
OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_803_), .B(_804_), .C(_66__1_), .Y(_805_) );
NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_805_), .B(_809_), .Y(_64__1_) );
OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_806_), .B(_803_), .C(_808_), .Y(_66__2_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(_66__2_), .Y(_813_) );
OR2X2 OR2X2_88 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_814_) );
NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_815_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_813_), .B(_815_), .C(_814_), .Y(_816_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_810_) );
AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_811_) );
OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_810_), .B(_811_), .C(_66__2_), .Y(_812_) );
NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_816_), .Y(_64__2_) );
OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_813_), .B(_810_), .C(_815_), .Y(_66__3_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(_67_), .Y(_817_) );
NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(w_cout_11_), .Y(_818_) );
OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_817_), .C(_818_), .Y(w_cout_12_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(_69__0_), .Y(_819_) );
NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_70__0_), .B(w_cout_11_), .Y(_820_) );
OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_819_), .C(_820_), .Y(_0__48_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(_69__1_), .Y(_821_) );
NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_70__1_), .Y(_822_) );
OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_821_), .C(_822_), .Y(_0__49_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(_69__2_), .Y(_823_) );
NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_70__2_), .Y(_824_) );
OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_823_), .C(_824_), .Y(_0__50_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(_69__3_), .Y(_825_) );
NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_70__3_), .Y(_826_) );
OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_825_), .C(_826_), .Y(_0__51_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_830_) );
OR2X2 OR2X2_89 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_831_) );
NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_832_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_830_), .B(_832_), .C(_831_), .Y(_833_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_827_) );
AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_828_) );
OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_827_), .B(_828_), .C(gnd), .Y(_829_) );
NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_829_), .B(_833_), .Y(_69__0_) );
OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_830_), .B(_827_), .C(_832_), .Y(_71__1_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(_71__3_), .Y(_837_) );
OR2X2 OR2X2_90 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_838_) );
NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_839_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_837_), .B(_839_), .C(_838_), .Y(_840_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_834_) );
AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_835_) );
OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_834_), .B(_835_), .C(_71__3_), .Y(_836_) );
NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_836_), .B(_840_), .Y(_69__3_) );
OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_837_), .B(_834_), .C(_839_), .Y(_67_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(_71__1_), .Y(_844_) );
OR2X2 OR2X2_91 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_845_) );
NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_846_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_844_), .B(_846_), .C(_845_), .Y(_847_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_841_) );
AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_842_) );
OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_841_), .B(_842_), .C(_71__1_), .Y(_843_) );
NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_847_), .Y(_69__1_) );
OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_844_), .B(_841_), .C(_846_), .Y(_71__2_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(_71__2_), .Y(_851_) );
OR2X2 OR2X2_92 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_852_) );
NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_853_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_851_), .B(_853_), .C(_852_), .Y(_854_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_848_) );
AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_849_) );
OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_849_), .C(_71__2_), .Y(_850_) );
NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_850_), .B(_854_), .Y(_69__2_) );
OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_851_), .B(_848_), .C(_853_), .Y(_71__3_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_858_) );
OR2X2 OR2X2_93 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_859_) );
NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_860_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_858_), .B(_860_), .C(_859_), .Y(_861_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_855_) );
AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_856_) );
OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_855_), .B(_856_), .C(vdd), .Y(_857_) );
NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_857_), .B(_861_), .Y(_70__0_) );
OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_858_), .B(_855_), .C(_860_), .Y(_72__1_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(_72__3_), .Y(_865_) );
OR2X2 OR2X2_94 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_866_) );
NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_867_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(_867_), .C(_866_), .Y(_868_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_862_) );
AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_863_) );
OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(_863_), .C(_72__3_), .Y(_864_) );
NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_864_), .B(_868_), .Y(_70__3_) );
OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(_862_), .C(_867_), .Y(_68_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(_72__1_), .Y(_872_) );
OR2X2 OR2X2_95 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_873_) );
NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_874_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_874_), .C(_873_), .Y(_875_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_869_) );
AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_870_) );
OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_869_), .B(_870_), .C(_72__1_), .Y(_871_) );
NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_871_), .B(_875_), .Y(_70__1_) );
OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_869_), .C(_874_), .Y(_72__2_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(_72__2_), .Y(_879_) );
OR2X2 OR2X2_96 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_880_) );
NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_881_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_879_), .B(_881_), .C(_880_), .Y(_882_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_876_) );
AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_877_) );
OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_876_), .B(_877_), .C(_72__2_), .Y(_878_) );
NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_878_), .B(_882_), .Y(_70__2_) );
OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_879_), .B(_876_), .C(_881_), .Y(_72__3_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(_73_), .Y(_883_) );
NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(w_cout_12_), .Y(_884_) );
OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_883_), .C(_884_), .Y(w_cout_13_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(_75__0_), .Y(_885_) );
NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_76__0_), .B(w_cout_12_), .Y(_886_) );
OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_885_), .C(_886_), .Y(_0__52_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(_75__1_), .Y(_887_) );
NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_76__1_), .Y(_888_) );
OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_887_), .C(_888_), .Y(_0__53_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(_75__2_), .Y(_889_) );
NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_76__2_), .Y(_890_) );
OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_889_), .C(_890_), .Y(_0__54_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(_75__3_), .Y(_891_) );
NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_76__3_), .Y(_892_) );
OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_891_), .C(_892_), .Y(_0__55_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_896_) );
OR2X2 OR2X2_97 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_897_) );
NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_898_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_896_), .B(_898_), .C(_897_), .Y(_899_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_893_) );
AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_894_) );
OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_893_), .B(_894_), .C(gnd), .Y(_895_) );
NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_895_), .B(_899_), .Y(_75__0_) );
OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_896_), .B(_893_), .C(_898_), .Y(_77__1_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(_77__3_), .Y(_903_) );
OR2X2 OR2X2_98 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_904_) );
NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_905_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_903_), .B(_905_), .C(_904_), .Y(_906_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_900_) );
AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_901_) );
OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_900_), .B(_901_), .C(_77__3_), .Y(_902_) );
NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_902_), .B(_906_), .Y(_75__3_) );
OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_903_), .B(_900_), .C(_905_), .Y(_73_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(_77__1_), .Y(_910_) );
OR2X2 OR2X2_99 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_911_) );
NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_912_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_912_), .C(_911_), .Y(_913_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_907_) );
AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_908_) );
OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_907_), .B(_908_), .C(_77__1_), .Y(_909_) );
NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_913_), .Y(_75__1_) );
OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_910_), .B(_907_), .C(_912_), .Y(_77__2_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(_77__2_), .Y(_917_) );
OR2X2 OR2X2_100 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_918_) );
NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_919_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_919_), .C(_918_), .Y(_920_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_914_) );
AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_915_) );
OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_914_), .B(_915_), .C(_77__2_), .Y(_916_) );
NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_916_), .B(_920_), .Y(_75__2_) );
OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_917_), .B(_914_), .C(_919_), .Y(_77__3_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_924_) );
OR2X2 OR2X2_101 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_925_) );
NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_926_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_924_), .B(_926_), .C(_925_), .Y(_927_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_921_) );
AND2X2 AND2X2_101 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_922_) );
OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_921_), .B(_922_), .C(vdd), .Y(_923_) );
NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_927_), .Y(_76__0_) );
OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_924_), .B(_921_), .C(_926_), .Y(_78__1_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(_78__3_), .Y(_931_) );
OR2X2 OR2X2_102 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_932_) );
NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_933_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_933_), .C(_932_), .Y(_934_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_928_) );
AND2X2 AND2X2_102 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_929_) );
OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_928_), .B(_929_), .C(_78__3_), .Y(_930_) );
NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_934_), .Y(_76__3_) );
OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_928_), .C(_933_), .Y(_74_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(_78__1_), .Y(_938_) );
OR2X2 OR2X2_103 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_939_) );
NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_940_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_938_), .B(_940_), .C(_939_), .Y(_941_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_935_) );
AND2X2 AND2X2_103 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_936_) );
OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(_936_), .C(_78__1_), .Y(_937_) );
NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_937_), .B(_941_), .Y(_76__1_) );
OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_938_), .B(_935_), .C(_940_), .Y(_78__2_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(_78__2_), .Y(_945_) );
OR2X2 OR2X2_104 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_946_) );
NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_947_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_945_), .B(_947_), .C(_946_), .Y(_948_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_942_) );
AND2X2 AND2X2_104 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_943_) );
OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_942_), .B(_943_), .C(_78__2_), .Y(_944_) );
NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_944_), .B(_948_), .Y(_76__2_) );
OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_945_), .B(_942_), .C(_947_), .Y(_78__3_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(_79_), .Y(_949_) );
NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(w_cout_13_), .Y(_950_) );
OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(w_cout_13_), .B(_949_), .C(_950_), .Y(w_cout_14_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(_81__0_), .Y(_951_) );
NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_82__0_), .B(w_cout_13_), .Y(_952_) );
OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(w_cout_13_), .B(_951_), .C(_952_), .Y(_0__56_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(_81__1_), .Y(_953_) );
NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(w_cout_13_), .B(_82__1_), .Y(_954_) );
OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(w_cout_13_), .B(_953_), .C(_954_), .Y(_0__57_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(_81__2_), .Y(_955_) );
NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(w_cout_13_), .B(_82__2_), .Y(_956_) );
OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(w_cout_13_), .B(_955_), .C(_956_), .Y(_0__58_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(_81__3_), .Y(_957_) );
NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(w_cout_13_), .B(_82__3_), .Y(_958_) );
OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(w_cout_13_), .B(_957_), .C(_958_), .Y(_0__59_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_962_) );
OR2X2 OR2X2_105 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_963_) );
NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_964_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_964_), .C(_963_), .Y(_965_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_959_) );
AND2X2 AND2X2_105 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_960_) );
OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_959_), .B(_960_), .C(gnd), .Y(_961_) );
NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_961_), .B(_965_), .Y(_81__0_) );
OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_959_), .C(_964_), .Y(_83__1_) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(_83__3_), .Y(_969_) );
OR2X2 OR2X2_106 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_970_) );
NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_971_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_969_), .B(_971_), .C(_970_), .Y(_972_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_966_) );
AND2X2 AND2X2_106 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_967_) );
OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_966_), .B(_967_), .C(_83__3_), .Y(_968_) );
NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_968_), .B(_972_), .Y(_81__3_) );
OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_969_), .B(_966_), .C(_971_), .Y(_79_) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(_83__1_), .Y(_976_) );
OR2X2 OR2X2_107 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_977_) );
NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_978_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(_978_), .C(_977_), .Y(_979_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_973_) );
AND2X2 AND2X2_107 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_974_) );
OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_973_), .B(_974_), .C(_83__1_), .Y(_975_) );
NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_975_), .B(_979_), .Y(_81__1_) );
OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(_973_), .C(_978_), .Y(_83__2_) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(_83__2_), .Y(_983_) );
OR2X2 OR2X2_108 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_984_) );
NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_985_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_985_), .C(_984_), .Y(_986_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_980_) );
AND2X2 AND2X2_108 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_981_) );
OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_980_), .B(_981_), .C(_83__2_), .Y(_982_) );
NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_982_), .B(_986_), .Y(_81__2_) );
OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_980_), .C(_985_), .Y(_83__3_) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_990_) );
OR2X2 OR2X2_109 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_991_) );
NAND2X1 NAND2X1_287 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_992_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_992_), .C(_991_), .Y(_993_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_987_) );
AND2X2 AND2X2_109 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_988_) );
OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_987_), .B(_988_), .C(vdd), .Y(_989_) );
NAND2X1 NAND2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_989_), .B(_993_), .Y(_82__0_) );
OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_987_), .C(_992_), .Y(_84__1_) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(_84__3_), .Y(_997_) );
OR2X2 OR2X2_110 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_998_) );
NAND2X1 NAND2X1_289 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_999_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_997_), .B(_999_), .C(_998_), .Y(_1000_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_994_) );
AND2X2 AND2X2_110 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_995_) );
OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_994_), .B(_995_), .C(_84__3_), .Y(_996_) );
NAND2X1 NAND2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_996_), .B(_1000_), .Y(_82__3_) );
OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_997_), .B(_994_), .C(_999_), .Y(_80_) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(_84__1_), .Y(_1004_) );
OR2X2 OR2X2_111 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_1005_) );
NAND2X1 NAND2X1_291 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_1006_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .B(_1006_), .C(_1005_), .Y(_1007_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_1001_) );
AND2X2 AND2X2_111 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_1002_) );
OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .B(_1002_), .C(_84__1_), .Y(_1003_) );
NAND2X1 NAND2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_1003_), .B(_1007_), .Y(_82__1_) );
OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .B(_1001_), .C(_1006_), .Y(_84__2_) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(_84__2_), .Y(_1011_) );
OR2X2 OR2X2_112 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1012_) );
NAND2X1 NAND2X1_293 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1013_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .B(_1013_), .C(_1012_), .Y(_1014_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1008_) );
AND2X2 AND2X2_112 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1009_) );
OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_1008_), .B(_1009_), .C(_84__2_), .Y(_1010_) );
NAND2X1 NAND2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1010_), .B(_1014_), .Y(_82__2_) );
OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .B(_1008_), .C(_1013_), .Y(_84__3_) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(_85_), .Y(_1015_) );
NAND2X1 NAND2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(w_cout_14_), .Y(_1016_) );
OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(w_cout_14_), .B(_1015_), .C(_1016_), .Y(w_cout_15_) );
INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(_87__0_), .Y(_1017_) );
NAND2X1 NAND2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_88__0_), .B(w_cout_14_), .Y(_1018_) );
OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(w_cout_14_), .B(_1017_), .C(_1018_), .Y(_0__60_) );
INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(_87__1_), .Y(_1019_) );
NAND2X1 NAND2X1_297 ( .gnd(gnd), .vdd(vdd), .A(w_cout_14_), .B(_88__1_), .Y(_1020_) );
OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(w_cout_14_), .B(_1019_), .C(_1020_), .Y(_0__61_) );
INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(_87__2_), .Y(_1021_) );
NAND2X1 NAND2X1_298 ( .gnd(gnd), .vdd(vdd), .A(w_cout_14_), .B(_88__2_), .Y(_1022_) );
OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(w_cout_14_), .B(_1021_), .C(_1022_), .Y(_0__62_) );
INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(_87__3_), .Y(_1023_) );
NAND2X1 NAND2X1_299 ( .gnd(gnd), .vdd(vdd), .A(w_cout_14_), .B(_88__3_), .Y(_1024_) );
OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(w_cout_14_), .B(_1023_), .C(_1024_), .Y(_0__63_) );
INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_1028_) );
OR2X2 OR2X2_113 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1029_) );
NAND2X1 NAND2X1_300 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1030_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1028_), .B(_1030_), .C(_1029_), .Y(_1031_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1025_) );
AND2X2 AND2X2_113 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1026_) );
OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .B(_1026_), .C(gnd), .Y(_1027_) );
NAND2X1 NAND2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1027_), .B(_1031_), .Y(_87__0_) );
OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1028_), .B(_1025_), .C(_1030_), .Y(_89__1_) );
INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(_89__3_), .Y(_1035_) );
OR2X2 OR2X2_114 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_1036_) );
NAND2X1 NAND2X1_302 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_1037_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .B(_1037_), .C(_1036_), .Y(_1038_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_1032_) );
AND2X2 AND2X2_114 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_1033_) );
OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_1032_), .B(_1033_), .C(_89__3_), .Y(_1034_) );
NAND2X1 NAND2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_1034_), .B(_1038_), .Y(_87__3_) );
OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .B(_1032_), .C(_1037_), .Y(_85_) );
INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(_89__1_), .Y(_1042_) );
OR2X2 OR2X2_115 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_1043_) );
NAND2X1 NAND2X1_304 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_1044_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1042_), .B(_1044_), .C(_1043_), .Y(_1045_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_1039_) );
AND2X2 AND2X2_115 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_1040_) );
OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .B(_1040_), .C(_89__1_), .Y(_1041_) );
NAND2X1 NAND2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_1041_), .B(_1045_), .Y(_87__1_) );
OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_1042_), .B(_1039_), .C(_1044_), .Y(_89__2_) );
INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(_89__2_), .Y(_1049_) );
OR2X2 OR2X2_116 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_1050_) );
NAND2X1 NAND2X1_306 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_1051_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_1051_), .C(_1050_), .Y(_1052_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_1046_) );
AND2X2 AND2X2_116 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_1047_) );
OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .B(_1047_), .C(_89__2_), .Y(_1048_) );
NAND2X1 NAND2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1048_), .B(_1052_), .Y(_87__2_) );
OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_1046_), .C(_1051_), .Y(_89__3_) );
INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_1056_) );
OR2X2 OR2X2_117 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1057_) );
NAND2X1 NAND2X1_308 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1058_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1056_), .B(_1058_), .C(_1057_), .Y(_1059_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1053_) );
AND2X2 AND2X2_117 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_1054_) );
OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_1053_), .B(_1054_), .C(vdd), .Y(_1055_) );
NAND2X1 NAND2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .B(_1059_), .Y(_88__0_) );
OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_1056_), .B(_1053_), .C(_1058_), .Y(_90__1_) );
INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(_90__3_), .Y(_1063_) );
OR2X2 OR2X2_118 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_1064_) );
NAND2X1 NAND2X1_310 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_1065_) );
NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .B(_1065_), .C(_1064_), .Y(_1066_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_1060_) );
AND2X2 AND2X2_118 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_1061_) );
OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_1060_), .B(_1061_), .C(_90__3_), .Y(_1062_) );
NAND2X1 NAND2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_1062_), .B(_1066_), .Y(_88__3_) );
OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .B(_1060_), .C(_1065_), .Y(_86_) );
INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(_90__1_), .Y(_1070_) );
OR2X2 OR2X2_119 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_1071_) );
NAND2X1 NAND2X1_312 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_1072_) );
NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .B(_1072_), .C(_1071_), .Y(_1073_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_1067_) );
AND2X2 AND2X2_119 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_1068_) );
OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .B(_1068_), .C(_90__1_), .Y(_1069_) );
NAND2X1 NAND2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .B(_1073_), .Y(_88__1_) );
OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .B(_1067_), .C(_1072_), .Y(_90__2_) );
INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(_90__2_), .Y(_1077_) );
OR2X2 OR2X2_120 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_1078_) );
NAND2X1 NAND2X1_314 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_1079_) );
NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .B(_1079_), .C(_1078_), .Y(_1080_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_1074_) );
AND2X2 AND2X2_120 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_1075_) );
OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_1074_), .B(_1075_), .C(_90__2_), .Y(_1076_) );
NAND2X1 NAND2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_1076_), .B(_1080_), .Y(_88__2_) );
OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .B(_1074_), .C(_1079_), .Y(_90__3_) );
INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_1084_) );
OR2X2 OR2X2_121 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1085_) );
NAND2X1 NAND2X1_316 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1086_) );
NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1084_), .B(_1086_), .C(_1085_), .Y(_1087_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1081_) );
AND2X2 AND2X2_121 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1082_) );
OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_1081_), .B(_1082_), .C(gnd), .Y(_1083_) );
NAND2X1 NAND2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_1083_), .B(_1087_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_1084_), .B(_1081_), .C(_1086_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_i_carry), .Y(_1091_) );
OR2X2 OR2X2_122 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_1092_) );
NAND2X1 NAND2X1_318 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_1093_) );
NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1091_), .B(_1093_), .C(_1092_), .Y(_1094_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_1088_) );
AND2X2 AND2X2_122 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_1089_) );
OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_1088_), .B(_1089_), .C(rca_inst_fa3_i_carry), .Y(_1090_) );
NAND2X1 NAND2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_1094_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_1091_), .B(_1088_), .C(_1093_), .Y(rca_inst_cout) );
INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_carry), .Y(_1098_) );
OR2X2 OR2X2_123 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1099_) );
NAND2X1 NAND2X1_320 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1100_) );
NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1098_), .B(_1100_), .C(_1099_), .Y(_1101_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1095_) );
AND2X2 AND2X2_123 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1096_) );
OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_1095_), .B(_1096_), .C(rca_inst_fa0_o_carry), .Y(_1097_) );
NAND2X1 NAND2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_1097_), .B(_1101_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_1098_), .B(_1095_), .C(_1100_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_carry), .Y(_1105_) );
OR2X2 OR2X2_124 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1106_) );
NAND2X1 NAND2X1_322 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1107_) );
NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .B(_1107_), .C(_1106_), .Y(_1108_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1102_) );
AND2X2 AND2X2_124 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1103_) );
OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1103_), .C(rca_inst_fa_1__o_carry), .Y(_1104_) );
NAND2X1 NAND2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .B(_1108_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .B(_1102_), .C(_1107_), .Y(rca_inst_fa3_i_carry) );
BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_67 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_68 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_69 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_70 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .Y(w_cout_0_) );
endmodule
