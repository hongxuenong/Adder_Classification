module CSkipA_25bit ( gnd, vdd, i_add_term1, i_add_term2, sum, cout);

input gnd, vdd;
output cout;
input [24:0] i_add_term1;
input [24:0] i_add_term2;
output [24:0] sum;

BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .Y(cout) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_sum), .Y(sum[24]) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .Y(_19_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(_19_), .Y(_20_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .Y(_21_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .B(_21_), .Y(_22_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .Y(_23_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(_23_), .Y(_24_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .Y(_25_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .B(_25_), .Y(_26_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_22_), .C(_24_), .D(_26_), .Y(_27_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_28_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_29_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_29_), .Y(_30_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_31_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_31_), .Y(_32_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_32_), .Y(_3_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_33_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_3_), .Y(_34_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_33_), .C(_34_), .Y(w_cout_1_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[4]), .Y(_35_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(_35_), .Y(_36_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .Y(_37_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[4]), .B(_37_), .Y(_38_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[5]), .Y(_39_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(_39_), .Y(_40_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .Y(_41_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[5]), .B(_41_), .Y(_42_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_38_), .C(_40_), .D(_42_), .Y(_43_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_44_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_45_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_45_), .Y(_46_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_47_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_47_), .Y(_48_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_48_), .Y(_6_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(_49_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_6_), .Y(_50_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_49_), .C(_50_), .Y(w_cout_2_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[8]), .Y(_51_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(_51_), .Y(_52_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .Y(_53_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[8]), .B(_53_), .Y(_54_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[9]), .Y(_55_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(_55_), .Y(_56_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .Y(_57_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[9]), .B(_57_), .Y(_58_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_54_), .C(_56_), .D(_58_), .Y(_59_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_60_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_61_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_61_), .Y(_62_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_63_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_63_), .Y(_64_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_64_), .Y(_9_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_65_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_9_), .Y(_66_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_65_), .C(_66_), .Y(w_cout_3_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[12]), .Y(_67_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(_67_), .Y(_68_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .Y(_69_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[12]), .B(_69_), .Y(_70_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[13]), .Y(_71_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(_71_), .Y(_72_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .Y(_73_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[13]), .B(_73_), .Y(_74_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_70_), .C(_72_), .D(_74_), .Y(_75_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_76_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_77_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_77_), .Y(_78_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_79_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_79_), .Y(_80_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_80_), .Y(_12_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(_81_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_12_), .Y(_82_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_81_), .C(_82_), .Y(w_cout_4_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[16]), .Y(_83_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(_83_), .Y(_84_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .Y(_85_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[16]), .B(_85_), .Y(_86_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[17]), .Y(_87_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(_87_), .Y(_88_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .Y(_89_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[17]), .B(_89_), .Y(_90_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_86_), .C(_88_), .D(_90_), .Y(_91_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_92_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_93_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_93_), .Y(_94_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_95_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_95_), .Y(_96_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_96_), .Y(_15_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_97_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_15_), .Y(_98_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_97_), .C(_98_), .Y(w_cout_5_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[20]), .Y(_99_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(_99_), .Y(_100_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .Y(_101_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[20]), .B(_101_), .Y(_102_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[21]), .Y(_103_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(_103_), .Y(_104_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .Y(_105_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[21]), .B(_105_), .Y(_106_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_102_), .C(_104_), .D(_106_), .Y(_107_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_108_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_109_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_109_), .Y(_110_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_111_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_111_), .Y(_112_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_112_), .Y(_18_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_113_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_18_), .Y(_114_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_113_), .C(_114_), .Y(cskip1_inst_cin) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_118_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_119_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_120_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_120_), .C(_119_), .Y(_121_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_115_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_116_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_116_), .C(gnd), .Y(_117_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_121_), .Y(_0__0_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_115_), .C(_120_), .Y(_2__1_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_2__1_), .Y(_125_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_126_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_127_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_127_), .C(_126_), .Y(_128_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_122_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_123_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_123_), .C(_2__1_), .Y(_124_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_128_), .Y(_0__1_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_122_), .C(_127_), .Y(_2__2_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_2__2_), .Y(_132_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_133_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_134_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_134_), .C(_133_), .Y(_135_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_129_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_130_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_129_), .B(_130_), .C(_2__2_), .Y(_131_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_135_), .Y(_0__2_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_129_), .C(_134_), .Y(_2__3_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_2__3_), .Y(_139_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_140_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_141_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_141_), .C(_140_), .Y(_142_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_136_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_137_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_137_), .C(_2__3_), .Y(_138_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_142_), .Y(_0__3_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_136_), .C(_141_), .Y(_1_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .Y(_146_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_147_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_148_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_148_), .C(_147_), .Y(_149_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_143_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_144_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_144_), .C(w_cout_1_), .Y(_145_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_149_), .Y(_0__4_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_143_), .C(_148_), .Y(_5__1_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_5__1_), .Y(_153_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_154_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_155_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_155_), .C(_154_), .Y(_156_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_150_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_151_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_151_), .C(_5__1_), .Y(_152_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_156_), .Y(_0__5_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_150_), .C(_155_), .Y(_5__2_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_5__2_), .Y(_160_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_161_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_162_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_162_), .C(_161_), .Y(_163_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_157_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_158_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_158_), .C(_5__2_), .Y(_159_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_159_), .B(_163_), .Y(_0__6_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_157_), .C(_162_), .Y(_5__3_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_5__3_), .Y(_167_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_168_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_169_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_169_), .C(_168_), .Y(_170_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_164_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_165_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_165_), .C(_5__3_), .Y(_166_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_170_), .Y(_0__7_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_164_), .C(_169_), .Y(_4_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .Y(_174_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_175_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_176_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_176_), .C(_175_), .Y(_177_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_171_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_172_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_172_), .C(w_cout_2_), .Y(_173_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(_177_), .Y(_0__8_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_171_), .C(_176_), .Y(_8__1_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_8__1_), .Y(_181_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_182_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_183_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_183_), .C(_182_), .Y(_184_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_178_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_179_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_179_), .C(_8__1_), .Y(_180_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_184_), .Y(_0__9_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_178_), .C(_183_), .Y(_8__2_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_8__2_), .Y(_188_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_189_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_190_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_190_), .C(_189_), .Y(_191_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_185_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_186_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_186_), .C(_8__2_), .Y(_187_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(_191_), .Y(_0__10_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_185_), .C(_190_), .Y(_8__3_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_8__3_), .Y(_195_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_196_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_197_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_197_), .C(_196_), .Y(_198_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_192_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_193_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(_193_), .C(_8__3_), .Y(_194_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_198_), .Y(_0__11_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_192_), .C(_197_), .Y(_7_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .Y(_202_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_203_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_204_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_204_), .C(_203_), .Y(_205_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_199_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_200_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_200_), .C(w_cout_3_), .Y(_201_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_205_), .Y(_0__12_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_199_), .C(_204_), .Y(_11__1_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_11__1_), .Y(_209_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_210_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_211_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_211_), .C(_210_), .Y(_212_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_206_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_207_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_207_), .C(_11__1_), .Y(_208_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_212_), .Y(_0__13_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_206_), .C(_211_), .Y(_11__2_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_11__2_), .Y(_216_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_217_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_218_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_218_), .C(_217_), .Y(_219_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_213_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_214_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_214_), .C(_11__2_), .Y(_215_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_219_), .Y(_0__14_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_213_), .C(_218_), .Y(_11__3_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_11__3_), .Y(_223_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_224_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_225_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_225_), .C(_224_), .Y(_226_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_220_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_221_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_221_), .C(_11__3_), .Y(_222_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_226_), .Y(_0__15_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_220_), .C(_225_), .Y(_10_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .Y(_230_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_231_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_232_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_232_), .C(_231_), .Y(_233_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_227_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_228_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_228_), .C(w_cout_4_), .Y(_229_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_233_), .Y(_0__16_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_227_), .C(_232_), .Y(_14__1_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_14__1_), .Y(_237_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_238_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_239_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_239_), .C(_238_), .Y(_240_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_234_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_235_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_235_), .C(_14__1_), .Y(_236_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_240_), .Y(_0__17_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_234_), .C(_239_), .Y(_14__2_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_14__2_), .Y(_244_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_245_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_246_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_246_), .C(_245_), .Y(_247_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_241_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_242_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_242_), .C(_14__2_), .Y(_243_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_247_), .Y(_0__18_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_241_), .C(_246_), .Y(_14__3_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_14__3_), .Y(_251_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_252_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_253_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_253_), .C(_252_), .Y(_254_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_248_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_249_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_249_), .C(_14__3_), .Y(_250_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_254_), .Y(_0__19_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_248_), .C(_253_), .Y(_13_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .Y(_258_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_259_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_260_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_260_), .C(_259_), .Y(_261_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_255_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_256_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_256_), .C(w_cout_5_), .Y(_257_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_261_), .Y(_0__20_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_255_), .C(_260_), .Y(_17__1_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_17__1_), .Y(_265_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_266_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_267_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_267_), .C(_266_), .Y(_268_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_262_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_263_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_263_), .C(_17__1_), .Y(_264_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_268_), .Y(_0__21_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_262_), .C(_267_), .Y(_17__2_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_17__2_), .Y(_272_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_273_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_274_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_274_), .C(_273_), .Y(_275_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_269_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_270_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_270_), .C(_17__2_), .Y(_271_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_275_), .Y(_0__22_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_269_), .C(_274_), .Y(_17__3_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_17__3_), .Y(_279_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_280_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_281_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_279_), .B(_281_), .C(_280_), .Y(_282_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_276_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_277_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_277_), .C(_17__3_), .Y(_278_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_282_), .Y(_0__23_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_279_), .B(_276_), .C(_281_), .Y(_16_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_cin), .Y(_286_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_287_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_288_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_288_), .C(_287_), .Y(_289_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_283_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_284_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_283_), .B(_284_), .C(cskip1_inst_cin), .Y(_285_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_289_), .Y(cskip1_inst_sum) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_283_), .C(_288_), .Y(cskip1_inst_rca0_w_CARRY_1_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_rca0_w_CARRY_1_), .Y(_291_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_292_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_290_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_290_), .C(_292_), .Y(cskip1_inst_rca0_w_CARRY_2_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_rca0_w_CARRY_2_), .Y(_294_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_295_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_293_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_293_), .C(_295_), .Y(cskip1_inst_rca0_w_CARRY_3_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_rca0_w_CARRY_3_), .Y(_297_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_298_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_296_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_296_), .C(_298_), .Y(cskip1_inst_cout0) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_299_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_300_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_300_), .Y(cskip1_inst_skip0_P) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_cout0), .Y(_301_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(cskip1_inst_skip0_P), .Y(_302_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_skip0_P), .B(_301_), .C(_302_), .Y(w_cout_7_) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_sum), .Y(_0__24_) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_2__0_) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .Y(_5__0_) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(_5__4_) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .Y(_8__0_) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .Y(_11__0_) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(_11__4_) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .Y(_14__0_) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .Y(_17__0_) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_17__4_) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_cin), .Y(cskip1_inst_rca0_w_CARRY_0_) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_cout0), .Y(cskip1_inst_rca0_w_CARRY_4_) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_cin), .Y(w_cout_6_) );
endmodule
