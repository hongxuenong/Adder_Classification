module csa_49bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [48:0] i_add_term1;
input [48:0] i_add_term2;
output [48:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

OR2X2 OR2X2_1 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_147_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_148_) );
NAND3X1 NAND3X1_1 ( .A(_146_), .B(_148_), .C(_147_), .Y(_149_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_143_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_144_) );
OAI21X1 OAI21X1_1 ( .A(_143_), .B(_144_), .C(gnd), .Y(_145_) );
NAND2X1 NAND2X1_2 ( .A(_145_), .B(_149_), .Y(_9__0_) );
OAI21X1 OAI21X1_2 ( .A(_146_), .B(_143_), .C(_148_), .Y(_11__1_) );
INVX1 INVX1_1 ( .A(_11__3_), .Y(_153_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_154_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_155_) );
NAND3X1 NAND3X1_2 ( .A(_153_), .B(_155_), .C(_154_), .Y(_156_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_150_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_151_) );
OAI21X1 OAI21X1_3 ( .A(_150_), .B(_151_), .C(_11__3_), .Y(_152_) );
NAND2X1 NAND2X1_4 ( .A(_152_), .B(_156_), .Y(_9__3_) );
OAI21X1 OAI21X1_4 ( .A(_153_), .B(_150_), .C(_155_), .Y(_7_) );
INVX1 INVX1_2 ( .A(_11__1_), .Y(_160_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_161_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_162_) );
NAND3X1 NAND3X1_3 ( .A(_160_), .B(_162_), .C(_161_), .Y(_163_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_157_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_158_) );
OAI21X1 OAI21X1_5 ( .A(_157_), .B(_158_), .C(_11__1_), .Y(_159_) );
NAND2X1 NAND2X1_6 ( .A(_159_), .B(_163_), .Y(_9__1_) );
OAI21X1 OAI21X1_6 ( .A(_160_), .B(_157_), .C(_162_), .Y(_11__2_) );
INVX1 INVX1_3 ( .A(_11__2_), .Y(_167_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_168_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_169_) );
NAND3X1 NAND3X1_4 ( .A(_167_), .B(_169_), .C(_168_), .Y(_170_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_164_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_165_) );
OAI21X1 OAI21X1_7 ( .A(_164_), .B(_165_), .C(_11__2_), .Y(_166_) );
NAND2X1 NAND2X1_8 ( .A(_166_), .B(_170_), .Y(_9__2_) );
OAI21X1 OAI21X1_8 ( .A(_167_), .B(_164_), .C(_169_), .Y(_11__3_) );
INVX1 INVX1_4 ( .A(vdd), .Y(_174_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_175_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_176_) );
NAND3X1 NAND3X1_5 ( .A(_174_), .B(_176_), .C(_175_), .Y(_177_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_171_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_172_) );
OAI21X1 OAI21X1_9 ( .A(_171_), .B(_172_), .C(vdd), .Y(_173_) );
NAND2X1 NAND2X1_10 ( .A(_173_), .B(_177_), .Y(_10__0_) );
OAI21X1 OAI21X1_10 ( .A(_174_), .B(_171_), .C(_176_), .Y(_12__1_) );
INVX1 INVX1_5 ( .A(_12__3_), .Y(_181_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_182_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_183_) );
NAND3X1 NAND3X1_6 ( .A(_181_), .B(_183_), .C(_182_), .Y(_184_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_178_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_179_) );
OAI21X1 OAI21X1_11 ( .A(_178_), .B(_179_), .C(_12__3_), .Y(_180_) );
NAND2X1 NAND2X1_12 ( .A(_180_), .B(_184_), .Y(_10__3_) );
OAI21X1 OAI21X1_12 ( .A(_181_), .B(_178_), .C(_183_), .Y(_8_) );
INVX1 INVX1_6 ( .A(_12__1_), .Y(_188_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_189_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_190_) );
NAND3X1 NAND3X1_7 ( .A(_188_), .B(_190_), .C(_189_), .Y(_191_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_185_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_186_) );
OAI21X1 OAI21X1_13 ( .A(_185_), .B(_186_), .C(_12__1_), .Y(_187_) );
NAND2X1 NAND2X1_14 ( .A(_187_), .B(_191_), .Y(_10__1_) );
OAI21X1 OAI21X1_14 ( .A(_188_), .B(_185_), .C(_190_), .Y(_12__2_) );
INVX1 INVX1_7 ( .A(_12__2_), .Y(_195_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_196_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_197_) );
NAND3X1 NAND3X1_8 ( .A(_195_), .B(_197_), .C(_196_), .Y(_198_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_192_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_193_) );
OAI21X1 OAI21X1_15 ( .A(_192_), .B(_193_), .C(_12__2_), .Y(_194_) );
NAND2X1 NAND2X1_16 ( .A(_194_), .B(_198_), .Y(_10__2_) );
OAI21X1 OAI21X1_16 ( .A(_195_), .B(_192_), .C(_197_), .Y(_12__3_) );
INVX1 INVX1_8 ( .A(_13_), .Y(_199_) );
NAND2X1 NAND2X1_17 ( .A(_14_), .B(w_cout_2_), .Y(_200_) );
OAI21X1 OAI21X1_17 ( .A(w_cout_2_), .B(_199_), .C(_200_), .Y(w_cout_3_) );
INVX1 INVX1_9 ( .A(_15__0_), .Y(_201_) );
NAND2X1 NAND2X1_18 ( .A(_16__0_), .B(w_cout_2_), .Y(_202_) );
OAI21X1 OAI21X1_18 ( .A(w_cout_2_), .B(_201_), .C(_202_), .Y(_0__12_) );
INVX1 INVX1_10 ( .A(_15__1_), .Y(_203_) );
NAND2X1 NAND2X1_19 ( .A(w_cout_2_), .B(_16__1_), .Y(_204_) );
OAI21X1 OAI21X1_19 ( .A(w_cout_2_), .B(_203_), .C(_204_), .Y(_0__13_) );
INVX1 INVX1_11 ( .A(_15__2_), .Y(_205_) );
NAND2X1 NAND2X1_20 ( .A(w_cout_2_), .B(_16__2_), .Y(_206_) );
OAI21X1 OAI21X1_20 ( .A(w_cout_2_), .B(_205_), .C(_206_), .Y(_0__14_) );
INVX1 INVX1_12 ( .A(_15__3_), .Y(_207_) );
NAND2X1 NAND2X1_21 ( .A(w_cout_2_), .B(_16__3_), .Y(_208_) );
OAI21X1 OAI21X1_21 ( .A(w_cout_2_), .B(_207_), .C(_208_), .Y(_0__15_) );
INVX1 INVX1_13 ( .A(gnd), .Y(_212_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_213_) );
NAND2X1 NAND2X1_22 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_214_) );
NAND3X1 NAND3X1_9 ( .A(_212_), .B(_214_), .C(_213_), .Y(_215_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_209_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_210_) );
OAI21X1 OAI21X1_22 ( .A(_209_), .B(_210_), .C(gnd), .Y(_211_) );
NAND2X1 NAND2X1_23 ( .A(_211_), .B(_215_), .Y(_15__0_) );
OAI21X1 OAI21X1_23 ( .A(_212_), .B(_209_), .C(_214_), .Y(_17__1_) );
INVX1 INVX1_14 ( .A(_17__3_), .Y(_219_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_220_) );
NAND2X1 NAND2X1_24 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_221_) );
NAND3X1 NAND3X1_10 ( .A(_219_), .B(_221_), .C(_220_), .Y(_222_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_216_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_217_) );
OAI21X1 OAI21X1_24 ( .A(_216_), .B(_217_), .C(_17__3_), .Y(_218_) );
NAND2X1 NAND2X1_25 ( .A(_218_), .B(_222_), .Y(_15__3_) );
OAI21X1 OAI21X1_25 ( .A(_219_), .B(_216_), .C(_221_), .Y(_13_) );
INVX1 INVX1_15 ( .A(_17__1_), .Y(_226_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_227_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_228_) );
NAND3X1 NAND3X1_11 ( .A(_226_), .B(_228_), .C(_227_), .Y(_229_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_223_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_224_) );
OAI21X1 OAI21X1_26 ( .A(_223_), .B(_224_), .C(_17__1_), .Y(_225_) );
NAND2X1 NAND2X1_27 ( .A(_225_), .B(_229_), .Y(_15__1_) );
OAI21X1 OAI21X1_27 ( .A(_226_), .B(_223_), .C(_228_), .Y(_17__2_) );
INVX1 INVX1_16 ( .A(_17__2_), .Y(_233_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_234_) );
NAND2X1 NAND2X1_28 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_235_) );
NAND3X1 NAND3X1_12 ( .A(_233_), .B(_235_), .C(_234_), .Y(_236_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_230_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_231_) );
OAI21X1 OAI21X1_28 ( .A(_230_), .B(_231_), .C(_17__2_), .Y(_232_) );
NAND2X1 NAND2X1_29 ( .A(_232_), .B(_236_), .Y(_15__2_) );
OAI21X1 OAI21X1_29 ( .A(_233_), .B(_230_), .C(_235_), .Y(_17__3_) );
INVX1 INVX1_17 ( .A(vdd), .Y(_240_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_241_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_242_) );
NAND3X1 NAND3X1_13 ( .A(_240_), .B(_242_), .C(_241_), .Y(_243_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_237_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_238_) );
OAI21X1 OAI21X1_30 ( .A(_237_), .B(_238_), .C(vdd), .Y(_239_) );
NAND2X1 NAND2X1_31 ( .A(_239_), .B(_243_), .Y(_16__0_) );
OAI21X1 OAI21X1_31 ( .A(_240_), .B(_237_), .C(_242_), .Y(_18__1_) );
INVX1 INVX1_18 ( .A(_18__3_), .Y(_247_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_248_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_249_) );
NAND3X1 NAND3X1_14 ( .A(_247_), .B(_249_), .C(_248_), .Y(_250_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_244_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_245_) );
OAI21X1 OAI21X1_32 ( .A(_244_), .B(_245_), .C(_18__3_), .Y(_246_) );
NAND2X1 NAND2X1_33 ( .A(_246_), .B(_250_), .Y(_16__3_) );
OAI21X1 OAI21X1_33 ( .A(_247_), .B(_244_), .C(_249_), .Y(_14_) );
INVX1 INVX1_19 ( .A(_18__1_), .Y(_254_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_255_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_256_) );
NAND3X1 NAND3X1_15 ( .A(_254_), .B(_256_), .C(_255_), .Y(_257_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_251_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_252_) );
OAI21X1 OAI21X1_34 ( .A(_251_), .B(_252_), .C(_18__1_), .Y(_253_) );
NAND2X1 NAND2X1_35 ( .A(_253_), .B(_257_), .Y(_16__1_) );
OAI21X1 OAI21X1_35 ( .A(_254_), .B(_251_), .C(_256_), .Y(_18__2_) );
INVX1 INVX1_20 ( .A(_18__2_), .Y(_261_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_262_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_263_) );
NAND3X1 NAND3X1_16 ( .A(_261_), .B(_263_), .C(_262_), .Y(_264_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_258_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_259_) );
OAI21X1 OAI21X1_36 ( .A(_258_), .B(_259_), .C(_18__2_), .Y(_260_) );
NAND2X1 NAND2X1_37 ( .A(_260_), .B(_264_), .Y(_16__2_) );
OAI21X1 OAI21X1_37 ( .A(_261_), .B(_258_), .C(_263_), .Y(_18__3_) );
INVX1 INVX1_21 ( .A(_19_), .Y(_265_) );
NAND2X1 NAND2X1_38 ( .A(_20_), .B(w_cout_3_), .Y(_266_) );
OAI21X1 OAI21X1_38 ( .A(w_cout_3_), .B(_265_), .C(_266_), .Y(w_cout_4_) );
INVX1 INVX1_22 ( .A(_21__0_), .Y(_267_) );
NAND2X1 NAND2X1_39 ( .A(_22__0_), .B(w_cout_3_), .Y(_268_) );
OAI21X1 OAI21X1_39 ( .A(w_cout_3_), .B(_267_), .C(_268_), .Y(_0__16_) );
INVX1 INVX1_23 ( .A(_21__1_), .Y(_269_) );
NAND2X1 NAND2X1_40 ( .A(w_cout_3_), .B(_22__1_), .Y(_270_) );
OAI21X1 OAI21X1_40 ( .A(w_cout_3_), .B(_269_), .C(_270_), .Y(_0__17_) );
INVX1 INVX1_24 ( .A(_21__2_), .Y(_271_) );
NAND2X1 NAND2X1_41 ( .A(w_cout_3_), .B(_22__2_), .Y(_272_) );
OAI21X1 OAI21X1_41 ( .A(w_cout_3_), .B(_271_), .C(_272_), .Y(_0__18_) );
INVX1 INVX1_25 ( .A(_21__3_), .Y(_273_) );
NAND2X1 NAND2X1_42 ( .A(w_cout_3_), .B(_22__3_), .Y(_274_) );
OAI21X1 OAI21X1_42 ( .A(w_cout_3_), .B(_273_), .C(_274_), .Y(_0__19_) );
INVX1 INVX1_26 ( .A(gnd), .Y(_278_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_279_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_280_) );
NAND3X1 NAND3X1_17 ( .A(_278_), .B(_280_), .C(_279_), .Y(_281_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_275_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_276_) );
OAI21X1 OAI21X1_43 ( .A(_275_), .B(_276_), .C(gnd), .Y(_277_) );
NAND2X1 NAND2X1_44 ( .A(_277_), .B(_281_), .Y(_21__0_) );
OAI21X1 OAI21X1_44 ( .A(_278_), .B(_275_), .C(_280_), .Y(_23__1_) );
INVX1 INVX1_27 ( .A(_23__3_), .Y(_285_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_286_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_287_) );
NAND3X1 NAND3X1_18 ( .A(_285_), .B(_287_), .C(_286_), .Y(_288_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_282_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_283_) );
OAI21X1 OAI21X1_45 ( .A(_282_), .B(_283_), .C(_23__3_), .Y(_284_) );
NAND2X1 NAND2X1_46 ( .A(_284_), .B(_288_), .Y(_21__3_) );
OAI21X1 OAI21X1_46 ( .A(_285_), .B(_282_), .C(_287_), .Y(_19_) );
INVX1 INVX1_28 ( .A(_23__1_), .Y(_292_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_293_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_294_) );
NAND3X1 NAND3X1_19 ( .A(_292_), .B(_294_), .C(_293_), .Y(_295_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_289_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_290_) );
OAI21X1 OAI21X1_47 ( .A(_289_), .B(_290_), .C(_23__1_), .Y(_291_) );
NAND2X1 NAND2X1_48 ( .A(_291_), .B(_295_), .Y(_21__1_) );
OAI21X1 OAI21X1_48 ( .A(_292_), .B(_289_), .C(_294_), .Y(_23__2_) );
INVX1 INVX1_29 ( .A(_23__2_), .Y(_299_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_300_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_301_) );
NAND3X1 NAND3X1_20 ( .A(_299_), .B(_301_), .C(_300_), .Y(_302_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_296_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_297_) );
OAI21X1 OAI21X1_49 ( .A(_296_), .B(_297_), .C(_23__2_), .Y(_298_) );
NAND2X1 NAND2X1_50 ( .A(_298_), .B(_302_), .Y(_21__2_) );
OAI21X1 OAI21X1_50 ( .A(_299_), .B(_296_), .C(_301_), .Y(_23__3_) );
INVX1 INVX1_30 ( .A(vdd), .Y(_306_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_307_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_308_) );
NAND3X1 NAND3X1_21 ( .A(_306_), .B(_308_), .C(_307_), .Y(_309_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_303_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_304_) );
OAI21X1 OAI21X1_51 ( .A(_303_), .B(_304_), .C(vdd), .Y(_305_) );
NAND2X1 NAND2X1_52 ( .A(_305_), .B(_309_), .Y(_22__0_) );
OAI21X1 OAI21X1_52 ( .A(_306_), .B(_303_), .C(_308_), .Y(_24__1_) );
INVX1 INVX1_31 ( .A(_24__3_), .Y(_313_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_314_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_315_) );
NAND3X1 NAND3X1_22 ( .A(_313_), .B(_315_), .C(_314_), .Y(_316_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_310_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_311_) );
OAI21X1 OAI21X1_53 ( .A(_310_), .B(_311_), .C(_24__3_), .Y(_312_) );
NAND2X1 NAND2X1_54 ( .A(_312_), .B(_316_), .Y(_22__3_) );
OAI21X1 OAI21X1_54 ( .A(_313_), .B(_310_), .C(_315_), .Y(_20_) );
INVX1 INVX1_32 ( .A(_24__1_), .Y(_320_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_321_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_322_) );
NAND3X1 NAND3X1_23 ( .A(_320_), .B(_322_), .C(_321_), .Y(_323_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_317_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_318_) );
OAI21X1 OAI21X1_55 ( .A(_317_), .B(_318_), .C(_24__1_), .Y(_319_) );
NAND2X1 NAND2X1_56 ( .A(_319_), .B(_323_), .Y(_22__1_) );
OAI21X1 OAI21X1_56 ( .A(_320_), .B(_317_), .C(_322_), .Y(_24__2_) );
INVX1 INVX1_33 ( .A(_24__2_), .Y(_327_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_328_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_329_) );
NAND3X1 NAND3X1_24 ( .A(_327_), .B(_329_), .C(_328_), .Y(_330_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_324_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_325_) );
OAI21X1 OAI21X1_57 ( .A(_324_), .B(_325_), .C(_24__2_), .Y(_326_) );
NAND2X1 NAND2X1_58 ( .A(_326_), .B(_330_), .Y(_22__2_) );
OAI21X1 OAI21X1_58 ( .A(_327_), .B(_324_), .C(_329_), .Y(_24__3_) );
INVX1 INVX1_34 ( .A(_25_), .Y(_331_) );
NAND2X1 NAND2X1_59 ( .A(_26_), .B(w_cout_4_), .Y(_332_) );
OAI21X1 OAI21X1_59 ( .A(w_cout_4_), .B(_331_), .C(_332_), .Y(w_cout_5_) );
INVX1 INVX1_35 ( .A(_27__0_), .Y(_333_) );
NAND2X1 NAND2X1_60 ( .A(_28__0_), .B(w_cout_4_), .Y(_334_) );
OAI21X1 OAI21X1_60 ( .A(w_cout_4_), .B(_333_), .C(_334_), .Y(_0__20_) );
INVX1 INVX1_36 ( .A(_27__1_), .Y(_335_) );
NAND2X1 NAND2X1_61 ( .A(w_cout_4_), .B(_28__1_), .Y(_336_) );
OAI21X1 OAI21X1_61 ( .A(w_cout_4_), .B(_335_), .C(_336_), .Y(_0__21_) );
INVX1 INVX1_37 ( .A(_27__2_), .Y(_337_) );
NAND2X1 NAND2X1_62 ( .A(w_cout_4_), .B(_28__2_), .Y(_338_) );
OAI21X1 OAI21X1_62 ( .A(w_cout_4_), .B(_337_), .C(_338_), .Y(_0__22_) );
INVX1 INVX1_38 ( .A(_27__3_), .Y(_339_) );
NAND2X1 NAND2X1_63 ( .A(w_cout_4_), .B(_28__3_), .Y(_340_) );
OAI21X1 OAI21X1_63 ( .A(w_cout_4_), .B(_339_), .C(_340_), .Y(_0__23_) );
INVX1 INVX1_39 ( .A(gnd), .Y(_344_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_345_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_346_) );
NAND3X1 NAND3X1_25 ( .A(_344_), .B(_346_), .C(_345_), .Y(_347_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_341_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_342_) );
OAI21X1 OAI21X1_64 ( .A(_341_), .B(_342_), .C(gnd), .Y(_343_) );
NAND2X1 NAND2X1_65 ( .A(_343_), .B(_347_), .Y(_27__0_) );
OAI21X1 OAI21X1_65 ( .A(_344_), .B(_341_), .C(_346_), .Y(_29__1_) );
INVX1 INVX1_40 ( .A(_29__3_), .Y(_351_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_352_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_353_) );
NAND3X1 NAND3X1_26 ( .A(_351_), .B(_353_), .C(_352_), .Y(_354_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_348_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_349_) );
OAI21X1 OAI21X1_66 ( .A(_348_), .B(_349_), .C(_29__3_), .Y(_350_) );
NAND2X1 NAND2X1_67 ( .A(_350_), .B(_354_), .Y(_27__3_) );
OAI21X1 OAI21X1_67 ( .A(_351_), .B(_348_), .C(_353_), .Y(_25_) );
INVX1 INVX1_41 ( .A(_29__1_), .Y(_358_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_359_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_360_) );
NAND3X1 NAND3X1_27 ( .A(_358_), .B(_360_), .C(_359_), .Y(_361_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_355_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_356_) );
OAI21X1 OAI21X1_68 ( .A(_355_), .B(_356_), .C(_29__1_), .Y(_357_) );
NAND2X1 NAND2X1_69 ( .A(_357_), .B(_361_), .Y(_27__1_) );
OAI21X1 OAI21X1_69 ( .A(_358_), .B(_355_), .C(_360_), .Y(_29__2_) );
INVX1 INVX1_42 ( .A(_29__2_), .Y(_365_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_366_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_367_) );
NAND3X1 NAND3X1_28 ( .A(_365_), .B(_367_), .C(_366_), .Y(_368_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_362_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_363_) );
OAI21X1 OAI21X1_70 ( .A(_362_), .B(_363_), .C(_29__2_), .Y(_364_) );
NAND2X1 NAND2X1_71 ( .A(_364_), .B(_368_), .Y(_27__2_) );
OAI21X1 OAI21X1_71 ( .A(_365_), .B(_362_), .C(_367_), .Y(_29__3_) );
INVX1 INVX1_43 ( .A(vdd), .Y(_372_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_373_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_374_) );
NAND3X1 NAND3X1_29 ( .A(_372_), .B(_374_), .C(_373_), .Y(_375_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_369_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_370_) );
OAI21X1 OAI21X1_72 ( .A(_369_), .B(_370_), .C(vdd), .Y(_371_) );
NAND2X1 NAND2X1_73 ( .A(_371_), .B(_375_), .Y(_28__0_) );
OAI21X1 OAI21X1_73 ( .A(_372_), .B(_369_), .C(_374_), .Y(_30__1_) );
INVX1 INVX1_44 ( .A(_30__3_), .Y(_379_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_380_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_381_) );
NAND3X1 NAND3X1_30 ( .A(_379_), .B(_381_), .C(_380_), .Y(_382_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_376_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_377_) );
OAI21X1 OAI21X1_74 ( .A(_376_), .B(_377_), .C(_30__3_), .Y(_378_) );
NAND2X1 NAND2X1_75 ( .A(_378_), .B(_382_), .Y(_28__3_) );
OAI21X1 OAI21X1_75 ( .A(_379_), .B(_376_), .C(_381_), .Y(_26_) );
INVX1 INVX1_45 ( .A(_30__1_), .Y(_386_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_387_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_388_) );
NAND3X1 NAND3X1_31 ( .A(_386_), .B(_388_), .C(_387_), .Y(_389_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_383_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_384_) );
OAI21X1 OAI21X1_76 ( .A(_383_), .B(_384_), .C(_30__1_), .Y(_385_) );
NAND2X1 NAND2X1_77 ( .A(_385_), .B(_389_), .Y(_28__1_) );
OAI21X1 OAI21X1_77 ( .A(_386_), .B(_383_), .C(_388_), .Y(_30__2_) );
INVX1 INVX1_46 ( .A(_30__2_), .Y(_393_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_394_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_395_) );
NAND3X1 NAND3X1_32 ( .A(_393_), .B(_395_), .C(_394_), .Y(_396_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_390_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_391_) );
OAI21X1 OAI21X1_78 ( .A(_390_), .B(_391_), .C(_30__2_), .Y(_392_) );
NAND2X1 NAND2X1_79 ( .A(_392_), .B(_396_), .Y(_28__2_) );
OAI21X1 OAI21X1_79 ( .A(_393_), .B(_390_), .C(_395_), .Y(_30__3_) );
INVX1 INVX1_47 ( .A(_31_), .Y(_397_) );
NAND2X1 NAND2X1_80 ( .A(_32_), .B(w_cout_5_), .Y(_398_) );
OAI21X1 OAI21X1_80 ( .A(w_cout_5_), .B(_397_), .C(_398_), .Y(w_cout_6_) );
INVX1 INVX1_48 ( .A(_33__0_), .Y(_399_) );
NAND2X1 NAND2X1_81 ( .A(_34__0_), .B(w_cout_5_), .Y(_400_) );
OAI21X1 OAI21X1_81 ( .A(w_cout_5_), .B(_399_), .C(_400_), .Y(_0__24_) );
INVX1 INVX1_49 ( .A(_33__1_), .Y(_401_) );
NAND2X1 NAND2X1_82 ( .A(w_cout_5_), .B(_34__1_), .Y(_402_) );
OAI21X1 OAI21X1_82 ( .A(w_cout_5_), .B(_401_), .C(_402_), .Y(_0__25_) );
INVX1 INVX1_50 ( .A(_33__2_), .Y(_403_) );
NAND2X1 NAND2X1_83 ( .A(w_cout_5_), .B(_34__2_), .Y(_404_) );
OAI21X1 OAI21X1_83 ( .A(w_cout_5_), .B(_403_), .C(_404_), .Y(_0__26_) );
INVX1 INVX1_51 ( .A(_33__3_), .Y(_405_) );
NAND2X1 NAND2X1_84 ( .A(w_cout_5_), .B(_34__3_), .Y(_406_) );
OAI21X1 OAI21X1_84 ( .A(w_cout_5_), .B(_405_), .C(_406_), .Y(_0__27_) );
INVX1 INVX1_52 ( .A(gnd), .Y(_410_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_411_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_412_) );
NAND3X1 NAND3X1_33 ( .A(_410_), .B(_412_), .C(_411_), .Y(_413_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_407_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_408_) );
OAI21X1 OAI21X1_85 ( .A(_407_), .B(_408_), .C(gnd), .Y(_409_) );
NAND2X1 NAND2X1_86 ( .A(_409_), .B(_413_), .Y(_33__0_) );
OAI21X1 OAI21X1_86 ( .A(_410_), .B(_407_), .C(_412_), .Y(_35__1_) );
INVX1 INVX1_53 ( .A(_35__3_), .Y(_417_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_418_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_419_) );
NAND3X1 NAND3X1_34 ( .A(_417_), .B(_419_), .C(_418_), .Y(_420_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_414_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_415_) );
OAI21X1 OAI21X1_87 ( .A(_414_), .B(_415_), .C(_35__3_), .Y(_416_) );
NAND2X1 NAND2X1_88 ( .A(_416_), .B(_420_), .Y(_33__3_) );
OAI21X1 OAI21X1_88 ( .A(_417_), .B(_414_), .C(_419_), .Y(_31_) );
INVX1 INVX1_54 ( .A(_35__1_), .Y(_424_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_425_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_426_) );
NAND3X1 NAND3X1_35 ( .A(_424_), .B(_426_), .C(_425_), .Y(_427_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_421_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_422_) );
OAI21X1 OAI21X1_89 ( .A(_421_), .B(_422_), .C(_35__1_), .Y(_423_) );
NAND2X1 NAND2X1_90 ( .A(_423_), .B(_427_), .Y(_33__1_) );
OAI21X1 OAI21X1_90 ( .A(_424_), .B(_421_), .C(_426_), .Y(_35__2_) );
INVX1 INVX1_55 ( .A(_35__2_), .Y(_431_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_432_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_433_) );
NAND3X1 NAND3X1_36 ( .A(_431_), .B(_433_), .C(_432_), .Y(_434_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_428_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_429_) );
OAI21X1 OAI21X1_91 ( .A(_428_), .B(_429_), .C(_35__2_), .Y(_430_) );
NAND2X1 NAND2X1_92 ( .A(_430_), .B(_434_), .Y(_33__2_) );
OAI21X1 OAI21X1_92 ( .A(_431_), .B(_428_), .C(_433_), .Y(_35__3_) );
INVX1 INVX1_56 ( .A(vdd), .Y(_438_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_439_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_440_) );
NAND3X1 NAND3X1_37 ( .A(_438_), .B(_440_), .C(_439_), .Y(_441_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_435_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_436_) );
OAI21X1 OAI21X1_93 ( .A(_435_), .B(_436_), .C(vdd), .Y(_437_) );
NAND2X1 NAND2X1_94 ( .A(_437_), .B(_441_), .Y(_34__0_) );
OAI21X1 OAI21X1_94 ( .A(_438_), .B(_435_), .C(_440_), .Y(_36__1_) );
INVX1 INVX1_57 ( .A(_36__3_), .Y(_445_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_446_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_447_) );
NAND3X1 NAND3X1_38 ( .A(_445_), .B(_447_), .C(_446_), .Y(_448_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_442_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_443_) );
OAI21X1 OAI21X1_95 ( .A(_442_), .B(_443_), .C(_36__3_), .Y(_444_) );
NAND2X1 NAND2X1_96 ( .A(_444_), .B(_448_), .Y(_34__3_) );
OAI21X1 OAI21X1_96 ( .A(_445_), .B(_442_), .C(_447_), .Y(_32_) );
INVX1 INVX1_58 ( .A(_36__1_), .Y(_452_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_453_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_454_) );
NAND3X1 NAND3X1_39 ( .A(_452_), .B(_454_), .C(_453_), .Y(_455_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_449_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_450_) );
OAI21X1 OAI21X1_97 ( .A(_449_), .B(_450_), .C(_36__1_), .Y(_451_) );
NAND2X1 NAND2X1_98 ( .A(_451_), .B(_455_), .Y(_34__1_) );
OAI21X1 OAI21X1_98 ( .A(_452_), .B(_449_), .C(_454_), .Y(_36__2_) );
INVX1 INVX1_59 ( .A(_36__2_), .Y(_459_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_460_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_461_) );
NAND3X1 NAND3X1_40 ( .A(_459_), .B(_461_), .C(_460_), .Y(_462_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_456_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_457_) );
OAI21X1 OAI21X1_99 ( .A(_456_), .B(_457_), .C(_36__2_), .Y(_458_) );
NAND2X1 NAND2X1_100 ( .A(_458_), .B(_462_), .Y(_34__2_) );
OAI21X1 OAI21X1_100 ( .A(_459_), .B(_456_), .C(_461_), .Y(_36__3_) );
INVX1 INVX1_60 ( .A(_37_), .Y(_463_) );
NAND2X1 NAND2X1_101 ( .A(_38_), .B(w_cout_6_), .Y(_464_) );
OAI21X1 OAI21X1_101 ( .A(w_cout_6_), .B(_463_), .C(_464_), .Y(w_cout_7_) );
INVX1 INVX1_61 ( .A(_39__0_), .Y(_465_) );
NAND2X1 NAND2X1_102 ( .A(_40__0_), .B(w_cout_6_), .Y(_466_) );
OAI21X1 OAI21X1_102 ( .A(w_cout_6_), .B(_465_), .C(_466_), .Y(_0__28_) );
INVX1 INVX1_62 ( .A(_39__1_), .Y(_467_) );
NAND2X1 NAND2X1_103 ( .A(w_cout_6_), .B(_40__1_), .Y(_468_) );
OAI21X1 OAI21X1_103 ( .A(w_cout_6_), .B(_467_), .C(_468_), .Y(_0__29_) );
INVX1 INVX1_63 ( .A(_39__2_), .Y(_469_) );
NAND2X1 NAND2X1_104 ( .A(w_cout_6_), .B(_40__2_), .Y(_470_) );
OAI21X1 OAI21X1_104 ( .A(w_cout_6_), .B(_469_), .C(_470_), .Y(_0__30_) );
INVX1 INVX1_64 ( .A(_39__3_), .Y(_471_) );
NAND2X1 NAND2X1_105 ( .A(w_cout_6_), .B(_40__3_), .Y(_472_) );
OAI21X1 OAI21X1_105 ( .A(w_cout_6_), .B(_471_), .C(_472_), .Y(_0__31_) );
INVX1 INVX1_65 ( .A(gnd), .Y(_476_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_477_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_478_) );
NAND3X1 NAND3X1_41 ( .A(_476_), .B(_478_), .C(_477_), .Y(_479_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_473_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_474_) );
OAI21X1 OAI21X1_106 ( .A(_473_), .B(_474_), .C(gnd), .Y(_475_) );
NAND2X1 NAND2X1_107 ( .A(_475_), .B(_479_), .Y(_39__0_) );
OAI21X1 OAI21X1_107 ( .A(_476_), .B(_473_), .C(_478_), .Y(_41__1_) );
INVX1 INVX1_66 ( .A(_41__3_), .Y(_483_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_484_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_485_) );
NAND3X1 NAND3X1_42 ( .A(_483_), .B(_485_), .C(_484_), .Y(_486_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_480_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_481_) );
OAI21X1 OAI21X1_108 ( .A(_480_), .B(_481_), .C(_41__3_), .Y(_482_) );
NAND2X1 NAND2X1_109 ( .A(_482_), .B(_486_), .Y(_39__3_) );
OAI21X1 OAI21X1_109 ( .A(_483_), .B(_480_), .C(_485_), .Y(_37_) );
INVX1 INVX1_67 ( .A(_41__1_), .Y(_490_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_491_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_492_) );
NAND3X1 NAND3X1_43 ( .A(_490_), .B(_492_), .C(_491_), .Y(_493_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_487_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_488_) );
OAI21X1 OAI21X1_110 ( .A(_487_), .B(_488_), .C(_41__1_), .Y(_489_) );
NAND2X1 NAND2X1_111 ( .A(_489_), .B(_493_), .Y(_39__1_) );
OAI21X1 OAI21X1_111 ( .A(_490_), .B(_487_), .C(_492_), .Y(_41__2_) );
INVX1 INVX1_68 ( .A(_41__2_), .Y(_497_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_498_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_499_) );
NAND3X1 NAND3X1_44 ( .A(_497_), .B(_499_), .C(_498_), .Y(_500_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_494_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_495_) );
OAI21X1 OAI21X1_112 ( .A(_494_), .B(_495_), .C(_41__2_), .Y(_496_) );
NAND2X1 NAND2X1_113 ( .A(_496_), .B(_500_), .Y(_39__2_) );
OAI21X1 OAI21X1_113 ( .A(_497_), .B(_494_), .C(_499_), .Y(_41__3_) );
INVX1 INVX1_69 ( .A(vdd), .Y(_504_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_505_) );
NAND2X1 NAND2X1_114 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_506_) );
NAND3X1 NAND3X1_45 ( .A(_504_), .B(_506_), .C(_505_), .Y(_507_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_501_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_502_) );
OAI21X1 OAI21X1_114 ( .A(_501_), .B(_502_), .C(vdd), .Y(_503_) );
NAND2X1 NAND2X1_115 ( .A(_503_), .B(_507_), .Y(_40__0_) );
OAI21X1 OAI21X1_115 ( .A(_504_), .B(_501_), .C(_506_), .Y(_42__1_) );
INVX1 INVX1_70 ( .A(_42__3_), .Y(_511_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_512_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_513_) );
NAND3X1 NAND3X1_46 ( .A(_511_), .B(_513_), .C(_512_), .Y(_514_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_508_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_509_) );
OAI21X1 OAI21X1_116 ( .A(_508_), .B(_509_), .C(_42__3_), .Y(_510_) );
NAND2X1 NAND2X1_117 ( .A(_510_), .B(_514_), .Y(_40__3_) );
OAI21X1 OAI21X1_117 ( .A(_511_), .B(_508_), .C(_513_), .Y(_38_) );
INVX1 INVX1_71 ( .A(_42__1_), .Y(_518_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_519_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_520_) );
NAND3X1 NAND3X1_47 ( .A(_518_), .B(_520_), .C(_519_), .Y(_521_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_515_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_516_) );
OAI21X1 OAI21X1_118 ( .A(_515_), .B(_516_), .C(_42__1_), .Y(_517_) );
NAND2X1 NAND2X1_119 ( .A(_517_), .B(_521_), .Y(_40__1_) );
OAI21X1 OAI21X1_119 ( .A(_518_), .B(_515_), .C(_520_), .Y(_42__2_) );
INVX1 INVX1_72 ( .A(_42__2_), .Y(_525_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_526_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_527_) );
NAND3X1 NAND3X1_48 ( .A(_525_), .B(_527_), .C(_526_), .Y(_528_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_522_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_523_) );
OAI21X1 OAI21X1_120 ( .A(_522_), .B(_523_), .C(_42__2_), .Y(_524_) );
NAND2X1 NAND2X1_121 ( .A(_524_), .B(_528_), .Y(_40__2_) );
OAI21X1 OAI21X1_121 ( .A(_525_), .B(_522_), .C(_527_), .Y(_42__3_) );
INVX1 INVX1_73 ( .A(_43_), .Y(_529_) );
NAND2X1 NAND2X1_122 ( .A(_44_), .B(w_cout_7_), .Y(_530_) );
OAI21X1 OAI21X1_122 ( .A(w_cout_7_), .B(_529_), .C(_530_), .Y(w_cout_8_) );
INVX1 INVX1_74 ( .A(_45__0_), .Y(_531_) );
NAND2X1 NAND2X1_123 ( .A(_46__0_), .B(w_cout_7_), .Y(_532_) );
OAI21X1 OAI21X1_123 ( .A(w_cout_7_), .B(_531_), .C(_532_), .Y(_0__32_) );
INVX1 INVX1_75 ( .A(_45__1_), .Y(_533_) );
NAND2X1 NAND2X1_124 ( .A(w_cout_7_), .B(_46__1_), .Y(_534_) );
OAI21X1 OAI21X1_124 ( .A(w_cout_7_), .B(_533_), .C(_534_), .Y(_0__33_) );
INVX1 INVX1_76 ( .A(_45__2_), .Y(_535_) );
NAND2X1 NAND2X1_125 ( .A(w_cout_7_), .B(_46__2_), .Y(_536_) );
OAI21X1 OAI21X1_125 ( .A(w_cout_7_), .B(_535_), .C(_536_), .Y(_0__34_) );
INVX1 INVX1_77 ( .A(_45__3_), .Y(_537_) );
NAND2X1 NAND2X1_126 ( .A(w_cout_7_), .B(_46__3_), .Y(_538_) );
OAI21X1 OAI21X1_126 ( .A(w_cout_7_), .B(_537_), .C(_538_), .Y(_0__35_) );
INVX1 INVX1_78 ( .A(gnd), .Y(_542_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_543_) );
NAND2X1 NAND2X1_127 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_544_) );
NAND3X1 NAND3X1_49 ( .A(_542_), .B(_544_), .C(_543_), .Y(_545_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_539_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_540_) );
OAI21X1 OAI21X1_127 ( .A(_539_), .B(_540_), .C(gnd), .Y(_541_) );
NAND2X1 NAND2X1_128 ( .A(_541_), .B(_545_), .Y(_45__0_) );
OAI21X1 OAI21X1_128 ( .A(_542_), .B(_539_), .C(_544_), .Y(_47__1_) );
INVX1 INVX1_79 ( .A(_47__3_), .Y(_549_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_550_) );
NAND2X1 NAND2X1_129 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_551_) );
NAND3X1 NAND3X1_50 ( .A(_549_), .B(_551_), .C(_550_), .Y(_552_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_546_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_547_) );
OAI21X1 OAI21X1_129 ( .A(_546_), .B(_547_), .C(_47__3_), .Y(_548_) );
NAND2X1 NAND2X1_130 ( .A(_548_), .B(_552_), .Y(_45__3_) );
OAI21X1 OAI21X1_130 ( .A(_549_), .B(_546_), .C(_551_), .Y(_43_) );
INVX1 INVX1_80 ( .A(_47__1_), .Y(_556_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_557_) );
NAND2X1 NAND2X1_131 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_558_) );
NAND3X1 NAND3X1_51 ( .A(_556_), .B(_558_), .C(_557_), .Y(_559_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_553_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_554_) );
OAI21X1 OAI21X1_131 ( .A(_553_), .B(_554_), .C(_47__1_), .Y(_555_) );
NAND2X1 NAND2X1_132 ( .A(_555_), .B(_559_), .Y(_45__1_) );
OAI21X1 OAI21X1_132 ( .A(_556_), .B(_553_), .C(_558_), .Y(_47__2_) );
INVX1 INVX1_81 ( .A(_47__2_), .Y(_563_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_564_) );
NAND2X1 NAND2X1_133 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_565_) );
NAND3X1 NAND3X1_52 ( .A(_563_), .B(_565_), .C(_564_), .Y(_566_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_560_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_561_) );
OAI21X1 OAI21X1_133 ( .A(_560_), .B(_561_), .C(_47__2_), .Y(_562_) );
NAND2X1 NAND2X1_134 ( .A(_562_), .B(_566_), .Y(_45__2_) );
OAI21X1 OAI21X1_134 ( .A(_563_), .B(_560_), .C(_565_), .Y(_47__3_) );
INVX1 INVX1_82 ( .A(vdd), .Y(_570_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_571_) );
NAND2X1 NAND2X1_135 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_572_) );
NAND3X1 NAND3X1_53 ( .A(_570_), .B(_572_), .C(_571_), .Y(_573_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_567_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_568_) );
OAI21X1 OAI21X1_135 ( .A(_567_), .B(_568_), .C(vdd), .Y(_569_) );
NAND2X1 NAND2X1_136 ( .A(_569_), .B(_573_), .Y(_46__0_) );
OAI21X1 OAI21X1_136 ( .A(_570_), .B(_567_), .C(_572_), .Y(_48__1_) );
INVX1 INVX1_83 ( .A(_48__3_), .Y(_577_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_578_) );
NAND2X1 NAND2X1_137 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_579_) );
NAND3X1 NAND3X1_54 ( .A(_577_), .B(_579_), .C(_578_), .Y(_580_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_574_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_575_) );
OAI21X1 OAI21X1_137 ( .A(_574_), .B(_575_), .C(_48__3_), .Y(_576_) );
NAND2X1 NAND2X1_138 ( .A(_576_), .B(_580_), .Y(_46__3_) );
OAI21X1 OAI21X1_138 ( .A(_577_), .B(_574_), .C(_579_), .Y(_44_) );
INVX1 INVX1_84 ( .A(_48__1_), .Y(_584_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_585_) );
NAND2X1 NAND2X1_139 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_586_) );
NAND3X1 NAND3X1_55 ( .A(_584_), .B(_586_), .C(_585_), .Y(_587_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_581_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_582_) );
OAI21X1 OAI21X1_139 ( .A(_581_), .B(_582_), .C(_48__1_), .Y(_583_) );
NAND2X1 NAND2X1_140 ( .A(_583_), .B(_587_), .Y(_46__1_) );
OAI21X1 OAI21X1_140 ( .A(_584_), .B(_581_), .C(_586_), .Y(_48__2_) );
INVX1 INVX1_85 ( .A(_48__2_), .Y(_591_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_592_) );
NAND2X1 NAND2X1_141 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_593_) );
NAND3X1 NAND3X1_56 ( .A(_591_), .B(_593_), .C(_592_), .Y(_594_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_588_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_589_) );
OAI21X1 OAI21X1_141 ( .A(_588_), .B(_589_), .C(_48__2_), .Y(_590_) );
NAND2X1 NAND2X1_142 ( .A(_590_), .B(_594_), .Y(_46__2_) );
OAI21X1 OAI21X1_142 ( .A(_591_), .B(_588_), .C(_593_), .Y(_48__3_) );
INVX1 INVX1_86 ( .A(_49_), .Y(_595_) );
NAND2X1 NAND2X1_143 ( .A(_50_), .B(w_cout_8_), .Y(_596_) );
OAI21X1 OAI21X1_143 ( .A(w_cout_8_), .B(_595_), .C(_596_), .Y(w_cout_9_) );
INVX1 INVX1_87 ( .A(_51__0_), .Y(_597_) );
NAND2X1 NAND2X1_144 ( .A(_52__0_), .B(w_cout_8_), .Y(_598_) );
OAI21X1 OAI21X1_144 ( .A(w_cout_8_), .B(_597_), .C(_598_), .Y(_0__36_) );
INVX1 INVX1_88 ( .A(_51__1_), .Y(_599_) );
NAND2X1 NAND2X1_145 ( .A(w_cout_8_), .B(_52__1_), .Y(_600_) );
OAI21X1 OAI21X1_145 ( .A(w_cout_8_), .B(_599_), .C(_600_), .Y(_0__37_) );
INVX1 INVX1_89 ( .A(_51__2_), .Y(_601_) );
NAND2X1 NAND2X1_146 ( .A(w_cout_8_), .B(_52__2_), .Y(_602_) );
OAI21X1 OAI21X1_146 ( .A(w_cout_8_), .B(_601_), .C(_602_), .Y(_0__38_) );
INVX1 INVX1_90 ( .A(_51__3_), .Y(_603_) );
NAND2X1 NAND2X1_147 ( .A(w_cout_8_), .B(_52__3_), .Y(_604_) );
OAI21X1 OAI21X1_147 ( .A(w_cout_8_), .B(_603_), .C(_604_), .Y(_0__39_) );
INVX1 INVX1_91 ( .A(gnd), .Y(_608_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_609_) );
NAND2X1 NAND2X1_148 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_610_) );
NAND3X1 NAND3X1_57 ( .A(_608_), .B(_610_), .C(_609_), .Y(_611_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_605_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_606_) );
OAI21X1 OAI21X1_148 ( .A(_605_), .B(_606_), .C(gnd), .Y(_607_) );
NAND2X1 NAND2X1_149 ( .A(_607_), .B(_611_), .Y(_51__0_) );
OAI21X1 OAI21X1_149 ( .A(_608_), .B(_605_), .C(_610_), .Y(_53__1_) );
INVX1 INVX1_92 ( .A(_53__3_), .Y(_615_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_616_) );
NAND2X1 NAND2X1_150 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_617_) );
NAND3X1 NAND3X1_58 ( .A(_615_), .B(_617_), .C(_616_), .Y(_618_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_612_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_613_) );
OAI21X1 OAI21X1_150 ( .A(_612_), .B(_613_), .C(_53__3_), .Y(_614_) );
NAND2X1 NAND2X1_151 ( .A(_614_), .B(_618_), .Y(_51__3_) );
OAI21X1 OAI21X1_151 ( .A(_615_), .B(_612_), .C(_617_), .Y(_49_) );
INVX1 INVX1_93 ( .A(_53__1_), .Y(_622_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_623_) );
NAND2X1 NAND2X1_152 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_624_) );
NAND3X1 NAND3X1_59 ( .A(_622_), .B(_624_), .C(_623_), .Y(_625_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_619_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_620_) );
OAI21X1 OAI21X1_152 ( .A(_619_), .B(_620_), .C(_53__1_), .Y(_621_) );
NAND2X1 NAND2X1_153 ( .A(_621_), .B(_625_), .Y(_51__1_) );
OAI21X1 OAI21X1_153 ( .A(_622_), .B(_619_), .C(_624_), .Y(_53__2_) );
INVX1 INVX1_94 ( .A(_53__2_), .Y(_629_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_630_) );
NAND2X1 NAND2X1_154 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_631_) );
NAND3X1 NAND3X1_60 ( .A(_629_), .B(_631_), .C(_630_), .Y(_632_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_626_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_627_) );
OAI21X1 OAI21X1_154 ( .A(_626_), .B(_627_), .C(_53__2_), .Y(_628_) );
NAND2X1 NAND2X1_155 ( .A(_628_), .B(_632_), .Y(_51__2_) );
OAI21X1 OAI21X1_155 ( .A(_629_), .B(_626_), .C(_631_), .Y(_53__3_) );
INVX1 INVX1_95 ( .A(vdd), .Y(_636_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_637_) );
NAND2X1 NAND2X1_156 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_638_) );
NAND3X1 NAND3X1_61 ( .A(_636_), .B(_638_), .C(_637_), .Y(_639_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_633_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_634_) );
OAI21X1 OAI21X1_156 ( .A(_633_), .B(_634_), .C(vdd), .Y(_635_) );
NAND2X1 NAND2X1_157 ( .A(_635_), .B(_639_), .Y(_52__0_) );
OAI21X1 OAI21X1_157 ( .A(_636_), .B(_633_), .C(_638_), .Y(_54__1_) );
INVX1 INVX1_96 ( .A(_54__3_), .Y(_643_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_644_) );
NAND2X1 NAND2X1_158 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_645_) );
NAND3X1 NAND3X1_62 ( .A(_643_), .B(_645_), .C(_644_), .Y(_646_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_640_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_641_) );
OAI21X1 OAI21X1_158 ( .A(_640_), .B(_641_), .C(_54__3_), .Y(_642_) );
NAND2X1 NAND2X1_159 ( .A(_642_), .B(_646_), .Y(_52__3_) );
OAI21X1 OAI21X1_159 ( .A(_643_), .B(_640_), .C(_645_), .Y(_50_) );
INVX1 INVX1_97 ( .A(_54__1_), .Y(_650_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_651_) );
NAND2X1 NAND2X1_160 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_652_) );
NAND3X1 NAND3X1_63 ( .A(_650_), .B(_652_), .C(_651_), .Y(_653_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_647_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_648_) );
OAI21X1 OAI21X1_160 ( .A(_647_), .B(_648_), .C(_54__1_), .Y(_649_) );
NAND2X1 NAND2X1_161 ( .A(_649_), .B(_653_), .Y(_52__1_) );
OAI21X1 OAI21X1_161 ( .A(_650_), .B(_647_), .C(_652_), .Y(_54__2_) );
INVX1 INVX1_98 ( .A(_54__2_), .Y(_657_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_658_) );
NAND2X1 NAND2X1_162 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_659_) );
NAND3X1 NAND3X1_64 ( .A(_657_), .B(_659_), .C(_658_), .Y(_660_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_654_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_655_) );
OAI21X1 OAI21X1_162 ( .A(_654_), .B(_655_), .C(_54__2_), .Y(_656_) );
NAND2X1 NAND2X1_163 ( .A(_656_), .B(_660_), .Y(_52__2_) );
OAI21X1 OAI21X1_163 ( .A(_657_), .B(_654_), .C(_659_), .Y(_54__3_) );
INVX1 INVX1_99 ( .A(_55_), .Y(_661_) );
NAND2X1 NAND2X1_164 ( .A(_56_), .B(w_cout_9_), .Y(_662_) );
OAI21X1 OAI21X1_164 ( .A(w_cout_9_), .B(_661_), .C(_662_), .Y(w_cout_10_) );
INVX1 INVX1_100 ( .A(_57__0_), .Y(_663_) );
NAND2X1 NAND2X1_165 ( .A(_58__0_), .B(w_cout_9_), .Y(_664_) );
OAI21X1 OAI21X1_165 ( .A(w_cout_9_), .B(_663_), .C(_664_), .Y(_0__40_) );
INVX1 INVX1_101 ( .A(_57__1_), .Y(_665_) );
NAND2X1 NAND2X1_166 ( .A(w_cout_9_), .B(_58__1_), .Y(_666_) );
OAI21X1 OAI21X1_166 ( .A(w_cout_9_), .B(_665_), .C(_666_), .Y(_0__41_) );
INVX1 INVX1_102 ( .A(_57__2_), .Y(_667_) );
NAND2X1 NAND2X1_167 ( .A(w_cout_9_), .B(_58__2_), .Y(_668_) );
OAI21X1 OAI21X1_167 ( .A(w_cout_9_), .B(_667_), .C(_668_), .Y(_0__42_) );
INVX1 INVX1_103 ( .A(_57__3_), .Y(_669_) );
NAND2X1 NAND2X1_168 ( .A(w_cout_9_), .B(_58__3_), .Y(_670_) );
OAI21X1 OAI21X1_168 ( .A(w_cout_9_), .B(_669_), .C(_670_), .Y(_0__43_) );
INVX1 INVX1_104 ( .A(gnd), .Y(_674_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_675_) );
NAND2X1 NAND2X1_169 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_676_) );
NAND3X1 NAND3X1_65 ( .A(_674_), .B(_676_), .C(_675_), .Y(_677_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_671_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_672_) );
OAI21X1 OAI21X1_169 ( .A(_671_), .B(_672_), .C(gnd), .Y(_673_) );
NAND2X1 NAND2X1_170 ( .A(_673_), .B(_677_), .Y(_57__0_) );
OAI21X1 OAI21X1_170 ( .A(_674_), .B(_671_), .C(_676_), .Y(_59__1_) );
INVX1 INVX1_105 ( .A(_59__3_), .Y(_681_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_682_) );
NAND2X1 NAND2X1_171 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_683_) );
NAND3X1 NAND3X1_66 ( .A(_681_), .B(_683_), .C(_682_), .Y(_684_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_678_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_679_) );
OAI21X1 OAI21X1_171 ( .A(_678_), .B(_679_), .C(_59__3_), .Y(_680_) );
NAND2X1 NAND2X1_172 ( .A(_680_), .B(_684_), .Y(_57__3_) );
OAI21X1 OAI21X1_172 ( .A(_681_), .B(_678_), .C(_683_), .Y(_55_) );
INVX1 INVX1_106 ( .A(_59__1_), .Y(_688_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_689_) );
NAND2X1 NAND2X1_173 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_690_) );
NAND3X1 NAND3X1_67 ( .A(_688_), .B(_690_), .C(_689_), .Y(_691_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_685_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_686_) );
OAI21X1 OAI21X1_173 ( .A(_685_), .B(_686_), .C(_59__1_), .Y(_687_) );
NAND2X1 NAND2X1_174 ( .A(_687_), .B(_691_), .Y(_57__1_) );
OAI21X1 OAI21X1_174 ( .A(_688_), .B(_685_), .C(_690_), .Y(_59__2_) );
INVX1 INVX1_107 ( .A(_59__2_), .Y(_695_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_696_) );
NAND2X1 NAND2X1_175 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_697_) );
NAND3X1 NAND3X1_68 ( .A(_695_), .B(_697_), .C(_696_), .Y(_698_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_692_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_693_) );
OAI21X1 OAI21X1_175 ( .A(_692_), .B(_693_), .C(_59__2_), .Y(_694_) );
NAND2X1 NAND2X1_176 ( .A(_694_), .B(_698_), .Y(_57__2_) );
OAI21X1 OAI21X1_176 ( .A(_695_), .B(_692_), .C(_697_), .Y(_59__3_) );
INVX1 INVX1_108 ( .A(vdd), .Y(_702_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_703_) );
NAND2X1 NAND2X1_177 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_704_) );
NAND3X1 NAND3X1_69 ( .A(_702_), .B(_704_), .C(_703_), .Y(_705_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_699_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_700_) );
OAI21X1 OAI21X1_177 ( .A(_699_), .B(_700_), .C(vdd), .Y(_701_) );
NAND2X1 NAND2X1_178 ( .A(_701_), .B(_705_), .Y(_58__0_) );
OAI21X1 OAI21X1_178 ( .A(_702_), .B(_699_), .C(_704_), .Y(_60__1_) );
INVX1 INVX1_109 ( .A(_60__3_), .Y(_709_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_710_) );
NAND2X1 NAND2X1_179 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_711_) );
NAND3X1 NAND3X1_70 ( .A(_709_), .B(_711_), .C(_710_), .Y(_712_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_706_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_707_) );
OAI21X1 OAI21X1_179 ( .A(_706_), .B(_707_), .C(_60__3_), .Y(_708_) );
NAND2X1 NAND2X1_180 ( .A(_708_), .B(_712_), .Y(_58__3_) );
OAI21X1 OAI21X1_180 ( .A(_709_), .B(_706_), .C(_711_), .Y(_56_) );
INVX1 INVX1_110 ( .A(_60__1_), .Y(_716_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_717_) );
NAND2X1 NAND2X1_181 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_718_) );
NAND3X1 NAND3X1_71 ( .A(_716_), .B(_718_), .C(_717_), .Y(_719_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_713_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_714_) );
OAI21X1 OAI21X1_181 ( .A(_713_), .B(_714_), .C(_60__1_), .Y(_715_) );
NAND2X1 NAND2X1_182 ( .A(_715_), .B(_719_), .Y(_58__1_) );
OAI21X1 OAI21X1_182 ( .A(_716_), .B(_713_), .C(_718_), .Y(_60__2_) );
INVX1 INVX1_111 ( .A(_60__2_), .Y(_723_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_724_) );
NAND2X1 NAND2X1_183 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_725_) );
NAND3X1 NAND3X1_72 ( .A(_723_), .B(_725_), .C(_724_), .Y(_726_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_720_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_721_) );
OAI21X1 OAI21X1_183 ( .A(_720_), .B(_721_), .C(_60__2_), .Y(_722_) );
NAND2X1 NAND2X1_184 ( .A(_722_), .B(_726_), .Y(_58__2_) );
OAI21X1 OAI21X1_184 ( .A(_723_), .B(_720_), .C(_725_), .Y(_60__3_) );
INVX1 INVX1_112 ( .A(_61_), .Y(_727_) );
NAND2X1 NAND2X1_185 ( .A(_62_), .B(w_cout_10_), .Y(_728_) );
OAI21X1 OAI21X1_185 ( .A(w_cout_10_), .B(_727_), .C(_728_), .Y(csa_inst_cin) );
INVX1 INVX1_113 ( .A(_63__0_), .Y(_729_) );
NAND2X1 NAND2X1_186 ( .A(_64__0_), .B(w_cout_10_), .Y(_730_) );
OAI21X1 OAI21X1_186 ( .A(w_cout_10_), .B(_729_), .C(_730_), .Y(_0__44_) );
INVX1 INVX1_114 ( .A(_63__1_), .Y(_731_) );
NAND2X1 NAND2X1_187 ( .A(w_cout_10_), .B(_64__1_), .Y(_732_) );
OAI21X1 OAI21X1_187 ( .A(w_cout_10_), .B(_731_), .C(_732_), .Y(_0__45_) );
INVX1 INVX1_115 ( .A(_63__2_), .Y(_733_) );
NAND2X1 NAND2X1_188 ( .A(w_cout_10_), .B(_64__2_), .Y(_734_) );
OAI21X1 OAI21X1_188 ( .A(w_cout_10_), .B(_733_), .C(_734_), .Y(_0__46_) );
INVX1 INVX1_116 ( .A(_63__3_), .Y(_735_) );
NAND2X1 NAND2X1_189 ( .A(w_cout_10_), .B(_64__3_), .Y(_736_) );
OAI21X1 OAI21X1_189 ( .A(w_cout_10_), .B(_735_), .C(_736_), .Y(_0__47_) );
INVX1 INVX1_117 ( .A(gnd), .Y(_740_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_741_) );
NAND2X1 NAND2X1_190 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_742_) );
NAND3X1 NAND3X1_73 ( .A(_740_), .B(_742_), .C(_741_), .Y(_743_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_737_) );
AND2X2 AND2X2_73 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_738_) );
OAI21X1 OAI21X1_190 ( .A(_737_), .B(_738_), .C(gnd), .Y(_739_) );
NAND2X1 NAND2X1_191 ( .A(_739_), .B(_743_), .Y(_63__0_) );
OAI21X1 OAI21X1_191 ( .A(_740_), .B(_737_), .C(_742_), .Y(_65__1_) );
INVX1 INVX1_118 ( .A(_65__3_), .Y(_747_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_748_) );
NAND2X1 NAND2X1_192 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_749_) );
NAND3X1 NAND3X1_74 ( .A(_747_), .B(_749_), .C(_748_), .Y(_750_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_744_) );
AND2X2 AND2X2_74 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_745_) );
OAI21X1 OAI21X1_192 ( .A(_744_), .B(_745_), .C(_65__3_), .Y(_746_) );
NAND2X1 NAND2X1_193 ( .A(_746_), .B(_750_), .Y(_63__3_) );
OAI21X1 OAI21X1_193 ( .A(_747_), .B(_744_), .C(_749_), .Y(_61_) );
INVX1 INVX1_119 ( .A(_65__1_), .Y(_754_) );
OR2X2 OR2X2_75 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_755_) );
NAND2X1 NAND2X1_194 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_756_) );
NAND3X1 NAND3X1_75 ( .A(_754_), .B(_756_), .C(_755_), .Y(_757_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_751_) );
AND2X2 AND2X2_75 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_752_) );
OAI21X1 OAI21X1_194 ( .A(_751_), .B(_752_), .C(_65__1_), .Y(_753_) );
NAND2X1 NAND2X1_195 ( .A(_753_), .B(_757_), .Y(_63__1_) );
OAI21X1 OAI21X1_195 ( .A(_754_), .B(_751_), .C(_756_), .Y(_65__2_) );
INVX1 INVX1_120 ( .A(_65__2_), .Y(_761_) );
OR2X2 OR2X2_76 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_762_) );
NAND2X1 NAND2X1_196 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_763_) );
NAND3X1 NAND3X1_76 ( .A(_761_), .B(_763_), .C(_762_), .Y(_764_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_758_) );
AND2X2 AND2X2_76 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_759_) );
OAI21X1 OAI21X1_196 ( .A(_758_), .B(_759_), .C(_65__2_), .Y(_760_) );
NAND2X1 NAND2X1_197 ( .A(_760_), .B(_764_), .Y(_63__2_) );
OAI21X1 OAI21X1_197 ( .A(_761_), .B(_758_), .C(_763_), .Y(_65__3_) );
INVX1 INVX1_121 ( .A(vdd), .Y(_768_) );
OR2X2 OR2X2_77 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_769_) );
NAND2X1 NAND2X1_198 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_770_) );
NAND3X1 NAND3X1_77 ( .A(_768_), .B(_770_), .C(_769_), .Y(_771_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_765_) );
AND2X2 AND2X2_77 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_766_) );
OAI21X1 OAI21X1_198 ( .A(_765_), .B(_766_), .C(vdd), .Y(_767_) );
NAND2X1 NAND2X1_199 ( .A(_767_), .B(_771_), .Y(_64__0_) );
OAI21X1 OAI21X1_199 ( .A(_768_), .B(_765_), .C(_770_), .Y(_66__1_) );
INVX1 INVX1_122 ( .A(_66__3_), .Y(_775_) );
OR2X2 OR2X2_78 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_776_) );
NAND2X1 NAND2X1_200 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_777_) );
NAND3X1 NAND3X1_78 ( .A(_775_), .B(_777_), .C(_776_), .Y(_778_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_772_) );
AND2X2 AND2X2_78 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_773_) );
OAI21X1 OAI21X1_200 ( .A(_772_), .B(_773_), .C(_66__3_), .Y(_774_) );
NAND2X1 NAND2X1_201 ( .A(_774_), .B(_778_), .Y(_64__3_) );
OAI21X1 OAI21X1_201 ( .A(_775_), .B(_772_), .C(_777_), .Y(_62_) );
INVX1 INVX1_123 ( .A(_66__1_), .Y(_782_) );
OR2X2 OR2X2_79 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_783_) );
NAND2X1 NAND2X1_202 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_784_) );
NAND3X1 NAND3X1_79 ( .A(_782_), .B(_784_), .C(_783_), .Y(_785_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_779_) );
AND2X2 AND2X2_79 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_780_) );
OAI21X1 OAI21X1_202 ( .A(_779_), .B(_780_), .C(_66__1_), .Y(_781_) );
NAND2X1 NAND2X1_203 ( .A(_781_), .B(_785_), .Y(_64__1_) );
OAI21X1 OAI21X1_203 ( .A(_782_), .B(_779_), .C(_784_), .Y(_66__2_) );
INVX1 INVX1_124 ( .A(_66__2_), .Y(_789_) );
OR2X2 OR2X2_80 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_790_) );
NAND2X1 NAND2X1_204 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_791_) );
NAND3X1 NAND3X1_80 ( .A(_789_), .B(_791_), .C(_790_), .Y(_792_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_786_) );
AND2X2 AND2X2_80 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_787_) );
OAI21X1 OAI21X1_204 ( .A(_786_), .B(_787_), .C(_66__2_), .Y(_788_) );
NAND2X1 NAND2X1_205 ( .A(_788_), .B(_792_), .Y(_64__2_) );
OAI21X1 OAI21X1_205 ( .A(_789_), .B(_786_), .C(_791_), .Y(_66__3_) );
INVX1 INVX1_125 ( .A(csa_inst_cout0_0), .Y(_793_) );
NAND2X1 NAND2X1_206 ( .A(csa_inst_cout0_1), .B(csa_inst_cin), .Y(_794_) );
OAI21X1 OAI21X1_206 ( .A(csa_inst_cin), .B(_793_), .C(_794_), .Y(w_cout_12_) );
INVX1 INVX1_126 ( .A(gnd), .Y(_796_) );
NAND2X1 NAND2X1_207 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_797_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_795_) );
OAI21X1 OAI21X1_207 ( .A(_796_), .B(_795_), .C(_797_), .Y(csa_inst_rca0_0_fa0_o_carry) );
INVX1 INVX1_127 ( .A(csa_inst_rca0_0_fa31_i_carry), .Y(_799_) );
NAND2X1 NAND2X1_208 ( .A(gnd), .B(gnd), .Y(_800_) );
NOR2X1 NOR2X1_82 ( .A(gnd), .B(gnd), .Y(_798_) );
OAI21X1 OAI21X1_208 ( .A(_799_), .B(_798_), .C(_800_), .Y(csa_inst_cout0_0) );
INVX1 INVX1_128 ( .A(csa_inst_rca0_0_fa0_o_carry), .Y(_802_) );
NAND2X1 NAND2X1_209 ( .A(gnd), .B(gnd), .Y(_803_) );
NOR2X1 NOR2X1_83 ( .A(gnd), .B(gnd), .Y(_801_) );
OAI21X1 OAI21X1_209 ( .A(_802_), .B(_801_), .C(_803_), .Y(csa_inst_rca0_0_fa_1__o_carry) );
INVX1 INVX1_129 ( .A(csa_inst_rca0_0_fa_1__o_carry), .Y(_805_) );
NAND2X1 NAND2X1_210 ( .A(gnd), .B(gnd), .Y(_806_) );
NOR2X1 NOR2X1_84 ( .A(gnd), .B(gnd), .Y(_804_) );
OAI21X1 OAI21X1_210 ( .A(_805_), .B(_804_), .C(_806_), .Y(csa_inst_rca0_0_fa31_i_carry) );
INVX1 INVX1_130 ( .A(vdd), .Y(_808_) );
NAND2X1 NAND2X1_211 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_809_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_807_) );
OAI21X1 OAI21X1_211 ( .A(_808_), .B(_807_), .C(_809_), .Y(csa_inst_rca0_1_fa0_o_carry) );
INVX1 INVX1_131 ( .A(csa_inst_rca0_1_fa31_i_carry), .Y(_811_) );
NAND2X1 NAND2X1_212 ( .A(gnd), .B(gnd), .Y(_812_) );
NOR2X1 NOR2X1_86 ( .A(gnd), .B(gnd), .Y(_810_) );
OAI21X1 OAI21X1_212 ( .A(_811_), .B(_810_), .C(_812_), .Y(csa_inst_cout0_1) );
INVX1 INVX1_132 ( .A(csa_inst_rca0_1_fa0_o_carry), .Y(_814_) );
NAND2X1 NAND2X1_213 ( .A(gnd), .B(gnd), .Y(_815_) );
NOR2X1 NOR2X1_87 ( .A(gnd), .B(gnd), .Y(_813_) );
OAI21X1 OAI21X1_213 ( .A(_814_), .B(_813_), .C(_815_), .Y(csa_inst_rca0_1_fa_1__o_carry) );
INVX1 INVX1_133 ( .A(csa_inst_rca0_1_fa_1__o_carry), .Y(_817_) );
NAND2X1 NAND2X1_214 ( .A(gnd), .B(gnd), .Y(_818_) );
NOR2X1 NOR2X1_88 ( .A(gnd), .B(gnd), .Y(_816_) );
OAI21X1 OAI21X1_214 ( .A(_817_), .B(_816_), .C(_818_), .Y(csa_inst_rca0_1_fa31_i_carry) );
INVX1 INVX1_134 ( .A(gnd), .Y(_822_) );
OR2X2 OR2X2_81 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_823_) );
NAND2X1 NAND2X1_215 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_824_) );
NAND3X1 NAND3X1_81 ( .A(_822_), .B(_824_), .C(_823_), .Y(_825_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_819_) );
AND2X2 AND2X2_81 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_820_) );
OAI21X1 OAI21X1_215 ( .A(_819_), .B(_820_), .C(gnd), .Y(_821_) );
NAND2X1 NAND2X1_216 ( .A(_821_), .B(_825_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_216 ( .A(_822_), .B(_819_), .C(_824_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_135 ( .A(rca_inst_fa31_i_carry), .Y(_829_) );
OR2X2 OR2X2_82 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_830_) );
NAND2X1 NAND2X1_217 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_831_) );
NAND3X1 NAND3X1_82 ( .A(_829_), .B(_831_), .C(_830_), .Y(_832_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_826_) );
AND2X2 AND2X2_82 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_827_) );
OAI21X1 OAI21X1_217 ( .A(_826_), .B(_827_), .C(rca_inst_fa31_i_carry), .Y(_828_) );
NAND2X1 NAND2X1_218 ( .A(_828_), .B(_832_), .Y(rca_inst_fa31_o_sum) );
OAI21X1 OAI21X1_218 ( .A(_829_), .B(_826_), .C(_831_), .Y(rca_inst_cout) );
INVX1 INVX1_136 ( .A(rca_inst_fa0_o_carry), .Y(_836_) );
OR2X2 OR2X2_83 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_837_) );
NAND2X1 NAND2X1_219 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_838_) );
NAND3X1 NAND3X1_83 ( .A(_836_), .B(_838_), .C(_837_), .Y(_839_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_833_) );
AND2X2 AND2X2_83 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_834_) );
OAI21X1 OAI21X1_219 ( .A(_833_), .B(_834_), .C(rca_inst_fa0_o_carry), .Y(_835_) );
NAND2X1 NAND2X1_220 ( .A(_835_), .B(_839_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_220 ( .A(_836_), .B(_833_), .C(_838_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_137 ( .A(rca_inst_fa_1__o_carry), .Y(_843_) );
OR2X2 OR2X2_84 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_844_) );
NAND2X1 NAND2X1_221 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_845_) );
NAND3X1 NAND3X1_84 ( .A(_843_), .B(_845_), .C(_844_), .Y(_846_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_840_) );
AND2X2 AND2X2_84 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_841_) );
OAI21X1 OAI21X1_221 ( .A(_840_), .B(_841_), .C(rca_inst_fa_1__o_carry), .Y(_842_) );
NAND2X1 NAND2X1_222 ( .A(_842_), .B(_846_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_222 ( .A(_843_), .B(_840_), .C(_845_), .Y(rca_inst_fa31_i_carry) );
BUFX2 BUFX2_1 ( .A(w_cout_12_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa31_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(gnd), .Y(sum[48]) );
INVX1 INVX1_138 ( .A(_1_), .Y(_67_) );
NAND2X1 NAND2X1_223 ( .A(_2_), .B(rca_inst_cout), .Y(_68_) );
OAI21X1 OAI21X1_223 ( .A(rca_inst_cout), .B(_67_), .C(_68_), .Y(w_cout_1_) );
INVX1 INVX1_139 ( .A(_3__0_), .Y(_69_) );
NAND2X1 NAND2X1_224 ( .A(_4__0_), .B(rca_inst_cout), .Y(_70_) );
OAI21X1 OAI21X1_224 ( .A(rca_inst_cout), .B(_69_), .C(_70_), .Y(_0__4_) );
INVX1 INVX1_140 ( .A(_3__1_), .Y(_71_) );
NAND2X1 NAND2X1_225 ( .A(rca_inst_cout), .B(_4__1_), .Y(_72_) );
OAI21X1 OAI21X1_225 ( .A(rca_inst_cout), .B(_71_), .C(_72_), .Y(_0__5_) );
INVX1 INVX1_141 ( .A(_3__2_), .Y(_73_) );
NAND2X1 NAND2X1_226 ( .A(rca_inst_cout), .B(_4__2_), .Y(_74_) );
OAI21X1 OAI21X1_226 ( .A(rca_inst_cout), .B(_73_), .C(_74_), .Y(_0__6_) );
INVX1 INVX1_142 ( .A(_3__3_), .Y(_75_) );
NAND2X1 NAND2X1_227 ( .A(rca_inst_cout), .B(_4__3_), .Y(_76_) );
OAI21X1 OAI21X1_227 ( .A(rca_inst_cout), .B(_75_), .C(_76_), .Y(_0__7_) );
INVX1 INVX1_143 ( .A(gnd), .Y(_80_) );
OR2X2 OR2X2_85 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_81_) );
NAND2X1 NAND2X1_228 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_82_) );
NAND3X1 NAND3X1_85 ( .A(_80_), .B(_82_), .C(_81_), .Y(_83_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_77_) );
AND2X2 AND2X2_85 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_78_) );
OAI21X1 OAI21X1_228 ( .A(_77_), .B(_78_), .C(gnd), .Y(_79_) );
NAND2X1 NAND2X1_229 ( .A(_79_), .B(_83_), .Y(_3__0_) );
OAI21X1 OAI21X1_229 ( .A(_80_), .B(_77_), .C(_82_), .Y(_5__1_) );
INVX1 INVX1_144 ( .A(_5__3_), .Y(_87_) );
OR2X2 OR2X2_86 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_88_) );
NAND2X1 NAND2X1_230 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_89_) );
NAND3X1 NAND3X1_86 ( .A(_87_), .B(_89_), .C(_88_), .Y(_90_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_84_) );
AND2X2 AND2X2_86 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_85_) );
OAI21X1 OAI21X1_230 ( .A(_84_), .B(_85_), .C(_5__3_), .Y(_86_) );
NAND2X1 NAND2X1_231 ( .A(_86_), .B(_90_), .Y(_3__3_) );
OAI21X1 OAI21X1_231 ( .A(_87_), .B(_84_), .C(_89_), .Y(_1_) );
INVX1 INVX1_145 ( .A(_5__1_), .Y(_94_) );
OR2X2 OR2X2_87 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_95_) );
NAND2X1 NAND2X1_232 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_96_) );
NAND3X1 NAND3X1_87 ( .A(_94_), .B(_96_), .C(_95_), .Y(_97_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_91_) );
AND2X2 AND2X2_87 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_92_) );
OAI21X1 OAI21X1_232 ( .A(_91_), .B(_92_), .C(_5__1_), .Y(_93_) );
NAND2X1 NAND2X1_233 ( .A(_93_), .B(_97_), .Y(_3__1_) );
OAI21X1 OAI21X1_233 ( .A(_94_), .B(_91_), .C(_96_), .Y(_5__2_) );
INVX1 INVX1_146 ( .A(_5__2_), .Y(_101_) );
OR2X2 OR2X2_88 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_102_) );
NAND2X1 NAND2X1_234 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_103_) );
NAND3X1 NAND3X1_88 ( .A(_101_), .B(_103_), .C(_102_), .Y(_104_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_98_) );
AND2X2 AND2X2_88 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_99_) );
OAI21X1 OAI21X1_234 ( .A(_98_), .B(_99_), .C(_5__2_), .Y(_100_) );
NAND2X1 NAND2X1_235 ( .A(_100_), .B(_104_), .Y(_3__2_) );
OAI21X1 OAI21X1_235 ( .A(_101_), .B(_98_), .C(_103_), .Y(_5__3_) );
INVX1 INVX1_147 ( .A(vdd), .Y(_108_) );
OR2X2 OR2X2_89 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_109_) );
NAND2X1 NAND2X1_236 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_110_) );
NAND3X1 NAND3X1_89 ( .A(_108_), .B(_110_), .C(_109_), .Y(_111_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_105_) );
AND2X2 AND2X2_89 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_106_) );
OAI21X1 OAI21X1_236 ( .A(_105_), .B(_106_), .C(vdd), .Y(_107_) );
NAND2X1 NAND2X1_237 ( .A(_107_), .B(_111_), .Y(_4__0_) );
OAI21X1 OAI21X1_237 ( .A(_108_), .B(_105_), .C(_110_), .Y(_6__1_) );
INVX1 INVX1_148 ( .A(_6__3_), .Y(_115_) );
OR2X2 OR2X2_90 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_116_) );
NAND2X1 NAND2X1_238 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_117_) );
NAND3X1 NAND3X1_90 ( .A(_115_), .B(_117_), .C(_116_), .Y(_118_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_112_) );
AND2X2 AND2X2_90 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_113_) );
OAI21X1 OAI21X1_238 ( .A(_112_), .B(_113_), .C(_6__3_), .Y(_114_) );
NAND2X1 NAND2X1_239 ( .A(_114_), .B(_118_), .Y(_4__3_) );
OAI21X1 OAI21X1_239 ( .A(_115_), .B(_112_), .C(_117_), .Y(_2_) );
INVX1 INVX1_149 ( .A(_6__1_), .Y(_122_) );
OR2X2 OR2X2_91 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_123_) );
NAND2X1 NAND2X1_240 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_124_) );
NAND3X1 NAND3X1_91 ( .A(_122_), .B(_124_), .C(_123_), .Y(_125_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_119_) );
AND2X2 AND2X2_91 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_120_) );
OAI21X1 OAI21X1_240 ( .A(_119_), .B(_120_), .C(_6__1_), .Y(_121_) );
NAND2X1 NAND2X1_241 ( .A(_121_), .B(_125_), .Y(_4__1_) );
OAI21X1 OAI21X1_241 ( .A(_122_), .B(_119_), .C(_124_), .Y(_6__2_) );
INVX1 INVX1_150 ( .A(_6__2_), .Y(_129_) );
OR2X2 OR2X2_92 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_130_) );
NAND2X1 NAND2X1_242 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_131_) );
NAND3X1 NAND3X1_92 ( .A(_129_), .B(_131_), .C(_130_), .Y(_132_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_126_) );
AND2X2 AND2X2_92 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_127_) );
OAI21X1 OAI21X1_242 ( .A(_126_), .B(_127_), .C(_6__2_), .Y(_128_) );
NAND2X1 NAND2X1_243 ( .A(_128_), .B(_132_), .Y(_4__2_) );
OAI21X1 OAI21X1_243 ( .A(_129_), .B(_126_), .C(_131_), .Y(_6__3_) );
INVX1 INVX1_151 ( .A(_7_), .Y(_133_) );
NAND2X1 NAND2X1_244 ( .A(_8_), .B(w_cout_1_), .Y(_134_) );
OAI21X1 OAI21X1_244 ( .A(w_cout_1_), .B(_133_), .C(_134_), .Y(w_cout_2_) );
INVX1 INVX1_152 ( .A(_9__0_), .Y(_135_) );
NAND2X1 NAND2X1_245 ( .A(_10__0_), .B(w_cout_1_), .Y(_136_) );
OAI21X1 OAI21X1_245 ( .A(w_cout_1_), .B(_135_), .C(_136_), .Y(_0__8_) );
INVX1 INVX1_153 ( .A(_9__1_), .Y(_137_) );
NAND2X1 NAND2X1_246 ( .A(w_cout_1_), .B(_10__1_), .Y(_138_) );
OAI21X1 OAI21X1_246 ( .A(w_cout_1_), .B(_137_), .C(_138_), .Y(_0__9_) );
INVX1 INVX1_154 ( .A(_9__2_), .Y(_139_) );
NAND2X1 NAND2X1_247 ( .A(w_cout_1_), .B(_10__2_), .Y(_140_) );
OAI21X1 OAI21X1_247 ( .A(w_cout_1_), .B(_139_), .C(_140_), .Y(_0__10_) );
INVX1 INVX1_155 ( .A(_9__3_), .Y(_141_) );
NAND2X1 NAND2X1_248 ( .A(w_cout_1_), .B(_10__3_), .Y(_142_) );
OAI21X1 OAI21X1_248 ( .A(w_cout_1_), .B(_141_), .C(_142_), .Y(_0__11_) );
INVX1 INVX1_156 ( .A(gnd), .Y(_146_) );
BUFX2 BUFX2_51 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_52 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_53 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_54 ( .A(rca_inst_fa31_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_55 ( .A(gnd), .Y(_0__48_) );
BUFX2 BUFX2_56 ( .A(rca_inst_cout), .Y(w_cout_0_) );
BUFX2 BUFX2_57 ( .A(csa_inst_cin), .Y(w_cout_11_) );
endmodule
