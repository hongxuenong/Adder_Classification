module csa_35bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output cout;

NAND3X1 NAND3X1_1 ( .A(_321_), .B(_323_), .C(_322_), .Y(_324_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_318_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_319_) );
OAI21X1 OAI21X1_1 ( .A(_318_), .B(_319_), .C(_23__3_), .Y(_320_) );
NAND2X1 NAND2X1_1 ( .A(_320_), .B(_324_), .Y(_21__3_) );
OAI21X1 OAI21X1_2 ( .A(_321_), .B(_318_), .C(_323_), .Y(_19_) );
INVX1 INVX1_1 ( .A(1'b1), .Y(_328_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_329_) );
NAND2X1 NAND2X1_2 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_330_) );
NAND3X1 NAND3X1_2 ( .A(_328_), .B(_330_), .C(_329_), .Y(_331_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_325_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_326_) );
OAI21X1 OAI21X1_3 ( .A(_325_), .B(_326_), .C(1'b1), .Y(_327_) );
NAND2X1 NAND2X1_3 ( .A(_327_), .B(_331_), .Y(_22__0_) );
OAI21X1 OAI21X1_4 ( .A(_328_), .B(_325_), .C(_330_), .Y(_24__1_) );
INVX1 INVX1_2 ( .A(_24__1_), .Y(_335_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_336_) );
NAND2X1 NAND2X1_4 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_337_) );
NAND3X1 NAND3X1_3 ( .A(_335_), .B(_337_), .C(_336_), .Y(_338_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_332_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_333_) );
OAI21X1 OAI21X1_5 ( .A(_332_), .B(_333_), .C(_24__1_), .Y(_334_) );
NAND2X1 NAND2X1_5 ( .A(_334_), .B(_338_), .Y(_22__1_) );
OAI21X1 OAI21X1_6 ( .A(_335_), .B(_332_), .C(_337_), .Y(_24__2_) );
INVX1 INVX1_3 ( .A(_24__2_), .Y(_342_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_343_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_344_) );
NAND3X1 NAND3X1_4 ( .A(_342_), .B(_344_), .C(_343_), .Y(_345_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_339_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_340_) );
OAI21X1 OAI21X1_7 ( .A(_339_), .B(_340_), .C(_24__2_), .Y(_341_) );
NAND2X1 NAND2X1_7 ( .A(_341_), .B(_345_), .Y(_22__2_) );
OAI21X1 OAI21X1_8 ( .A(_342_), .B(_339_), .C(_344_), .Y(_24__3_) );
INVX1 INVX1_4 ( .A(_24__3_), .Y(_349_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_350_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_351_) );
NAND3X1 NAND3X1_5 ( .A(_349_), .B(_351_), .C(_350_), .Y(_352_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_346_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_347_) );
OAI21X1 OAI21X1_9 ( .A(_346_), .B(_347_), .C(_24__3_), .Y(_348_) );
NAND2X1 NAND2X1_9 ( .A(_348_), .B(_352_), .Y(_22__3_) );
OAI21X1 OAI21X1_10 ( .A(_349_), .B(_346_), .C(_351_), .Y(_20_) );
INVX1 INVX1_5 ( .A(1'b0), .Y(_356_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_357_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_358_) );
NAND3X1 NAND3X1_6 ( .A(_356_), .B(_358_), .C(_357_), .Y(_359_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_353_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_354_) );
OAI21X1 OAI21X1_11 ( .A(_353_), .B(_354_), .C(1'b0), .Y(_355_) );
NAND2X1 NAND2X1_11 ( .A(_355_), .B(_359_), .Y(_27__0_) );
OAI21X1 OAI21X1_12 ( .A(_356_), .B(_353_), .C(_358_), .Y(_29__1_) );
INVX1 INVX1_6 ( .A(_29__1_), .Y(_363_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_364_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_365_) );
NAND3X1 NAND3X1_7 ( .A(_363_), .B(_365_), .C(_364_), .Y(_366_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_360_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_361_) );
OAI21X1 OAI21X1_13 ( .A(_360_), .B(_361_), .C(_29__1_), .Y(_362_) );
NAND2X1 NAND2X1_13 ( .A(_362_), .B(_366_), .Y(_27__1_) );
OAI21X1 OAI21X1_14 ( .A(_363_), .B(_360_), .C(_365_), .Y(_29__2_) );
INVX1 INVX1_7 ( .A(_29__2_), .Y(_370_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_371_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_372_) );
NAND3X1 NAND3X1_8 ( .A(_370_), .B(_372_), .C(_371_), .Y(_373_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_367_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_368_) );
OAI21X1 OAI21X1_15 ( .A(_367_), .B(_368_), .C(_29__2_), .Y(_369_) );
NAND2X1 NAND2X1_15 ( .A(_369_), .B(_373_), .Y(_27__2_) );
OAI21X1 OAI21X1_16 ( .A(_370_), .B(_367_), .C(_372_), .Y(_29__3_) );
INVX1 INVX1_8 ( .A(_29__3_), .Y(_377_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_378_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_379_) );
NAND3X1 NAND3X1_9 ( .A(_377_), .B(_379_), .C(_378_), .Y(_380_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_374_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_375_) );
OAI21X1 OAI21X1_17 ( .A(_374_), .B(_375_), .C(_29__3_), .Y(_376_) );
NAND2X1 NAND2X1_17 ( .A(_376_), .B(_380_), .Y(_27__3_) );
OAI21X1 OAI21X1_18 ( .A(_377_), .B(_374_), .C(_379_), .Y(_25_) );
INVX1 INVX1_9 ( .A(1'b1), .Y(_384_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_385_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_386_) );
NAND3X1 NAND3X1_10 ( .A(_384_), .B(_386_), .C(_385_), .Y(_387_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_381_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_382_) );
OAI21X1 OAI21X1_19 ( .A(_381_), .B(_382_), .C(1'b1), .Y(_383_) );
NAND2X1 NAND2X1_19 ( .A(_383_), .B(_387_), .Y(_28__0_) );
OAI21X1 OAI21X1_20 ( .A(_384_), .B(_381_), .C(_386_), .Y(_30__1_) );
INVX1 INVX1_10 ( .A(_30__1_), .Y(_391_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_392_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_393_) );
NAND3X1 NAND3X1_11 ( .A(_391_), .B(_393_), .C(_392_), .Y(_394_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_388_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_389_) );
OAI21X1 OAI21X1_21 ( .A(_388_), .B(_389_), .C(_30__1_), .Y(_390_) );
NAND2X1 NAND2X1_21 ( .A(_390_), .B(_394_), .Y(_28__1_) );
OAI21X1 OAI21X1_22 ( .A(_391_), .B(_388_), .C(_393_), .Y(_30__2_) );
INVX1 INVX1_11 ( .A(_30__2_), .Y(_398_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_399_) );
NAND2X1 NAND2X1_22 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_400_) );
NAND3X1 NAND3X1_12 ( .A(_398_), .B(_400_), .C(_399_), .Y(_401_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_395_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_396_) );
OAI21X1 OAI21X1_23 ( .A(_395_), .B(_396_), .C(_30__2_), .Y(_397_) );
NAND2X1 NAND2X1_23 ( .A(_397_), .B(_401_), .Y(_28__2_) );
OAI21X1 OAI21X1_24 ( .A(_398_), .B(_395_), .C(_400_), .Y(_30__3_) );
INVX1 INVX1_12 ( .A(_30__3_), .Y(_405_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_406_) );
NAND2X1 NAND2X1_24 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_407_) );
NAND3X1 NAND3X1_13 ( .A(_405_), .B(_407_), .C(_406_), .Y(_408_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_402_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_403_) );
OAI21X1 OAI21X1_25 ( .A(_402_), .B(_403_), .C(_30__3_), .Y(_404_) );
NAND2X1 NAND2X1_25 ( .A(_404_), .B(_408_), .Y(_28__3_) );
OAI21X1 OAI21X1_26 ( .A(_405_), .B(_402_), .C(_407_), .Y(_26_) );
INVX1 INVX1_13 ( .A(1'b0), .Y(_412_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_413_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_414_) );
NAND3X1 NAND3X1_14 ( .A(_412_), .B(_414_), .C(_413_), .Y(_415_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_409_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_410_) );
OAI21X1 OAI21X1_27 ( .A(_409_), .B(_410_), .C(1'b0), .Y(_411_) );
NAND2X1 NAND2X1_27 ( .A(_411_), .B(_415_), .Y(_33__0_) );
OAI21X1 OAI21X1_28 ( .A(_412_), .B(_409_), .C(_414_), .Y(_35__1_) );
INVX1 INVX1_14 ( .A(_35__1_), .Y(_419_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_420_) );
NAND2X1 NAND2X1_28 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_421_) );
NAND3X1 NAND3X1_15 ( .A(_419_), .B(_421_), .C(_420_), .Y(_422_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_416_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_417_) );
OAI21X1 OAI21X1_29 ( .A(_416_), .B(_417_), .C(_35__1_), .Y(_418_) );
NAND2X1 NAND2X1_29 ( .A(_418_), .B(_422_), .Y(_33__1_) );
OAI21X1 OAI21X1_30 ( .A(_419_), .B(_416_), .C(_421_), .Y(_35__2_) );
INVX1 INVX1_15 ( .A(_35__2_), .Y(_426_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_427_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_428_) );
NAND3X1 NAND3X1_16 ( .A(_426_), .B(_428_), .C(_427_), .Y(_429_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_423_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_424_) );
OAI21X1 OAI21X1_31 ( .A(_423_), .B(_424_), .C(_35__2_), .Y(_425_) );
NAND2X1 NAND2X1_31 ( .A(_425_), .B(_429_), .Y(_33__2_) );
OAI21X1 OAI21X1_32 ( .A(_426_), .B(_423_), .C(_428_), .Y(_35__3_) );
INVX1 INVX1_16 ( .A(_35__3_), .Y(_433_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_434_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_435_) );
NAND3X1 NAND3X1_17 ( .A(_433_), .B(_435_), .C(_434_), .Y(_436_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_430_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_431_) );
OAI21X1 OAI21X1_33 ( .A(_430_), .B(_431_), .C(_35__3_), .Y(_432_) );
NAND2X1 NAND2X1_33 ( .A(_432_), .B(_436_), .Y(_33__3_) );
OAI21X1 OAI21X1_34 ( .A(_433_), .B(_430_), .C(_435_), .Y(_31_) );
INVX1 INVX1_17 ( .A(1'b1), .Y(_440_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_441_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_442_) );
NAND3X1 NAND3X1_18 ( .A(_440_), .B(_442_), .C(_441_), .Y(_443_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_437_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_438_) );
OAI21X1 OAI21X1_35 ( .A(_437_), .B(_438_), .C(1'b1), .Y(_439_) );
NAND2X1 NAND2X1_35 ( .A(_439_), .B(_443_), .Y(_34__0_) );
OAI21X1 OAI21X1_36 ( .A(_440_), .B(_437_), .C(_442_), .Y(_36__1_) );
INVX1 INVX1_18 ( .A(_36__1_), .Y(_447_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_448_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_449_) );
NAND3X1 NAND3X1_19 ( .A(_447_), .B(_449_), .C(_448_), .Y(_450_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_444_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_445_) );
OAI21X1 OAI21X1_37 ( .A(_444_), .B(_445_), .C(_36__1_), .Y(_446_) );
NAND2X1 NAND2X1_37 ( .A(_446_), .B(_450_), .Y(_34__1_) );
OAI21X1 OAI21X1_38 ( .A(_447_), .B(_444_), .C(_449_), .Y(_36__2_) );
INVX1 INVX1_19 ( .A(_36__2_), .Y(_454_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_455_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_456_) );
NAND3X1 NAND3X1_20 ( .A(_454_), .B(_456_), .C(_455_), .Y(_457_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_451_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_452_) );
OAI21X1 OAI21X1_39 ( .A(_451_), .B(_452_), .C(_36__2_), .Y(_453_) );
NAND2X1 NAND2X1_39 ( .A(_453_), .B(_457_), .Y(_34__2_) );
OAI21X1 OAI21X1_40 ( .A(_454_), .B(_451_), .C(_456_), .Y(_36__3_) );
INVX1 INVX1_20 ( .A(_36__3_), .Y(_461_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_462_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_463_) );
NAND3X1 NAND3X1_21 ( .A(_461_), .B(_463_), .C(_462_), .Y(_464_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_458_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_459_) );
OAI21X1 OAI21X1_41 ( .A(_458_), .B(_459_), .C(_36__3_), .Y(_460_) );
NAND2X1 NAND2X1_41 ( .A(_460_), .B(_464_), .Y(_34__3_) );
OAI21X1 OAI21X1_42 ( .A(_461_), .B(_458_), .C(_463_), .Y(_32_) );
INVX1 INVX1_21 ( .A(1'b0), .Y(_468_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_469_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_470_) );
NAND3X1 NAND3X1_22 ( .A(_468_), .B(_470_), .C(_469_), .Y(_471_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_465_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_466_) );
OAI21X1 OAI21X1_43 ( .A(_465_), .B(_466_), .C(1'b0), .Y(_467_) );
NAND2X1 NAND2X1_43 ( .A(_467_), .B(_471_), .Y(_39__0_) );
OAI21X1 OAI21X1_44 ( .A(_468_), .B(_465_), .C(_470_), .Y(_41__1_) );
INVX1 INVX1_22 ( .A(_41__1_), .Y(_475_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_476_) );
NAND2X1 NAND2X1_44 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_477_) );
NAND3X1 NAND3X1_23 ( .A(_475_), .B(_477_), .C(_476_), .Y(_478_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_472_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_473_) );
OAI21X1 OAI21X1_45 ( .A(_472_), .B(_473_), .C(_41__1_), .Y(_474_) );
NAND2X1 NAND2X1_45 ( .A(_474_), .B(_478_), .Y(_39__1_) );
OAI21X1 OAI21X1_46 ( .A(_475_), .B(_472_), .C(_477_), .Y(_41__2_) );
INVX1 INVX1_23 ( .A(_41__2_), .Y(_482_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_483_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_484_) );
NAND3X1 NAND3X1_24 ( .A(_482_), .B(_484_), .C(_483_), .Y(_485_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_479_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_480_) );
OAI21X1 OAI21X1_47 ( .A(_479_), .B(_480_), .C(_41__2_), .Y(_481_) );
NAND2X1 NAND2X1_47 ( .A(_481_), .B(_485_), .Y(_39__2_) );
OAI21X1 OAI21X1_48 ( .A(_482_), .B(_479_), .C(_484_), .Y(_41__3_) );
INVX1 INVX1_24 ( .A(_41__3_), .Y(_489_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_490_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_491_) );
NAND3X1 NAND3X1_25 ( .A(_489_), .B(_491_), .C(_490_), .Y(_492_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_486_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_487_) );
OAI21X1 OAI21X1_49 ( .A(_486_), .B(_487_), .C(_41__3_), .Y(_488_) );
NAND2X1 NAND2X1_49 ( .A(_488_), .B(_492_), .Y(_39__3_) );
OAI21X1 OAI21X1_50 ( .A(_489_), .B(_486_), .C(_491_), .Y(_37_) );
INVX1 INVX1_25 ( .A(1'b1), .Y(_496_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_497_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_498_) );
NAND3X1 NAND3X1_26 ( .A(_496_), .B(_498_), .C(_497_), .Y(_499_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_493_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_494_) );
OAI21X1 OAI21X1_51 ( .A(_493_), .B(_494_), .C(1'b1), .Y(_495_) );
NAND2X1 NAND2X1_51 ( .A(_495_), .B(_499_), .Y(_40__0_) );
OAI21X1 OAI21X1_52 ( .A(_496_), .B(_493_), .C(_498_), .Y(_42__1_) );
INVX1 INVX1_26 ( .A(_42__1_), .Y(_503_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_504_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_505_) );
NAND3X1 NAND3X1_27 ( .A(_503_), .B(_505_), .C(_504_), .Y(_506_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_500_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_501_) );
OAI21X1 OAI21X1_53 ( .A(_500_), .B(_501_), .C(_42__1_), .Y(_502_) );
NAND2X1 NAND2X1_53 ( .A(_502_), .B(_506_), .Y(_40__1_) );
OAI21X1 OAI21X1_54 ( .A(_503_), .B(_500_), .C(_505_), .Y(_42__2_) );
INVX1 INVX1_27 ( .A(_42__2_), .Y(_510_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_511_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_512_) );
NAND3X1 NAND3X1_28 ( .A(_510_), .B(_512_), .C(_511_), .Y(_513_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_507_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_508_) );
OAI21X1 OAI21X1_55 ( .A(_507_), .B(_508_), .C(_42__2_), .Y(_509_) );
NAND2X1 NAND2X1_55 ( .A(_509_), .B(_513_), .Y(_40__2_) );
OAI21X1 OAI21X1_56 ( .A(_510_), .B(_507_), .C(_512_), .Y(_42__3_) );
INVX1 INVX1_28 ( .A(_42__3_), .Y(_517_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_518_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_519_) );
NAND3X1 NAND3X1_29 ( .A(_517_), .B(_519_), .C(_518_), .Y(_520_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_514_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_515_) );
OAI21X1 OAI21X1_57 ( .A(_514_), .B(_515_), .C(_42__3_), .Y(_516_) );
NAND2X1 NAND2X1_57 ( .A(_516_), .B(_520_), .Y(_40__3_) );
OAI21X1 OAI21X1_58 ( .A(_517_), .B(_514_), .C(_519_), .Y(_38_) );
INVX1 INVX1_29 ( .A(1'b0), .Y(_524_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_525_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_526_) );
NAND3X1 NAND3X1_30 ( .A(_524_), .B(_526_), .C(_525_), .Y(_527_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_521_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_522_) );
OAI21X1 OAI21X1_59 ( .A(_521_), .B(_522_), .C(1'b0), .Y(_523_) );
NAND2X1 NAND2X1_59 ( .A(_523_), .B(_527_), .Y(_45__0_) );
OAI21X1 OAI21X1_60 ( .A(_524_), .B(_521_), .C(_526_), .Y(_47__1_) );
INVX1 INVX1_30 ( .A(_47__1_), .Y(_531_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_532_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_533_) );
NAND3X1 NAND3X1_31 ( .A(_531_), .B(_533_), .C(_532_), .Y(_534_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_528_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_529_) );
OAI21X1 OAI21X1_61 ( .A(_528_), .B(_529_), .C(_47__1_), .Y(_530_) );
NAND2X1 NAND2X1_61 ( .A(_530_), .B(_534_), .Y(_45__1_) );
OAI21X1 OAI21X1_62 ( .A(_531_), .B(_528_), .C(_533_), .Y(_47__2_) );
INVX1 INVX1_31 ( .A(_47__2_), .Y(_538_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_539_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_540_) );
NAND3X1 NAND3X1_32 ( .A(_538_), .B(_540_), .C(_539_), .Y(_541_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_535_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_536_) );
OAI21X1 OAI21X1_63 ( .A(_535_), .B(_536_), .C(_47__2_), .Y(_537_) );
NAND2X1 NAND2X1_63 ( .A(_537_), .B(_541_), .Y(_45__2_) );
OAI21X1 OAI21X1_64 ( .A(_538_), .B(_535_), .C(_540_), .Y(_47__3_) );
INVX1 INVX1_32 ( .A(_47__3_), .Y(_545_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_546_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_547_) );
NAND3X1 NAND3X1_33 ( .A(_545_), .B(_547_), .C(_546_), .Y(_548_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_542_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_543_) );
OAI21X1 OAI21X1_65 ( .A(_542_), .B(_543_), .C(_47__3_), .Y(_544_) );
NAND2X1 NAND2X1_65 ( .A(_544_), .B(_548_), .Y(_45__3_) );
OAI21X1 OAI21X1_66 ( .A(_545_), .B(_542_), .C(_547_), .Y(_43_) );
INVX1 INVX1_33 ( .A(1'b1), .Y(_552_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_553_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_554_) );
NAND3X1 NAND3X1_34 ( .A(_552_), .B(_554_), .C(_553_), .Y(_555_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_549_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_550_) );
OAI21X1 OAI21X1_67 ( .A(_549_), .B(_550_), .C(1'b1), .Y(_551_) );
NAND2X1 NAND2X1_67 ( .A(_551_), .B(_555_), .Y(_46__0_) );
OAI21X1 OAI21X1_68 ( .A(_552_), .B(_549_), .C(_554_), .Y(_48__1_) );
INVX1 INVX1_34 ( .A(_48__1_), .Y(_559_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_560_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_561_) );
NAND3X1 NAND3X1_35 ( .A(_559_), .B(_561_), .C(_560_), .Y(_562_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_556_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_557_) );
OAI21X1 OAI21X1_69 ( .A(_556_), .B(_557_), .C(_48__1_), .Y(_558_) );
NAND2X1 NAND2X1_69 ( .A(_558_), .B(_562_), .Y(_46__1_) );
OAI21X1 OAI21X1_70 ( .A(_559_), .B(_556_), .C(_561_), .Y(_48__2_) );
INVX1 INVX1_35 ( .A(_48__2_), .Y(_566_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_567_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_568_) );
NAND3X1 NAND3X1_36 ( .A(_566_), .B(_568_), .C(_567_), .Y(_569_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_563_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_564_) );
OAI21X1 OAI21X1_71 ( .A(_563_), .B(_564_), .C(_48__2_), .Y(_565_) );
NAND2X1 NAND2X1_71 ( .A(_565_), .B(_569_), .Y(_46__2_) );
OAI21X1 OAI21X1_72 ( .A(_566_), .B(_563_), .C(_568_), .Y(_48__3_) );
INVX1 INVX1_36 ( .A(_48__3_), .Y(_573_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_574_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_575_) );
NAND3X1 NAND3X1_37 ( .A(_573_), .B(_575_), .C(_574_), .Y(_576_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_570_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_571_) );
OAI21X1 OAI21X1_73 ( .A(_570_), .B(_571_), .C(_48__3_), .Y(_572_) );
NAND2X1 NAND2X1_73 ( .A(_572_), .B(_576_), .Y(_46__3_) );
OAI21X1 OAI21X1_74 ( .A(_573_), .B(_570_), .C(_575_), .Y(_44_) );
INVX1 INVX1_37 ( .A(1'b0), .Y(_580_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_581_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_582_) );
NAND3X1 NAND3X1_38 ( .A(_580_), .B(_582_), .C(_581_), .Y(_583_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_577_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_578_) );
OAI21X1 OAI21X1_75 ( .A(_577_), .B(_578_), .C(1'b0), .Y(_579_) );
NAND2X1 NAND2X1_75 ( .A(_579_), .B(_583_), .Y(_0__0_) );
OAI21X1 OAI21X1_76 ( .A(_580_), .B(_577_), .C(_582_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_38 ( .A(rca_inst_w_CARRY_1_), .Y(_587_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_588_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_589_) );
NAND3X1 NAND3X1_39 ( .A(_587_), .B(_589_), .C(_588_), .Y(_590_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_584_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_585_) );
OAI21X1 OAI21X1_77 ( .A(_584_), .B(_585_), .C(rca_inst_w_CARRY_1_), .Y(_586_) );
NAND2X1 NAND2X1_77 ( .A(_586_), .B(_590_), .Y(_0__1_) );
OAI21X1 OAI21X1_78 ( .A(_587_), .B(_584_), .C(_589_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_39 ( .A(rca_inst_w_CARRY_2_), .Y(_594_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_595_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_596_) );
NAND3X1 NAND3X1_40 ( .A(_594_), .B(_596_), .C(_595_), .Y(_597_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_591_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_592_) );
OAI21X1 OAI21X1_79 ( .A(_591_), .B(_592_), .C(rca_inst_w_CARRY_2_), .Y(_593_) );
NAND2X1 NAND2X1_79 ( .A(_593_), .B(_597_), .Y(_0__2_) );
BUFX2 BUFX2_1 ( .A(w_cout_8_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
INVX1 INVX1_40 ( .A(_1_), .Y(_49_) );
NAND2X1 NAND2X1_80 ( .A(_2_), .B(1'b0), .Y(_50_) );
OAI21X1 OAI21X1_80 ( .A(1'b0), .B(_49_), .C(_50_), .Y(w_cout_1_) );
INVX1 INVX1_41 ( .A(_3__0_), .Y(_51_) );
NAND2X1 NAND2X1_81 ( .A(_4__0_), .B(1'b0), .Y(_52_) );
OAI21X1 OAI21X1_81 ( .A(1'b0), .B(_51_), .C(_52_), .Y(_0__3_) );
INVX1 INVX1_42 ( .A(_3__1_), .Y(_53_) );
NAND2X1 NAND2X1_82 ( .A(1'b0), .B(_4__1_), .Y(_54_) );
OAI21X1 OAI21X1_82 ( .A(1'b0), .B(_53_), .C(_54_), .Y(_0__4_) );
INVX1 INVX1_43 ( .A(_3__2_), .Y(_55_) );
NAND2X1 NAND2X1_83 ( .A(1'b0), .B(_4__2_), .Y(_56_) );
OAI21X1 OAI21X1_83 ( .A(1'b0), .B(_55_), .C(_56_), .Y(_0__5_) );
INVX1 INVX1_44 ( .A(_3__3_), .Y(_57_) );
NAND2X1 NAND2X1_84 ( .A(1'b0), .B(_4__3_), .Y(_58_) );
OAI21X1 OAI21X1_84 ( .A(1'b0), .B(_57_), .C(_58_), .Y(_0__6_) );
INVX1 INVX1_45 ( .A(_7_), .Y(_59_) );
NAND2X1 NAND2X1_85 ( .A(_8_), .B(w_cout_1_), .Y(_60_) );
OAI21X1 OAI21X1_85 ( .A(w_cout_1_), .B(_59_), .C(_60_), .Y(w_cout_2_) );
INVX1 INVX1_46 ( .A(_9__0_), .Y(_61_) );
NAND2X1 NAND2X1_86 ( .A(_10__0_), .B(w_cout_1_), .Y(_62_) );
OAI21X1 OAI21X1_86 ( .A(w_cout_1_), .B(_61_), .C(_62_), .Y(_0__7_) );
INVX1 INVX1_47 ( .A(_9__1_), .Y(_63_) );
NAND2X1 NAND2X1_87 ( .A(w_cout_1_), .B(_10__1_), .Y(_64_) );
OAI21X1 OAI21X1_87 ( .A(w_cout_1_), .B(_63_), .C(_64_), .Y(_0__8_) );
INVX1 INVX1_48 ( .A(_9__2_), .Y(_65_) );
NAND2X1 NAND2X1_88 ( .A(w_cout_1_), .B(_10__2_), .Y(_66_) );
OAI21X1 OAI21X1_88 ( .A(w_cout_1_), .B(_65_), .C(_66_), .Y(_0__9_) );
INVX1 INVX1_49 ( .A(_9__3_), .Y(_67_) );
NAND2X1 NAND2X1_89 ( .A(w_cout_1_), .B(_10__3_), .Y(_68_) );
OAI21X1 OAI21X1_89 ( .A(w_cout_1_), .B(_67_), .C(_68_), .Y(_0__10_) );
INVX1 INVX1_50 ( .A(_13_), .Y(_69_) );
NAND2X1 NAND2X1_90 ( .A(_14_), .B(w_cout_2_), .Y(_70_) );
OAI21X1 OAI21X1_90 ( .A(w_cout_2_), .B(_69_), .C(_70_), .Y(w_cout_3_) );
INVX1 INVX1_51 ( .A(_15__0_), .Y(_71_) );
NAND2X1 NAND2X1_91 ( .A(_16__0_), .B(w_cout_2_), .Y(_72_) );
OAI21X1 OAI21X1_91 ( .A(w_cout_2_), .B(_71_), .C(_72_), .Y(_0__11_) );
INVX1 INVX1_52 ( .A(_15__1_), .Y(_73_) );
NAND2X1 NAND2X1_92 ( .A(w_cout_2_), .B(_16__1_), .Y(_74_) );
OAI21X1 OAI21X1_92 ( .A(w_cout_2_), .B(_73_), .C(_74_), .Y(_0__12_) );
INVX1 INVX1_53 ( .A(_15__2_), .Y(_75_) );
NAND2X1 NAND2X1_93 ( .A(w_cout_2_), .B(_16__2_), .Y(_76_) );
OAI21X1 OAI21X1_93 ( .A(w_cout_2_), .B(_75_), .C(_76_), .Y(_0__13_) );
INVX1 INVX1_54 ( .A(_15__3_), .Y(_77_) );
NAND2X1 NAND2X1_94 ( .A(w_cout_2_), .B(_16__3_), .Y(_78_) );
OAI21X1 OAI21X1_94 ( .A(w_cout_2_), .B(_77_), .C(_78_), .Y(_0__14_) );
INVX1 INVX1_55 ( .A(_19_), .Y(_79_) );
NAND2X1 NAND2X1_95 ( .A(_20_), .B(w_cout_3_), .Y(_80_) );
OAI21X1 OAI21X1_95 ( .A(w_cout_3_), .B(_79_), .C(_80_), .Y(w_cout_4_) );
INVX1 INVX1_56 ( .A(_21__0_), .Y(_81_) );
NAND2X1 NAND2X1_96 ( .A(_22__0_), .B(w_cout_3_), .Y(_82_) );
OAI21X1 OAI21X1_96 ( .A(w_cout_3_), .B(_81_), .C(_82_), .Y(_0__15_) );
INVX1 INVX1_57 ( .A(_21__1_), .Y(_83_) );
NAND2X1 NAND2X1_97 ( .A(w_cout_3_), .B(_22__1_), .Y(_84_) );
OAI21X1 OAI21X1_97 ( .A(w_cout_3_), .B(_83_), .C(_84_), .Y(_0__16_) );
INVX1 INVX1_58 ( .A(_21__2_), .Y(_85_) );
NAND2X1 NAND2X1_98 ( .A(w_cout_3_), .B(_22__2_), .Y(_86_) );
OAI21X1 OAI21X1_98 ( .A(w_cout_3_), .B(_85_), .C(_86_), .Y(_0__17_) );
INVX1 INVX1_59 ( .A(_21__3_), .Y(_87_) );
NAND2X1 NAND2X1_99 ( .A(w_cout_3_), .B(_22__3_), .Y(_88_) );
OAI21X1 OAI21X1_99 ( .A(w_cout_3_), .B(_87_), .C(_88_), .Y(_0__18_) );
INVX1 INVX1_60 ( .A(_25_), .Y(_89_) );
NAND2X1 NAND2X1_100 ( .A(_26_), .B(w_cout_4_), .Y(_90_) );
OAI21X1 OAI21X1_100 ( .A(w_cout_4_), .B(_89_), .C(_90_), .Y(w_cout_5_) );
INVX1 INVX1_61 ( .A(_27__0_), .Y(_91_) );
NAND2X1 NAND2X1_101 ( .A(_28__0_), .B(w_cout_4_), .Y(_92_) );
OAI21X1 OAI21X1_101 ( .A(w_cout_4_), .B(_91_), .C(_92_), .Y(_0__19_) );
INVX1 INVX1_62 ( .A(_27__1_), .Y(_93_) );
NAND2X1 NAND2X1_102 ( .A(w_cout_4_), .B(_28__1_), .Y(_94_) );
OAI21X1 OAI21X1_102 ( .A(w_cout_4_), .B(_93_), .C(_94_), .Y(_0__20_) );
INVX1 INVX1_63 ( .A(_27__2_), .Y(_95_) );
NAND2X1 NAND2X1_103 ( .A(w_cout_4_), .B(_28__2_), .Y(_96_) );
OAI21X1 OAI21X1_103 ( .A(w_cout_4_), .B(_95_), .C(_96_), .Y(_0__21_) );
INVX1 INVX1_64 ( .A(_27__3_), .Y(_97_) );
NAND2X1 NAND2X1_104 ( .A(w_cout_4_), .B(_28__3_), .Y(_98_) );
OAI21X1 OAI21X1_104 ( .A(w_cout_4_), .B(_97_), .C(_98_), .Y(_0__22_) );
INVX1 INVX1_65 ( .A(_31_), .Y(_99_) );
NAND2X1 NAND2X1_105 ( .A(_32_), .B(w_cout_5_), .Y(_100_) );
OAI21X1 OAI21X1_105 ( .A(w_cout_5_), .B(_99_), .C(_100_), .Y(w_cout_6_) );
INVX1 INVX1_66 ( .A(_33__0_), .Y(_101_) );
NAND2X1 NAND2X1_106 ( .A(_34__0_), .B(w_cout_5_), .Y(_102_) );
OAI21X1 OAI21X1_106 ( .A(w_cout_5_), .B(_101_), .C(_102_), .Y(_0__23_) );
INVX1 INVX1_67 ( .A(_33__1_), .Y(_103_) );
NAND2X1 NAND2X1_107 ( .A(w_cout_5_), .B(_34__1_), .Y(_104_) );
OAI21X1 OAI21X1_107 ( .A(w_cout_5_), .B(_103_), .C(_104_), .Y(_0__24_) );
INVX1 INVX1_68 ( .A(_33__2_), .Y(_105_) );
NAND2X1 NAND2X1_108 ( .A(w_cout_5_), .B(_34__2_), .Y(_106_) );
OAI21X1 OAI21X1_108 ( .A(w_cout_5_), .B(_105_), .C(_106_), .Y(_0__25_) );
INVX1 INVX1_69 ( .A(_33__3_), .Y(_107_) );
NAND2X1 NAND2X1_109 ( .A(w_cout_5_), .B(_34__3_), .Y(_108_) );
OAI21X1 OAI21X1_109 ( .A(w_cout_5_), .B(_107_), .C(_108_), .Y(_0__26_) );
INVX1 INVX1_70 ( .A(_37_), .Y(_109_) );
NAND2X1 NAND2X1_110 ( .A(_38_), .B(w_cout_6_), .Y(_110_) );
OAI21X1 OAI21X1_110 ( .A(w_cout_6_), .B(_109_), .C(_110_), .Y(w_cout_7_) );
INVX1 INVX1_71 ( .A(_39__0_), .Y(_111_) );
NAND2X1 NAND2X1_111 ( .A(_40__0_), .B(w_cout_6_), .Y(_112_) );
OAI21X1 OAI21X1_111 ( .A(w_cout_6_), .B(_111_), .C(_112_), .Y(_0__27_) );
INVX1 INVX1_72 ( .A(_39__1_), .Y(_113_) );
NAND2X1 NAND2X1_112 ( .A(w_cout_6_), .B(_40__1_), .Y(_114_) );
OAI21X1 OAI21X1_112 ( .A(w_cout_6_), .B(_113_), .C(_114_), .Y(_0__28_) );
INVX1 INVX1_73 ( .A(_39__2_), .Y(_115_) );
NAND2X1 NAND2X1_113 ( .A(w_cout_6_), .B(_40__2_), .Y(_116_) );
OAI21X1 OAI21X1_113 ( .A(w_cout_6_), .B(_115_), .C(_116_), .Y(_0__29_) );
INVX1 INVX1_74 ( .A(_39__3_), .Y(_117_) );
NAND2X1 NAND2X1_114 ( .A(w_cout_6_), .B(_40__3_), .Y(_118_) );
OAI21X1 OAI21X1_114 ( .A(w_cout_6_), .B(_117_), .C(_118_), .Y(_0__30_) );
INVX1 INVX1_75 ( .A(_43_), .Y(_119_) );
NAND2X1 NAND2X1_115 ( .A(_44_), .B(w_cout_7_), .Y(_120_) );
OAI21X1 OAI21X1_115 ( .A(w_cout_7_), .B(_119_), .C(_120_), .Y(w_cout_8_) );
INVX1 INVX1_76 ( .A(_45__0_), .Y(_121_) );
NAND2X1 NAND2X1_116 ( .A(_46__0_), .B(w_cout_7_), .Y(_122_) );
OAI21X1 OAI21X1_116 ( .A(w_cout_7_), .B(_121_), .C(_122_), .Y(_0__31_) );
INVX1 INVX1_77 ( .A(_45__1_), .Y(_123_) );
NAND2X1 NAND2X1_117 ( .A(w_cout_7_), .B(_46__1_), .Y(_124_) );
OAI21X1 OAI21X1_117 ( .A(w_cout_7_), .B(_123_), .C(_124_), .Y(_0__32_) );
INVX1 INVX1_78 ( .A(_45__2_), .Y(_125_) );
NAND2X1 NAND2X1_118 ( .A(w_cout_7_), .B(_46__2_), .Y(_126_) );
OAI21X1 OAI21X1_118 ( .A(w_cout_7_), .B(_125_), .C(_126_), .Y(_0__33_) );
INVX1 INVX1_79 ( .A(_45__3_), .Y(_127_) );
NAND2X1 NAND2X1_119 ( .A(w_cout_7_), .B(_46__3_), .Y(_128_) );
OAI21X1 OAI21X1_119 ( .A(w_cout_7_), .B(_127_), .C(_128_), .Y(_0__34_) );
INVX1 INVX1_80 ( .A(1'b0), .Y(_132_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_133_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_134_) );
NAND3X1 NAND3X1_41 ( .A(_132_), .B(_134_), .C(_133_), .Y(_135_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_129_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_130_) );
OAI21X1 OAI21X1_120 ( .A(_129_), .B(_130_), .C(1'b0), .Y(_131_) );
NAND2X1 NAND2X1_121 ( .A(_131_), .B(_135_), .Y(_3__0_) );
OAI21X1 OAI21X1_121 ( .A(_132_), .B(_129_), .C(_134_), .Y(_5__1_) );
INVX1 INVX1_81 ( .A(_5__1_), .Y(_139_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_140_) );
NAND2X1 NAND2X1_122 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_141_) );
NAND3X1 NAND3X1_42 ( .A(_139_), .B(_141_), .C(_140_), .Y(_142_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_136_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_137_) );
OAI21X1 OAI21X1_122 ( .A(_136_), .B(_137_), .C(_5__1_), .Y(_138_) );
NAND2X1 NAND2X1_123 ( .A(_138_), .B(_142_), .Y(_3__1_) );
OAI21X1 OAI21X1_123 ( .A(_139_), .B(_136_), .C(_141_), .Y(_5__2_) );
INVX1 INVX1_82 ( .A(_5__2_), .Y(_146_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_147_) );
NAND2X1 NAND2X1_124 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_148_) );
NAND3X1 NAND3X1_43 ( .A(_146_), .B(_148_), .C(_147_), .Y(_149_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_143_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_144_) );
OAI21X1 OAI21X1_124 ( .A(_143_), .B(_144_), .C(_5__2_), .Y(_145_) );
NAND2X1 NAND2X1_125 ( .A(_145_), .B(_149_), .Y(_3__2_) );
OAI21X1 OAI21X1_125 ( .A(_146_), .B(_143_), .C(_148_), .Y(_5__3_) );
INVX1 INVX1_83 ( .A(_5__3_), .Y(_153_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_154_) );
NAND2X1 NAND2X1_126 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_155_) );
NAND3X1 NAND3X1_44 ( .A(_153_), .B(_155_), .C(_154_), .Y(_156_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_150_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_151_) );
OAI21X1 OAI21X1_126 ( .A(_150_), .B(_151_), .C(_5__3_), .Y(_152_) );
NAND2X1 NAND2X1_127 ( .A(_152_), .B(_156_), .Y(_3__3_) );
OAI21X1 OAI21X1_127 ( .A(_153_), .B(_150_), .C(_155_), .Y(_1_) );
INVX1 INVX1_84 ( .A(1'b1), .Y(_160_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_161_) );
NAND2X1 NAND2X1_128 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_162_) );
NAND3X1 NAND3X1_45 ( .A(_160_), .B(_162_), .C(_161_), .Y(_163_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_157_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_158_) );
OAI21X1 OAI21X1_128 ( .A(_157_), .B(_158_), .C(1'b1), .Y(_159_) );
NAND2X1 NAND2X1_129 ( .A(_159_), .B(_163_), .Y(_4__0_) );
OAI21X1 OAI21X1_129 ( .A(_160_), .B(_157_), .C(_162_), .Y(_6__1_) );
INVX1 INVX1_85 ( .A(_6__1_), .Y(_167_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_168_) );
NAND2X1 NAND2X1_130 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_169_) );
NAND3X1 NAND3X1_46 ( .A(_167_), .B(_169_), .C(_168_), .Y(_170_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_164_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_165_) );
OAI21X1 OAI21X1_130 ( .A(_164_), .B(_165_), .C(_6__1_), .Y(_166_) );
NAND2X1 NAND2X1_131 ( .A(_166_), .B(_170_), .Y(_4__1_) );
OAI21X1 OAI21X1_131 ( .A(_167_), .B(_164_), .C(_169_), .Y(_6__2_) );
INVX1 INVX1_86 ( .A(_6__2_), .Y(_174_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_175_) );
NAND2X1 NAND2X1_132 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_176_) );
NAND3X1 NAND3X1_47 ( .A(_174_), .B(_176_), .C(_175_), .Y(_177_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_171_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_172_) );
OAI21X1 OAI21X1_132 ( .A(_171_), .B(_172_), .C(_6__2_), .Y(_173_) );
NAND2X1 NAND2X1_133 ( .A(_173_), .B(_177_), .Y(_4__2_) );
OAI21X1 OAI21X1_133 ( .A(_174_), .B(_171_), .C(_176_), .Y(_6__3_) );
INVX1 INVX1_87 ( .A(_6__3_), .Y(_181_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_182_) );
NAND2X1 NAND2X1_134 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_183_) );
NAND3X1 NAND3X1_48 ( .A(_181_), .B(_183_), .C(_182_), .Y(_184_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_178_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_179_) );
OAI21X1 OAI21X1_134 ( .A(_178_), .B(_179_), .C(_6__3_), .Y(_180_) );
NAND2X1 NAND2X1_135 ( .A(_180_), .B(_184_), .Y(_4__3_) );
OAI21X1 OAI21X1_135 ( .A(_181_), .B(_178_), .C(_183_), .Y(_2_) );
INVX1 INVX1_88 ( .A(1'b0), .Y(_188_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_189_) );
NAND2X1 NAND2X1_136 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_190_) );
NAND3X1 NAND3X1_49 ( .A(_188_), .B(_190_), .C(_189_), .Y(_191_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_185_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_186_) );
OAI21X1 OAI21X1_136 ( .A(_185_), .B(_186_), .C(1'b0), .Y(_187_) );
NAND2X1 NAND2X1_137 ( .A(_187_), .B(_191_), .Y(_9__0_) );
OAI21X1 OAI21X1_137 ( .A(_188_), .B(_185_), .C(_190_), .Y(_11__1_) );
INVX1 INVX1_89 ( .A(_11__1_), .Y(_195_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_196_) );
NAND2X1 NAND2X1_138 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_197_) );
NAND3X1 NAND3X1_50 ( .A(_195_), .B(_197_), .C(_196_), .Y(_198_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_192_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_193_) );
OAI21X1 OAI21X1_138 ( .A(_192_), .B(_193_), .C(_11__1_), .Y(_194_) );
NAND2X1 NAND2X1_139 ( .A(_194_), .B(_198_), .Y(_9__1_) );
OAI21X1 OAI21X1_139 ( .A(_195_), .B(_192_), .C(_197_), .Y(_11__2_) );
INVX1 INVX1_90 ( .A(_11__2_), .Y(_202_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_203_) );
NAND2X1 NAND2X1_140 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_204_) );
NAND3X1 NAND3X1_51 ( .A(_202_), .B(_204_), .C(_203_), .Y(_205_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_199_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_200_) );
OAI21X1 OAI21X1_140 ( .A(_199_), .B(_200_), .C(_11__2_), .Y(_201_) );
NAND2X1 NAND2X1_141 ( .A(_201_), .B(_205_), .Y(_9__2_) );
OAI21X1 OAI21X1_141 ( .A(_202_), .B(_199_), .C(_204_), .Y(_11__3_) );
INVX1 INVX1_91 ( .A(_11__3_), .Y(_209_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_210_) );
NAND2X1 NAND2X1_142 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_211_) );
NAND3X1 NAND3X1_52 ( .A(_209_), .B(_211_), .C(_210_), .Y(_212_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_206_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_207_) );
OAI21X1 OAI21X1_142 ( .A(_206_), .B(_207_), .C(_11__3_), .Y(_208_) );
NAND2X1 NAND2X1_143 ( .A(_208_), .B(_212_), .Y(_9__3_) );
OAI21X1 OAI21X1_143 ( .A(_209_), .B(_206_), .C(_211_), .Y(_7_) );
INVX1 INVX1_92 ( .A(1'b1), .Y(_216_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_217_) );
NAND2X1 NAND2X1_144 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_218_) );
NAND3X1 NAND3X1_53 ( .A(_216_), .B(_218_), .C(_217_), .Y(_219_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_213_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_214_) );
OAI21X1 OAI21X1_144 ( .A(_213_), .B(_214_), .C(1'b1), .Y(_215_) );
NAND2X1 NAND2X1_145 ( .A(_215_), .B(_219_), .Y(_10__0_) );
OAI21X1 OAI21X1_145 ( .A(_216_), .B(_213_), .C(_218_), .Y(_12__1_) );
INVX1 INVX1_93 ( .A(_12__1_), .Y(_223_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_224_) );
NAND2X1 NAND2X1_146 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_225_) );
NAND3X1 NAND3X1_54 ( .A(_223_), .B(_225_), .C(_224_), .Y(_226_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_220_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_221_) );
OAI21X1 OAI21X1_146 ( .A(_220_), .B(_221_), .C(_12__1_), .Y(_222_) );
NAND2X1 NAND2X1_147 ( .A(_222_), .B(_226_), .Y(_10__1_) );
OAI21X1 OAI21X1_147 ( .A(_223_), .B(_220_), .C(_225_), .Y(_12__2_) );
INVX1 INVX1_94 ( .A(_12__2_), .Y(_230_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_231_) );
NAND2X1 NAND2X1_148 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_232_) );
NAND3X1 NAND3X1_55 ( .A(_230_), .B(_232_), .C(_231_), .Y(_233_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_227_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_228_) );
OAI21X1 OAI21X1_148 ( .A(_227_), .B(_228_), .C(_12__2_), .Y(_229_) );
NAND2X1 NAND2X1_149 ( .A(_229_), .B(_233_), .Y(_10__2_) );
OAI21X1 OAI21X1_149 ( .A(_230_), .B(_227_), .C(_232_), .Y(_12__3_) );
INVX1 INVX1_95 ( .A(_12__3_), .Y(_237_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_238_) );
NAND2X1 NAND2X1_150 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_239_) );
NAND3X1 NAND3X1_56 ( .A(_237_), .B(_239_), .C(_238_), .Y(_240_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_234_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_235_) );
OAI21X1 OAI21X1_150 ( .A(_234_), .B(_235_), .C(_12__3_), .Y(_236_) );
NAND2X1 NAND2X1_151 ( .A(_236_), .B(_240_), .Y(_10__3_) );
OAI21X1 OAI21X1_151 ( .A(_237_), .B(_234_), .C(_239_), .Y(_8_) );
INVX1 INVX1_96 ( .A(1'b0), .Y(_244_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_245_) );
NAND2X1 NAND2X1_152 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_246_) );
NAND3X1 NAND3X1_57 ( .A(_244_), .B(_246_), .C(_245_), .Y(_247_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_241_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_242_) );
OAI21X1 OAI21X1_152 ( .A(_241_), .B(_242_), .C(1'b0), .Y(_243_) );
NAND2X1 NAND2X1_153 ( .A(_243_), .B(_247_), .Y(_15__0_) );
OAI21X1 OAI21X1_153 ( .A(_244_), .B(_241_), .C(_246_), .Y(_17__1_) );
INVX1 INVX1_97 ( .A(_17__1_), .Y(_251_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_252_) );
NAND2X1 NAND2X1_154 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_253_) );
NAND3X1 NAND3X1_58 ( .A(_251_), .B(_253_), .C(_252_), .Y(_254_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_248_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_249_) );
OAI21X1 OAI21X1_154 ( .A(_248_), .B(_249_), .C(_17__1_), .Y(_250_) );
NAND2X1 NAND2X1_155 ( .A(_250_), .B(_254_), .Y(_15__1_) );
OAI21X1 OAI21X1_155 ( .A(_251_), .B(_248_), .C(_253_), .Y(_17__2_) );
INVX1 INVX1_98 ( .A(_17__2_), .Y(_258_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_259_) );
NAND2X1 NAND2X1_156 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_260_) );
NAND3X1 NAND3X1_59 ( .A(_258_), .B(_260_), .C(_259_), .Y(_261_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_255_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_256_) );
OAI21X1 OAI21X1_156 ( .A(_255_), .B(_256_), .C(_17__2_), .Y(_257_) );
NAND2X1 NAND2X1_157 ( .A(_257_), .B(_261_), .Y(_15__2_) );
OAI21X1 OAI21X1_157 ( .A(_258_), .B(_255_), .C(_260_), .Y(_17__3_) );
INVX1 INVX1_99 ( .A(_17__3_), .Y(_265_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_266_) );
NAND2X1 NAND2X1_158 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_267_) );
NAND3X1 NAND3X1_60 ( .A(_265_), .B(_267_), .C(_266_), .Y(_268_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_262_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_263_) );
OAI21X1 OAI21X1_158 ( .A(_262_), .B(_263_), .C(_17__3_), .Y(_264_) );
NAND2X1 NAND2X1_159 ( .A(_264_), .B(_268_), .Y(_15__3_) );
OAI21X1 OAI21X1_159 ( .A(_265_), .B(_262_), .C(_267_), .Y(_13_) );
INVX1 INVX1_100 ( .A(1'b1), .Y(_272_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_273_) );
NAND2X1 NAND2X1_160 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_274_) );
NAND3X1 NAND3X1_61 ( .A(_272_), .B(_274_), .C(_273_), .Y(_275_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_269_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_270_) );
OAI21X1 OAI21X1_160 ( .A(_269_), .B(_270_), .C(1'b1), .Y(_271_) );
NAND2X1 NAND2X1_161 ( .A(_271_), .B(_275_), .Y(_16__0_) );
OAI21X1 OAI21X1_161 ( .A(_272_), .B(_269_), .C(_274_), .Y(_18__1_) );
INVX1 INVX1_101 ( .A(_18__1_), .Y(_279_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_280_) );
NAND2X1 NAND2X1_162 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_281_) );
NAND3X1 NAND3X1_62 ( .A(_279_), .B(_281_), .C(_280_), .Y(_282_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_276_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_277_) );
OAI21X1 OAI21X1_162 ( .A(_276_), .B(_277_), .C(_18__1_), .Y(_278_) );
NAND2X1 NAND2X1_163 ( .A(_278_), .B(_282_), .Y(_16__1_) );
OAI21X1 OAI21X1_163 ( .A(_279_), .B(_276_), .C(_281_), .Y(_18__2_) );
INVX1 INVX1_102 ( .A(_18__2_), .Y(_286_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_287_) );
NAND2X1 NAND2X1_164 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_288_) );
NAND3X1 NAND3X1_63 ( .A(_286_), .B(_288_), .C(_287_), .Y(_289_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_283_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_284_) );
OAI21X1 OAI21X1_164 ( .A(_283_), .B(_284_), .C(_18__2_), .Y(_285_) );
NAND2X1 NAND2X1_165 ( .A(_285_), .B(_289_), .Y(_16__2_) );
OAI21X1 OAI21X1_165 ( .A(_286_), .B(_283_), .C(_288_), .Y(_18__3_) );
INVX1 INVX1_103 ( .A(_18__3_), .Y(_293_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_294_) );
NAND2X1 NAND2X1_166 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_295_) );
NAND3X1 NAND3X1_64 ( .A(_293_), .B(_295_), .C(_294_), .Y(_296_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_290_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_291_) );
OAI21X1 OAI21X1_166 ( .A(_290_), .B(_291_), .C(_18__3_), .Y(_292_) );
NAND2X1 NAND2X1_167 ( .A(_292_), .B(_296_), .Y(_16__3_) );
OAI21X1 OAI21X1_167 ( .A(_293_), .B(_290_), .C(_295_), .Y(_14_) );
INVX1 INVX1_104 ( .A(1'b0), .Y(_300_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_301_) );
NAND2X1 NAND2X1_168 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_302_) );
NAND3X1 NAND3X1_65 ( .A(_300_), .B(_302_), .C(_301_), .Y(_303_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_297_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_298_) );
OAI21X1 OAI21X1_168 ( .A(_297_), .B(_298_), .C(1'b0), .Y(_299_) );
NAND2X1 NAND2X1_169 ( .A(_299_), .B(_303_), .Y(_21__0_) );
OAI21X1 OAI21X1_169 ( .A(_300_), .B(_297_), .C(_302_), .Y(_23__1_) );
INVX1 INVX1_105 ( .A(_23__1_), .Y(_307_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_308_) );
NAND2X1 NAND2X1_170 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_309_) );
NAND3X1 NAND3X1_66 ( .A(_307_), .B(_309_), .C(_308_), .Y(_310_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_304_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_305_) );
OAI21X1 OAI21X1_170 ( .A(_304_), .B(_305_), .C(_23__1_), .Y(_306_) );
NAND2X1 NAND2X1_171 ( .A(_306_), .B(_310_), .Y(_21__1_) );
OAI21X1 OAI21X1_171 ( .A(_307_), .B(_304_), .C(_309_), .Y(_23__2_) );
INVX1 INVX1_106 ( .A(_23__2_), .Y(_314_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_315_) );
NAND2X1 NAND2X1_172 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_316_) );
NAND3X1 NAND3X1_67 ( .A(_314_), .B(_316_), .C(_315_), .Y(_317_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_311_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_312_) );
OAI21X1 OAI21X1_172 ( .A(_311_), .B(_312_), .C(_23__2_), .Y(_313_) );
NAND2X1 NAND2X1_173 ( .A(_313_), .B(_317_), .Y(_21__2_) );
OAI21X1 OAI21X1_173 ( .A(_314_), .B(_311_), .C(_316_), .Y(_23__3_) );
INVX1 INVX1_107 ( .A(_23__3_), .Y(_321_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_322_) );
NAND2X1 NAND2X1_174 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_323_) );
BUFX2 BUFX2_37 ( .A(1'b0), .Y(_5__0_) );
BUFX2 BUFX2_38 ( .A(_1_), .Y(_5__4_) );
BUFX2 BUFX2_39 ( .A(1'b1), .Y(_6__0_) );
BUFX2 BUFX2_40 ( .A(_2_), .Y(_6__4_) );
BUFX2 BUFX2_41 ( .A(1'b0), .Y(_11__0_) );
BUFX2 BUFX2_42 ( .A(_7_), .Y(_11__4_) );
BUFX2 BUFX2_43 ( .A(1'b1), .Y(_12__0_) );
BUFX2 BUFX2_44 ( .A(_8_), .Y(_12__4_) );
BUFX2 BUFX2_45 ( .A(1'b0), .Y(_17__0_) );
BUFX2 BUFX2_46 ( .A(_13_), .Y(_17__4_) );
BUFX2 BUFX2_47 ( .A(1'b1), .Y(_18__0_) );
BUFX2 BUFX2_48 ( .A(_14_), .Y(_18__4_) );
BUFX2 BUFX2_49 ( .A(1'b0), .Y(_23__0_) );
BUFX2 BUFX2_50 ( .A(_19_), .Y(_23__4_) );
BUFX2 BUFX2_51 ( .A(1'b1), .Y(_24__0_) );
BUFX2 BUFX2_52 ( .A(_20_), .Y(_24__4_) );
BUFX2 BUFX2_53 ( .A(1'b0), .Y(_29__0_) );
BUFX2 BUFX2_54 ( .A(_25_), .Y(_29__4_) );
BUFX2 BUFX2_55 ( .A(1'b1), .Y(_30__0_) );
BUFX2 BUFX2_56 ( .A(_26_), .Y(_30__4_) );
BUFX2 BUFX2_57 ( .A(1'b0), .Y(_35__0_) );
BUFX2 BUFX2_58 ( .A(_31_), .Y(_35__4_) );
BUFX2 BUFX2_59 ( .A(1'b1), .Y(_36__0_) );
BUFX2 BUFX2_60 ( .A(_32_), .Y(_36__4_) );
BUFX2 BUFX2_61 ( .A(1'b0), .Y(_41__0_) );
BUFX2 BUFX2_62 ( .A(_37_), .Y(_41__4_) );
BUFX2 BUFX2_63 ( .A(1'b1), .Y(_42__0_) );
BUFX2 BUFX2_64 ( .A(_38_), .Y(_42__4_) );
BUFX2 BUFX2_65 ( .A(1'b0), .Y(_47__0_) );
BUFX2 BUFX2_66 ( .A(_43_), .Y(_47__4_) );
BUFX2 BUFX2_67 ( .A(1'b1), .Y(_48__0_) );
BUFX2 BUFX2_68 ( .A(_44_), .Y(_48__4_) );
BUFX2 BUFX2_69 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_70 ( .A(1'b0), .Y(w_cout_0_) );
endmodule
