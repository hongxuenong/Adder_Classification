module csa_55bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term1[45], i_add_term1[46], i_add_term1[47], i_add_term1[48], i_add_term1[49], i_add_term1[50], i_add_term1[51], i_add_term1[52], i_add_term1[53], i_add_term1[54], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], i_add_term2[45], i_add_term2[46], i_add_term2[47], i_add_term2[48], i_add_term2[49], i_add_term2[50], i_add_term2[51], i_add_term2[52], i_add_term2[53], i_add_term2[54], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], sum[45], sum[46], sum[47], sum[48], sum[49], sum[50], sum[51], sum[52], sum[53], sum[54], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term1[45];
input i_add_term1[46];
input i_add_term1[47];
input i_add_term1[48];
input i_add_term1[49];
input i_add_term1[50];
input i_add_term1[51];
input i_add_term1[52];
input i_add_term1[53];
input i_add_term1[54];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
input i_add_term2[45];
input i_add_term2[46];
input i_add_term2[47];
input i_add_term2[48];
input i_add_term2[49];
input i_add_term2[50];
input i_add_term2[51];
input i_add_term2[52];
input i_add_term2[53];
input i_add_term2[54];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output sum[45];
output sum[46];
output sum[47];
output sum[48];
output sum[49];
output sum[50];
output sum[51];
output sum[52];
output sum[53];
output sum[54];
output cout;

BUFX2 BUFX2_1 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_2 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_3 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_4 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_5 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_6 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_7 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_8 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_9 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_10 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_11 ( .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_12 ( .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_13 ( .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_14 ( .A(_0__54_), .Y(sum[54]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_79_) );
NAND2X1 NAND2X1_1 ( .A(_2_), .B(1'b0), .Y(_80_) );
OAI21X1 OAI21X1_1 ( .A(1'b0), .B(_79_), .C(_80_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3__0_), .Y(_81_) );
NAND2X1 NAND2X1_2 ( .A(_4__0_), .B(1'b0), .Y(_82_) );
OAI21X1 OAI21X1_2 ( .A(1'b0), .B(_81_), .C(_82_), .Y(_0__3_) );
INVX1 INVX1_3 ( .A(_3__1_), .Y(_83_) );
NAND2X1 NAND2X1_3 ( .A(1'b0), .B(_4__1_), .Y(_84_) );
OAI21X1 OAI21X1_3 ( .A(1'b0), .B(_83_), .C(_84_), .Y(_0__4_) );
INVX1 INVX1_4 ( .A(_3__2_), .Y(_85_) );
NAND2X1 NAND2X1_4 ( .A(1'b0), .B(_4__2_), .Y(_86_) );
OAI21X1 OAI21X1_4 ( .A(1'b0), .B(_85_), .C(_86_), .Y(_0__5_) );
INVX1 INVX1_5 ( .A(_3__3_), .Y(_87_) );
NAND2X1 NAND2X1_5 ( .A(1'b0), .B(_4__3_), .Y(_88_) );
OAI21X1 OAI21X1_5 ( .A(1'b0), .B(_87_), .C(_88_), .Y(_0__6_) );
INVX1 INVX1_6 ( .A(_7_), .Y(_89_) );
NAND2X1 NAND2X1_6 ( .A(_8_), .B(w_cout_1_), .Y(_90_) );
OAI21X1 OAI21X1_6 ( .A(w_cout_1_), .B(_89_), .C(_90_), .Y(w_cout_2_) );
INVX1 INVX1_7 ( .A(_9__0_), .Y(_91_) );
NAND2X1 NAND2X1_7 ( .A(_10__0_), .B(w_cout_1_), .Y(_92_) );
OAI21X1 OAI21X1_7 ( .A(w_cout_1_), .B(_91_), .C(_92_), .Y(_0__7_) );
INVX1 INVX1_8 ( .A(_9__1_), .Y(_93_) );
NAND2X1 NAND2X1_8 ( .A(w_cout_1_), .B(_10__1_), .Y(_94_) );
OAI21X1 OAI21X1_8 ( .A(w_cout_1_), .B(_93_), .C(_94_), .Y(_0__8_) );
INVX1 INVX1_9 ( .A(_9__2_), .Y(_95_) );
NAND2X1 NAND2X1_9 ( .A(w_cout_1_), .B(_10__2_), .Y(_96_) );
OAI21X1 OAI21X1_9 ( .A(w_cout_1_), .B(_95_), .C(_96_), .Y(_0__9_) );
INVX1 INVX1_10 ( .A(_9__3_), .Y(_97_) );
NAND2X1 NAND2X1_10 ( .A(w_cout_1_), .B(_10__3_), .Y(_98_) );
OAI21X1 OAI21X1_10 ( .A(w_cout_1_), .B(_97_), .C(_98_), .Y(_0__10_) );
INVX1 INVX1_11 ( .A(_13_), .Y(_99_) );
NAND2X1 NAND2X1_11 ( .A(_14_), .B(w_cout_2_), .Y(_100_) );
OAI21X1 OAI21X1_11 ( .A(w_cout_2_), .B(_99_), .C(_100_), .Y(w_cout_3_) );
INVX1 INVX1_12 ( .A(_15__0_), .Y(_101_) );
NAND2X1 NAND2X1_12 ( .A(_16__0_), .B(w_cout_2_), .Y(_102_) );
OAI21X1 OAI21X1_12 ( .A(w_cout_2_), .B(_101_), .C(_102_), .Y(_0__11_) );
INVX1 INVX1_13 ( .A(_15__1_), .Y(_103_) );
NAND2X1 NAND2X1_13 ( .A(w_cout_2_), .B(_16__1_), .Y(_104_) );
OAI21X1 OAI21X1_13 ( .A(w_cout_2_), .B(_103_), .C(_104_), .Y(_0__12_) );
INVX1 INVX1_14 ( .A(_15__2_), .Y(_105_) );
NAND2X1 NAND2X1_14 ( .A(w_cout_2_), .B(_16__2_), .Y(_106_) );
OAI21X1 OAI21X1_14 ( .A(w_cout_2_), .B(_105_), .C(_106_), .Y(_0__13_) );
INVX1 INVX1_15 ( .A(_15__3_), .Y(_107_) );
NAND2X1 NAND2X1_15 ( .A(w_cout_2_), .B(_16__3_), .Y(_108_) );
OAI21X1 OAI21X1_15 ( .A(w_cout_2_), .B(_107_), .C(_108_), .Y(_0__14_) );
INVX1 INVX1_16 ( .A(_19_), .Y(_109_) );
NAND2X1 NAND2X1_16 ( .A(_20_), .B(w_cout_3_), .Y(_110_) );
OAI21X1 OAI21X1_16 ( .A(w_cout_3_), .B(_109_), .C(_110_), .Y(w_cout_4_) );
INVX1 INVX1_17 ( .A(_21__0_), .Y(_111_) );
NAND2X1 NAND2X1_17 ( .A(_22__0_), .B(w_cout_3_), .Y(_112_) );
OAI21X1 OAI21X1_17 ( .A(w_cout_3_), .B(_111_), .C(_112_), .Y(_0__15_) );
INVX1 INVX1_18 ( .A(_21__1_), .Y(_113_) );
NAND2X1 NAND2X1_18 ( .A(w_cout_3_), .B(_22__1_), .Y(_114_) );
OAI21X1 OAI21X1_18 ( .A(w_cout_3_), .B(_113_), .C(_114_), .Y(_0__16_) );
INVX1 INVX1_19 ( .A(_21__2_), .Y(_115_) );
NAND2X1 NAND2X1_19 ( .A(w_cout_3_), .B(_22__2_), .Y(_116_) );
OAI21X1 OAI21X1_19 ( .A(w_cout_3_), .B(_115_), .C(_116_), .Y(_0__17_) );
INVX1 INVX1_20 ( .A(_21__3_), .Y(_117_) );
NAND2X1 NAND2X1_20 ( .A(w_cout_3_), .B(_22__3_), .Y(_118_) );
OAI21X1 OAI21X1_20 ( .A(w_cout_3_), .B(_117_), .C(_118_), .Y(_0__18_) );
INVX1 INVX1_21 ( .A(_25_), .Y(_119_) );
NAND2X1 NAND2X1_21 ( .A(_26_), .B(w_cout_4_), .Y(_120_) );
OAI21X1 OAI21X1_21 ( .A(w_cout_4_), .B(_119_), .C(_120_), .Y(w_cout_5_) );
INVX1 INVX1_22 ( .A(_27__0_), .Y(_121_) );
NAND2X1 NAND2X1_22 ( .A(_28__0_), .B(w_cout_4_), .Y(_122_) );
OAI21X1 OAI21X1_22 ( .A(w_cout_4_), .B(_121_), .C(_122_), .Y(_0__19_) );
INVX1 INVX1_23 ( .A(_27__1_), .Y(_123_) );
NAND2X1 NAND2X1_23 ( .A(w_cout_4_), .B(_28__1_), .Y(_124_) );
OAI21X1 OAI21X1_23 ( .A(w_cout_4_), .B(_123_), .C(_124_), .Y(_0__20_) );
INVX1 INVX1_24 ( .A(_27__2_), .Y(_125_) );
NAND2X1 NAND2X1_24 ( .A(w_cout_4_), .B(_28__2_), .Y(_126_) );
OAI21X1 OAI21X1_24 ( .A(w_cout_4_), .B(_125_), .C(_126_), .Y(_0__21_) );
INVX1 INVX1_25 ( .A(_27__3_), .Y(_127_) );
NAND2X1 NAND2X1_25 ( .A(w_cout_4_), .B(_28__3_), .Y(_128_) );
OAI21X1 OAI21X1_25 ( .A(w_cout_4_), .B(_127_), .C(_128_), .Y(_0__22_) );
INVX1 INVX1_26 ( .A(_31_), .Y(_129_) );
NAND2X1 NAND2X1_26 ( .A(_32_), .B(w_cout_5_), .Y(_130_) );
OAI21X1 OAI21X1_26 ( .A(w_cout_5_), .B(_129_), .C(_130_), .Y(w_cout_6_) );
INVX1 INVX1_27 ( .A(_33__0_), .Y(_131_) );
NAND2X1 NAND2X1_27 ( .A(_34__0_), .B(w_cout_5_), .Y(_132_) );
OAI21X1 OAI21X1_27 ( .A(w_cout_5_), .B(_131_), .C(_132_), .Y(_0__23_) );
INVX1 INVX1_28 ( .A(_33__1_), .Y(_133_) );
NAND2X1 NAND2X1_28 ( .A(w_cout_5_), .B(_34__1_), .Y(_134_) );
OAI21X1 OAI21X1_28 ( .A(w_cout_5_), .B(_133_), .C(_134_), .Y(_0__24_) );
INVX1 INVX1_29 ( .A(_33__2_), .Y(_135_) );
NAND2X1 NAND2X1_29 ( .A(w_cout_5_), .B(_34__2_), .Y(_136_) );
OAI21X1 OAI21X1_29 ( .A(w_cout_5_), .B(_135_), .C(_136_), .Y(_0__25_) );
INVX1 INVX1_30 ( .A(_33__3_), .Y(_137_) );
NAND2X1 NAND2X1_30 ( .A(w_cout_5_), .B(_34__3_), .Y(_138_) );
OAI21X1 OAI21X1_30 ( .A(w_cout_5_), .B(_137_), .C(_138_), .Y(_0__26_) );
INVX1 INVX1_31 ( .A(_37_), .Y(_139_) );
NAND2X1 NAND2X1_31 ( .A(_38_), .B(w_cout_6_), .Y(_140_) );
OAI21X1 OAI21X1_31 ( .A(w_cout_6_), .B(_139_), .C(_140_), .Y(w_cout_7_) );
INVX1 INVX1_32 ( .A(_39__0_), .Y(_141_) );
NAND2X1 NAND2X1_32 ( .A(_40__0_), .B(w_cout_6_), .Y(_142_) );
OAI21X1 OAI21X1_32 ( .A(w_cout_6_), .B(_141_), .C(_142_), .Y(_0__27_) );
INVX1 INVX1_33 ( .A(_39__1_), .Y(_143_) );
NAND2X1 NAND2X1_33 ( .A(w_cout_6_), .B(_40__1_), .Y(_144_) );
OAI21X1 OAI21X1_33 ( .A(w_cout_6_), .B(_143_), .C(_144_), .Y(_0__28_) );
INVX1 INVX1_34 ( .A(_39__2_), .Y(_145_) );
NAND2X1 NAND2X1_34 ( .A(w_cout_6_), .B(_40__2_), .Y(_146_) );
OAI21X1 OAI21X1_34 ( .A(w_cout_6_), .B(_145_), .C(_146_), .Y(_0__29_) );
INVX1 INVX1_35 ( .A(_39__3_), .Y(_147_) );
NAND2X1 NAND2X1_35 ( .A(w_cout_6_), .B(_40__3_), .Y(_148_) );
OAI21X1 OAI21X1_35 ( .A(w_cout_6_), .B(_147_), .C(_148_), .Y(_0__30_) );
INVX1 INVX1_36 ( .A(_43_), .Y(_149_) );
NAND2X1 NAND2X1_36 ( .A(_44_), .B(w_cout_7_), .Y(_150_) );
OAI21X1 OAI21X1_36 ( .A(w_cout_7_), .B(_149_), .C(_150_), .Y(w_cout_8_) );
INVX1 INVX1_37 ( .A(_45__0_), .Y(_151_) );
NAND2X1 NAND2X1_37 ( .A(_46__0_), .B(w_cout_7_), .Y(_152_) );
OAI21X1 OAI21X1_37 ( .A(w_cout_7_), .B(_151_), .C(_152_), .Y(_0__31_) );
INVX1 INVX1_38 ( .A(_45__1_), .Y(_153_) );
NAND2X1 NAND2X1_38 ( .A(w_cout_7_), .B(_46__1_), .Y(_154_) );
OAI21X1 OAI21X1_38 ( .A(w_cout_7_), .B(_153_), .C(_154_), .Y(_0__32_) );
INVX1 INVX1_39 ( .A(_45__2_), .Y(_155_) );
NAND2X1 NAND2X1_39 ( .A(w_cout_7_), .B(_46__2_), .Y(_156_) );
OAI21X1 OAI21X1_39 ( .A(w_cout_7_), .B(_155_), .C(_156_), .Y(_0__33_) );
INVX1 INVX1_40 ( .A(_45__3_), .Y(_157_) );
NAND2X1 NAND2X1_40 ( .A(w_cout_7_), .B(_46__3_), .Y(_158_) );
OAI21X1 OAI21X1_40 ( .A(w_cout_7_), .B(_157_), .C(_158_), .Y(_0__34_) );
INVX1 INVX1_41 ( .A(_49_), .Y(_159_) );
NAND2X1 NAND2X1_41 ( .A(_50_), .B(w_cout_8_), .Y(_160_) );
OAI21X1 OAI21X1_41 ( .A(w_cout_8_), .B(_159_), .C(_160_), .Y(w_cout_9_) );
INVX1 INVX1_42 ( .A(_51__0_), .Y(_161_) );
NAND2X1 NAND2X1_42 ( .A(_52__0_), .B(w_cout_8_), .Y(_162_) );
OAI21X1 OAI21X1_42 ( .A(w_cout_8_), .B(_161_), .C(_162_), .Y(_0__35_) );
INVX1 INVX1_43 ( .A(_51__1_), .Y(_163_) );
NAND2X1 NAND2X1_43 ( .A(w_cout_8_), .B(_52__1_), .Y(_164_) );
OAI21X1 OAI21X1_43 ( .A(w_cout_8_), .B(_163_), .C(_164_), .Y(_0__36_) );
INVX1 INVX1_44 ( .A(_51__2_), .Y(_165_) );
NAND2X1 NAND2X1_44 ( .A(w_cout_8_), .B(_52__2_), .Y(_166_) );
OAI21X1 OAI21X1_44 ( .A(w_cout_8_), .B(_165_), .C(_166_), .Y(_0__37_) );
INVX1 INVX1_45 ( .A(_51__3_), .Y(_167_) );
NAND2X1 NAND2X1_45 ( .A(w_cout_8_), .B(_52__3_), .Y(_168_) );
OAI21X1 OAI21X1_45 ( .A(w_cout_8_), .B(_167_), .C(_168_), .Y(_0__38_) );
INVX1 INVX1_46 ( .A(_55_), .Y(_169_) );
NAND2X1 NAND2X1_46 ( .A(_56_), .B(w_cout_9_), .Y(_170_) );
OAI21X1 OAI21X1_46 ( .A(w_cout_9_), .B(_169_), .C(_170_), .Y(w_cout_10_) );
INVX1 INVX1_47 ( .A(_57__0_), .Y(_171_) );
NAND2X1 NAND2X1_47 ( .A(_58__0_), .B(w_cout_9_), .Y(_172_) );
OAI21X1 OAI21X1_47 ( .A(w_cout_9_), .B(_171_), .C(_172_), .Y(_0__39_) );
INVX1 INVX1_48 ( .A(_57__1_), .Y(_173_) );
NAND2X1 NAND2X1_48 ( .A(w_cout_9_), .B(_58__1_), .Y(_174_) );
OAI21X1 OAI21X1_48 ( .A(w_cout_9_), .B(_173_), .C(_174_), .Y(_0__40_) );
INVX1 INVX1_49 ( .A(_57__2_), .Y(_175_) );
NAND2X1 NAND2X1_49 ( .A(w_cout_9_), .B(_58__2_), .Y(_176_) );
OAI21X1 OAI21X1_49 ( .A(w_cout_9_), .B(_175_), .C(_176_), .Y(_0__41_) );
INVX1 INVX1_50 ( .A(_57__3_), .Y(_177_) );
NAND2X1 NAND2X1_50 ( .A(w_cout_9_), .B(_58__3_), .Y(_178_) );
OAI21X1 OAI21X1_50 ( .A(w_cout_9_), .B(_177_), .C(_178_), .Y(_0__42_) );
INVX1 INVX1_51 ( .A(_61_), .Y(_179_) );
NAND2X1 NAND2X1_51 ( .A(_62_), .B(w_cout_10_), .Y(_180_) );
OAI21X1 OAI21X1_51 ( .A(w_cout_10_), .B(_179_), .C(_180_), .Y(w_cout_11_) );
INVX1 INVX1_52 ( .A(_63__0_), .Y(_181_) );
NAND2X1 NAND2X1_52 ( .A(_64__0_), .B(w_cout_10_), .Y(_182_) );
OAI21X1 OAI21X1_52 ( .A(w_cout_10_), .B(_181_), .C(_182_), .Y(_0__43_) );
INVX1 INVX1_53 ( .A(_63__1_), .Y(_183_) );
NAND2X1 NAND2X1_53 ( .A(w_cout_10_), .B(_64__1_), .Y(_184_) );
OAI21X1 OAI21X1_53 ( .A(w_cout_10_), .B(_183_), .C(_184_), .Y(_0__44_) );
INVX1 INVX1_54 ( .A(_63__2_), .Y(_185_) );
NAND2X1 NAND2X1_54 ( .A(w_cout_10_), .B(_64__2_), .Y(_186_) );
OAI21X1 OAI21X1_54 ( .A(w_cout_10_), .B(_185_), .C(_186_), .Y(_0__45_) );
INVX1 INVX1_55 ( .A(_63__3_), .Y(_187_) );
NAND2X1 NAND2X1_55 ( .A(w_cout_10_), .B(_64__3_), .Y(_188_) );
OAI21X1 OAI21X1_55 ( .A(w_cout_10_), .B(_187_), .C(_188_), .Y(_0__46_) );
INVX1 INVX1_56 ( .A(_67_), .Y(_189_) );
NAND2X1 NAND2X1_56 ( .A(_68_), .B(w_cout_11_), .Y(_190_) );
OAI21X1 OAI21X1_56 ( .A(w_cout_11_), .B(_189_), .C(_190_), .Y(w_cout_12_) );
INVX1 INVX1_57 ( .A(_69__0_), .Y(_191_) );
NAND2X1 NAND2X1_57 ( .A(_70__0_), .B(w_cout_11_), .Y(_192_) );
OAI21X1 OAI21X1_57 ( .A(w_cout_11_), .B(_191_), .C(_192_), .Y(_0__47_) );
INVX1 INVX1_58 ( .A(_69__1_), .Y(_193_) );
NAND2X1 NAND2X1_58 ( .A(w_cout_11_), .B(_70__1_), .Y(_194_) );
OAI21X1 OAI21X1_58 ( .A(w_cout_11_), .B(_193_), .C(_194_), .Y(_0__48_) );
INVX1 INVX1_59 ( .A(_69__2_), .Y(_195_) );
NAND2X1 NAND2X1_59 ( .A(w_cout_11_), .B(_70__2_), .Y(_196_) );
OAI21X1 OAI21X1_59 ( .A(w_cout_11_), .B(_195_), .C(_196_), .Y(_0__49_) );
INVX1 INVX1_60 ( .A(_69__3_), .Y(_197_) );
NAND2X1 NAND2X1_60 ( .A(w_cout_11_), .B(_70__3_), .Y(_198_) );
OAI21X1 OAI21X1_60 ( .A(w_cout_11_), .B(_197_), .C(_198_), .Y(_0__50_) );
INVX1 INVX1_61 ( .A(_73_), .Y(_199_) );
NAND2X1 NAND2X1_61 ( .A(_74_), .B(w_cout_12_), .Y(_200_) );
OAI21X1 OAI21X1_61 ( .A(w_cout_12_), .B(_199_), .C(_200_), .Y(w_cout_13_) );
INVX1 INVX1_62 ( .A(_75__0_), .Y(_201_) );
NAND2X1 NAND2X1_62 ( .A(_76__0_), .B(w_cout_12_), .Y(_202_) );
OAI21X1 OAI21X1_62 ( .A(w_cout_12_), .B(_201_), .C(_202_), .Y(_0__51_) );
INVX1 INVX1_63 ( .A(_75__1_), .Y(_203_) );
NAND2X1 NAND2X1_63 ( .A(w_cout_12_), .B(_76__1_), .Y(_204_) );
OAI21X1 OAI21X1_63 ( .A(w_cout_12_), .B(_203_), .C(_204_), .Y(_0__52_) );
INVX1 INVX1_64 ( .A(_75__2_), .Y(_205_) );
NAND2X1 NAND2X1_64 ( .A(w_cout_12_), .B(_76__2_), .Y(_206_) );
OAI21X1 OAI21X1_64 ( .A(w_cout_12_), .B(_205_), .C(_206_), .Y(_0__53_) );
INVX1 INVX1_65 ( .A(_75__3_), .Y(_207_) );
NAND2X1 NAND2X1_65 ( .A(w_cout_12_), .B(_76__3_), .Y(_208_) );
OAI21X1 OAI21X1_65 ( .A(w_cout_12_), .B(_207_), .C(_208_), .Y(_0__54_) );
INVX1 INVX1_66 ( .A(1'b0), .Y(_212_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_213_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_214_) );
NAND3X1 NAND3X1_1 ( .A(_212_), .B(_214_), .C(_213_), .Y(_215_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_209_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_210_) );
OAI21X1 OAI21X1_66 ( .A(_209_), .B(_210_), .C(1'b0), .Y(_211_) );
NAND2X1 NAND2X1_67 ( .A(_211_), .B(_215_), .Y(_3__0_) );
OAI21X1 OAI21X1_67 ( .A(_212_), .B(_209_), .C(_214_), .Y(_5__1_) );
INVX1 INVX1_67 ( .A(_5__1_), .Y(_219_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_220_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_221_) );
NAND3X1 NAND3X1_2 ( .A(_219_), .B(_221_), .C(_220_), .Y(_222_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_216_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_217_) );
OAI21X1 OAI21X1_68 ( .A(_216_), .B(_217_), .C(_5__1_), .Y(_218_) );
NAND2X1 NAND2X1_69 ( .A(_218_), .B(_222_), .Y(_3__1_) );
OAI21X1 OAI21X1_69 ( .A(_219_), .B(_216_), .C(_221_), .Y(_5__2_) );
INVX1 INVX1_68 ( .A(_5__2_), .Y(_226_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_227_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_228_) );
NAND3X1 NAND3X1_3 ( .A(_226_), .B(_228_), .C(_227_), .Y(_229_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_223_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_224_) );
OAI21X1 OAI21X1_70 ( .A(_223_), .B(_224_), .C(_5__2_), .Y(_225_) );
NAND2X1 NAND2X1_71 ( .A(_225_), .B(_229_), .Y(_3__2_) );
OAI21X1 OAI21X1_71 ( .A(_226_), .B(_223_), .C(_228_), .Y(_5__3_) );
INVX1 INVX1_69 ( .A(_5__3_), .Y(_233_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_234_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_235_) );
NAND3X1 NAND3X1_4 ( .A(_233_), .B(_235_), .C(_234_), .Y(_236_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_230_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_231_) );
OAI21X1 OAI21X1_72 ( .A(_230_), .B(_231_), .C(_5__3_), .Y(_232_) );
NAND2X1 NAND2X1_73 ( .A(_232_), .B(_236_), .Y(_3__3_) );
OAI21X1 OAI21X1_73 ( .A(_233_), .B(_230_), .C(_235_), .Y(_1_) );
INVX1 INVX1_70 ( .A(1'b1), .Y(_240_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_241_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_242_) );
NAND3X1 NAND3X1_5 ( .A(_240_), .B(_242_), .C(_241_), .Y(_243_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_237_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_238_) );
OAI21X1 OAI21X1_74 ( .A(_237_), .B(_238_), .C(1'b1), .Y(_239_) );
NAND2X1 NAND2X1_75 ( .A(_239_), .B(_243_), .Y(_4__0_) );
OAI21X1 OAI21X1_75 ( .A(_240_), .B(_237_), .C(_242_), .Y(_6__1_) );
INVX1 INVX1_71 ( .A(_6__1_), .Y(_247_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_248_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_249_) );
NAND3X1 NAND3X1_6 ( .A(_247_), .B(_249_), .C(_248_), .Y(_250_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_244_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_245_) );
OAI21X1 OAI21X1_76 ( .A(_244_), .B(_245_), .C(_6__1_), .Y(_246_) );
NAND2X1 NAND2X1_77 ( .A(_246_), .B(_250_), .Y(_4__1_) );
OAI21X1 OAI21X1_77 ( .A(_247_), .B(_244_), .C(_249_), .Y(_6__2_) );
INVX1 INVX1_72 ( .A(_6__2_), .Y(_254_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_255_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_256_) );
NAND3X1 NAND3X1_7 ( .A(_254_), .B(_256_), .C(_255_), .Y(_257_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_251_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_252_) );
OAI21X1 OAI21X1_78 ( .A(_251_), .B(_252_), .C(_6__2_), .Y(_253_) );
NAND2X1 NAND2X1_79 ( .A(_253_), .B(_257_), .Y(_4__2_) );
OAI21X1 OAI21X1_79 ( .A(_254_), .B(_251_), .C(_256_), .Y(_6__3_) );
INVX1 INVX1_73 ( .A(_6__3_), .Y(_261_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_262_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_263_) );
NAND3X1 NAND3X1_8 ( .A(_261_), .B(_263_), .C(_262_), .Y(_264_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_258_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_259_) );
OAI21X1 OAI21X1_80 ( .A(_258_), .B(_259_), .C(_6__3_), .Y(_260_) );
NAND2X1 NAND2X1_81 ( .A(_260_), .B(_264_), .Y(_4__3_) );
OAI21X1 OAI21X1_81 ( .A(_261_), .B(_258_), .C(_263_), .Y(_2_) );
INVX1 INVX1_74 ( .A(1'b0), .Y(_268_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_269_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_270_) );
NAND3X1 NAND3X1_9 ( .A(_268_), .B(_270_), .C(_269_), .Y(_271_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_265_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_266_) );
OAI21X1 OAI21X1_82 ( .A(_265_), .B(_266_), .C(1'b0), .Y(_267_) );
NAND2X1 NAND2X1_83 ( .A(_267_), .B(_271_), .Y(_9__0_) );
OAI21X1 OAI21X1_83 ( .A(_268_), .B(_265_), .C(_270_), .Y(_11__1_) );
INVX1 INVX1_75 ( .A(_11__1_), .Y(_275_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_276_) );
NAND2X1 NAND2X1_84 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_277_) );
NAND3X1 NAND3X1_10 ( .A(_275_), .B(_277_), .C(_276_), .Y(_278_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_272_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_273_) );
OAI21X1 OAI21X1_84 ( .A(_272_), .B(_273_), .C(_11__1_), .Y(_274_) );
NAND2X1 NAND2X1_85 ( .A(_274_), .B(_278_), .Y(_9__1_) );
OAI21X1 OAI21X1_85 ( .A(_275_), .B(_272_), .C(_277_), .Y(_11__2_) );
INVX1 INVX1_76 ( .A(_11__2_), .Y(_282_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_283_) );
NAND2X1 NAND2X1_86 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_284_) );
NAND3X1 NAND3X1_11 ( .A(_282_), .B(_284_), .C(_283_), .Y(_285_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_279_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_280_) );
OAI21X1 OAI21X1_86 ( .A(_279_), .B(_280_), .C(_11__2_), .Y(_281_) );
NAND2X1 NAND2X1_87 ( .A(_281_), .B(_285_), .Y(_9__2_) );
OAI21X1 OAI21X1_87 ( .A(_282_), .B(_279_), .C(_284_), .Y(_11__3_) );
INVX1 INVX1_77 ( .A(_11__3_), .Y(_289_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_290_) );
NAND2X1 NAND2X1_88 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_291_) );
NAND3X1 NAND3X1_12 ( .A(_289_), .B(_291_), .C(_290_), .Y(_292_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_286_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_287_) );
OAI21X1 OAI21X1_88 ( .A(_286_), .B(_287_), .C(_11__3_), .Y(_288_) );
NAND2X1 NAND2X1_89 ( .A(_288_), .B(_292_), .Y(_9__3_) );
OAI21X1 OAI21X1_89 ( .A(_289_), .B(_286_), .C(_291_), .Y(_7_) );
INVX1 INVX1_78 ( .A(1'b1), .Y(_296_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_297_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_298_) );
NAND3X1 NAND3X1_13 ( .A(_296_), .B(_298_), .C(_297_), .Y(_299_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_293_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_294_) );
OAI21X1 OAI21X1_90 ( .A(_293_), .B(_294_), .C(1'b1), .Y(_295_) );
NAND2X1 NAND2X1_91 ( .A(_295_), .B(_299_), .Y(_10__0_) );
OAI21X1 OAI21X1_91 ( .A(_296_), .B(_293_), .C(_298_), .Y(_12__1_) );
INVX1 INVX1_79 ( .A(_12__1_), .Y(_303_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_304_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_305_) );
NAND3X1 NAND3X1_14 ( .A(_303_), .B(_305_), .C(_304_), .Y(_306_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_300_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_301_) );
OAI21X1 OAI21X1_92 ( .A(_300_), .B(_301_), .C(_12__1_), .Y(_302_) );
NAND2X1 NAND2X1_93 ( .A(_302_), .B(_306_), .Y(_10__1_) );
OAI21X1 OAI21X1_93 ( .A(_303_), .B(_300_), .C(_305_), .Y(_12__2_) );
INVX1 INVX1_80 ( .A(_12__2_), .Y(_310_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_311_) );
NAND2X1 NAND2X1_94 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_312_) );
NAND3X1 NAND3X1_15 ( .A(_310_), .B(_312_), .C(_311_), .Y(_313_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_307_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_308_) );
OAI21X1 OAI21X1_94 ( .A(_307_), .B(_308_), .C(_12__2_), .Y(_309_) );
NAND2X1 NAND2X1_95 ( .A(_309_), .B(_313_), .Y(_10__2_) );
OAI21X1 OAI21X1_95 ( .A(_310_), .B(_307_), .C(_312_), .Y(_12__3_) );
INVX1 INVX1_81 ( .A(_12__3_), .Y(_317_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_318_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_319_) );
NAND3X1 NAND3X1_16 ( .A(_317_), .B(_319_), .C(_318_), .Y(_320_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_314_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_315_) );
OAI21X1 OAI21X1_96 ( .A(_314_), .B(_315_), .C(_12__3_), .Y(_316_) );
NAND2X1 NAND2X1_97 ( .A(_316_), .B(_320_), .Y(_10__3_) );
OAI21X1 OAI21X1_97 ( .A(_317_), .B(_314_), .C(_319_), .Y(_8_) );
INVX1 INVX1_82 ( .A(1'b0), .Y(_324_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_325_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_326_) );
NAND3X1 NAND3X1_17 ( .A(_324_), .B(_326_), .C(_325_), .Y(_327_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_321_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_322_) );
OAI21X1 OAI21X1_98 ( .A(_321_), .B(_322_), .C(1'b0), .Y(_323_) );
NAND2X1 NAND2X1_99 ( .A(_323_), .B(_327_), .Y(_15__0_) );
OAI21X1 OAI21X1_99 ( .A(_324_), .B(_321_), .C(_326_), .Y(_17__1_) );
INVX1 INVX1_83 ( .A(_17__1_), .Y(_331_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_332_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_333_) );
NAND3X1 NAND3X1_18 ( .A(_331_), .B(_333_), .C(_332_), .Y(_334_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_328_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_329_) );
OAI21X1 OAI21X1_100 ( .A(_328_), .B(_329_), .C(_17__1_), .Y(_330_) );
NAND2X1 NAND2X1_101 ( .A(_330_), .B(_334_), .Y(_15__1_) );
OAI21X1 OAI21X1_101 ( .A(_331_), .B(_328_), .C(_333_), .Y(_17__2_) );
INVX1 INVX1_84 ( .A(_17__2_), .Y(_338_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_339_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_340_) );
NAND3X1 NAND3X1_19 ( .A(_338_), .B(_340_), .C(_339_), .Y(_341_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_335_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_336_) );
OAI21X1 OAI21X1_102 ( .A(_335_), .B(_336_), .C(_17__2_), .Y(_337_) );
NAND2X1 NAND2X1_103 ( .A(_337_), .B(_341_), .Y(_15__2_) );
OAI21X1 OAI21X1_103 ( .A(_338_), .B(_335_), .C(_340_), .Y(_17__3_) );
INVX1 INVX1_85 ( .A(_17__3_), .Y(_345_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_346_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_347_) );
NAND3X1 NAND3X1_20 ( .A(_345_), .B(_347_), .C(_346_), .Y(_348_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_342_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_343_) );
OAI21X1 OAI21X1_104 ( .A(_342_), .B(_343_), .C(_17__3_), .Y(_344_) );
NAND2X1 NAND2X1_105 ( .A(_344_), .B(_348_), .Y(_15__3_) );
OAI21X1 OAI21X1_105 ( .A(_345_), .B(_342_), .C(_347_), .Y(_13_) );
INVX1 INVX1_86 ( .A(1'b1), .Y(_352_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_353_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_354_) );
NAND3X1 NAND3X1_21 ( .A(_352_), .B(_354_), .C(_353_), .Y(_355_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_349_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_350_) );
OAI21X1 OAI21X1_106 ( .A(_349_), .B(_350_), .C(1'b1), .Y(_351_) );
NAND2X1 NAND2X1_107 ( .A(_351_), .B(_355_), .Y(_16__0_) );
OAI21X1 OAI21X1_107 ( .A(_352_), .B(_349_), .C(_354_), .Y(_18__1_) );
INVX1 INVX1_87 ( .A(_18__1_), .Y(_359_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_360_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_361_) );
NAND3X1 NAND3X1_22 ( .A(_359_), .B(_361_), .C(_360_), .Y(_362_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_356_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_357_) );
OAI21X1 OAI21X1_108 ( .A(_356_), .B(_357_), .C(_18__1_), .Y(_358_) );
NAND2X1 NAND2X1_109 ( .A(_358_), .B(_362_), .Y(_16__1_) );
OAI21X1 OAI21X1_109 ( .A(_359_), .B(_356_), .C(_361_), .Y(_18__2_) );
INVX1 INVX1_88 ( .A(_18__2_), .Y(_366_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_367_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_368_) );
NAND3X1 NAND3X1_23 ( .A(_366_), .B(_368_), .C(_367_), .Y(_369_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_363_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_364_) );
OAI21X1 OAI21X1_110 ( .A(_363_), .B(_364_), .C(_18__2_), .Y(_365_) );
NAND2X1 NAND2X1_111 ( .A(_365_), .B(_369_), .Y(_16__2_) );
OAI21X1 OAI21X1_111 ( .A(_366_), .B(_363_), .C(_368_), .Y(_18__3_) );
INVX1 INVX1_89 ( .A(_18__3_), .Y(_373_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_374_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_375_) );
NAND3X1 NAND3X1_24 ( .A(_373_), .B(_375_), .C(_374_), .Y(_376_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_370_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_371_) );
OAI21X1 OAI21X1_112 ( .A(_370_), .B(_371_), .C(_18__3_), .Y(_372_) );
NAND2X1 NAND2X1_113 ( .A(_372_), .B(_376_), .Y(_16__3_) );
OAI21X1 OAI21X1_113 ( .A(_373_), .B(_370_), .C(_375_), .Y(_14_) );
INVX1 INVX1_90 ( .A(1'b0), .Y(_380_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_381_) );
NAND2X1 NAND2X1_114 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_382_) );
NAND3X1 NAND3X1_25 ( .A(_380_), .B(_382_), .C(_381_), .Y(_383_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_377_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_378_) );
OAI21X1 OAI21X1_114 ( .A(_377_), .B(_378_), .C(1'b0), .Y(_379_) );
NAND2X1 NAND2X1_115 ( .A(_379_), .B(_383_), .Y(_21__0_) );
OAI21X1 OAI21X1_115 ( .A(_380_), .B(_377_), .C(_382_), .Y(_23__1_) );
INVX1 INVX1_91 ( .A(_23__1_), .Y(_387_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_388_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_389_) );
NAND3X1 NAND3X1_26 ( .A(_387_), .B(_389_), .C(_388_), .Y(_390_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_384_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_385_) );
OAI21X1 OAI21X1_116 ( .A(_384_), .B(_385_), .C(_23__1_), .Y(_386_) );
NAND2X1 NAND2X1_117 ( .A(_386_), .B(_390_), .Y(_21__1_) );
OAI21X1 OAI21X1_117 ( .A(_387_), .B(_384_), .C(_389_), .Y(_23__2_) );
INVX1 INVX1_92 ( .A(_23__2_), .Y(_394_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_395_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_396_) );
NAND3X1 NAND3X1_27 ( .A(_394_), .B(_396_), .C(_395_), .Y(_397_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_391_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_392_) );
OAI21X1 OAI21X1_118 ( .A(_391_), .B(_392_), .C(_23__2_), .Y(_393_) );
NAND2X1 NAND2X1_119 ( .A(_393_), .B(_397_), .Y(_21__2_) );
OAI21X1 OAI21X1_119 ( .A(_394_), .B(_391_), .C(_396_), .Y(_23__3_) );
INVX1 INVX1_93 ( .A(_23__3_), .Y(_401_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_402_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_403_) );
NAND3X1 NAND3X1_28 ( .A(_401_), .B(_403_), .C(_402_), .Y(_404_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_398_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_399_) );
OAI21X1 OAI21X1_120 ( .A(_398_), .B(_399_), .C(_23__3_), .Y(_400_) );
NAND2X1 NAND2X1_121 ( .A(_400_), .B(_404_), .Y(_21__3_) );
OAI21X1 OAI21X1_121 ( .A(_401_), .B(_398_), .C(_403_), .Y(_19_) );
INVX1 INVX1_94 ( .A(1'b1), .Y(_408_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_409_) );
NAND2X1 NAND2X1_122 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_410_) );
NAND3X1 NAND3X1_29 ( .A(_408_), .B(_410_), .C(_409_), .Y(_411_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_405_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_406_) );
OAI21X1 OAI21X1_122 ( .A(_405_), .B(_406_), .C(1'b1), .Y(_407_) );
NAND2X1 NAND2X1_123 ( .A(_407_), .B(_411_), .Y(_22__0_) );
OAI21X1 OAI21X1_123 ( .A(_408_), .B(_405_), .C(_410_), .Y(_24__1_) );
INVX1 INVX1_95 ( .A(_24__1_), .Y(_415_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_416_) );
NAND2X1 NAND2X1_124 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_417_) );
NAND3X1 NAND3X1_30 ( .A(_415_), .B(_417_), .C(_416_), .Y(_418_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_412_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_413_) );
OAI21X1 OAI21X1_124 ( .A(_412_), .B(_413_), .C(_24__1_), .Y(_414_) );
NAND2X1 NAND2X1_125 ( .A(_414_), .B(_418_), .Y(_22__1_) );
OAI21X1 OAI21X1_125 ( .A(_415_), .B(_412_), .C(_417_), .Y(_24__2_) );
INVX1 INVX1_96 ( .A(_24__2_), .Y(_422_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_423_) );
NAND2X1 NAND2X1_126 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_424_) );
NAND3X1 NAND3X1_31 ( .A(_422_), .B(_424_), .C(_423_), .Y(_425_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_419_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_420_) );
OAI21X1 OAI21X1_126 ( .A(_419_), .B(_420_), .C(_24__2_), .Y(_421_) );
NAND2X1 NAND2X1_127 ( .A(_421_), .B(_425_), .Y(_22__2_) );
OAI21X1 OAI21X1_127 ( .A(_422_), .B(_419_), .C(_424_), .Y(_24__3_) );
INVX1 INVX1_97 ( .A(_24__3_), .Y(_429_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_430_) );
NAND2X1 NAND2X1_128 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_431_) );
NAND3X1 NAND3X1_32 ( .A(_429_), .B(_431_), .C(_430_), .Y(_432_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_426_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_427_) );
OAI21X1 OAI21X1_128 ( .A(_426_), .B(_427_), .C(_24__3_), .Y(_428_) );
NAND2X1 NAND2X1_129 ( .A(_428_), .B(_432_), .Y(_22__3_) );
OAI21X1 OAI21X1_129 ( .A(_429_), .B(_426_), .C(_431_), .Y(_20_) );
INVX1 INVX1_98 ( .A(1'b0), .Y(_436_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_437_) );
NAND2X1 NAND2X1_130 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_438_) );
NAND3X1 NAND3X1_33 ( .A(_436_), .B(_438_), .C(_437_), .Y(_439_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_433_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_434_) );
OAI21X1 OAI21X1_130 ( .A(_433_), .B(_434_), .C(1'b0), .Y(_435_) );
NAND2X1 NAND2X1_131 ( .A(_435_), .B(_439_), .Y(_27__0_) );
OAI21X1 OAI21X1_131 ( .A(_436_), .B(_433_), .C(_438_), .Y(_29__1_) );
INVX1 INVX1_99 ( .A(_29__1_), .Y(_443_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_444_) );
NAND2X1 NAND2X1_132 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_445_) );
NAND3X1 NAND3X1_34 ( .A(_443_), .B(_445_), .C(_444_), .Y(_446_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_440_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_441_) );
OAI21X1 OAI21X1_132 ( .A(_440_), .B(_441_), .C(_29__1_), .Y(_442_) );
NAND2X1 NAND2X1_133 ( .A(_442_), .B(_446_), .Y(_27__1_) );
OAI21X1 OAI21X1_133 ( .A(_443_), .B(_440_), .C(_445_), .Y(_29__2_) );
INVX1 INVX1_100 ( .A(_29__2_), .Y(_450_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_451_) );
NAND2X1 NAND2X1_134 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_452_) );
NAND3X1 NAND3X1_35 ( .A(_450_), .B(_452_), .C(_451_), .Y(_453_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_447_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_448_) );
OAI21X1 OAI21X1_134 ( .A(_447_), .B(_448_), .C(_29__2_), .Y(_449_) );
NAND2X1 NAND2X1_135 ( .A(_449_), .B(_453_), .Y(_27__2_) );
OAI21X1 OAI21X1_135 ( .A(_450_), .B(_447_), .C(_452_), .Y(_29__3_) );
INVX1 INVX1_101 ( .A(_29__3_), .Y(_457_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_458_) );
NAND2X1 NAND2X1_136 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_459_) );
NAND3X1 NAND3X1_36 ( .A(_457_), .B(_459_), .C(_458_), .Y(_460_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_454_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_455_) );
OAI21X1 OAI21X1_136 ( .A(_454_), .B(_455_), .C(_29__3_), .Y(_456_) );
NAND2X1 NAND2X1_137 ( .A(_456_), .B(_460_), .Y(_27__3_) );
OAI21X1 OAI21X1_137 ( .A(_457_), .B(_454_), .C(_459_), .Y(_25_) );
INVX1 INVX1_102 ( .A(1'b1), .Y(_464_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_465_) );
NAND2X1 NAND2X1_138 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_466_) );
NAND3X1 NAND3X1_37 ( .A(_464_), .B(_466_), .C(_465_), .Y(_467_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_461_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_462_) );
OAI21X1 OAI21X1_138 ( .A(_461_), .B(_462_), .C(1'b1), .Y(_463_) );
NAND2X1 NAND2X1_139 ( .A(_463_), .B(_467_), .Y(_28__0_) );
OAI21X1 OAI21X1_139 ( .A(_464_), .B(_461_), .C(_466_), .Y(_30__1_) );
INVX1 INVX1_103 ( .A(_30__1_), .Y(_471_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_472_) );
NAND2X1 NAND2X1_140 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_473_) );
NAND3X1 NAND3X1_38 ( .A(_471_), .B(_473_), .C(_472_), .Y(_474_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_468_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_469_) );
OAI21X1 OAI21X1_140 ( .A(_468_), .B(_469_), .C(_30__1_), .Y(_470_) );
NAND2X1 NAND2X1_141 ( .A(_470_), .B(_474_), .Y(_28__1_) );
OAI21X1 OAI21X1_141 ( .A(_471_), .B(_468_), .C(_473_), .Y(_30__2_) );
INVX1 INVX1_104 ( .A(_30__2_), .Y(_478_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_479_) );
NAND2X1 NAND2X1_142 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_480_) );
NAND3X1 NAND3X1_39 ( .A(_478_), .B(_480_), .C(_479_), .Y(_481_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_475_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_476_) );
OAI21X1 OAI21X1_142 ( .A(_475_), .B(_476_), .C(_30__2_), .Y(_477_) );
NAND2X1 NAND2X1_143 ( .A(_477_), .B(_481_), .Y(_28__2_) );
OAI21X1 OAI21X1_143 ( .A(_478_), .B(_475_), .C(_480_), .Y(_30__3_) );
INVX1 INVX1_105 ( .A(_30__3_), .Y(_485_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_486_) );
NAND2X1 NAND2X1_144 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_487_) );
NAND3X1 NAND3X1_40 ( .A(_485_), .B(_487_), .C(_486_), .Y(_488_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_482_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_483_) );
OAI21X1 OAI21X1_144 ( .A(_482_), .B(_483_), .C(_30__3_), .Y(_484_) );
NAND2X1 NAND2X1_145 ( .A(_484_), .B(_488_), .Y(_28__3_) );
OAI21X1 OAI21X1_145 ( .A(_485_), .B(_482_), .C(_487_), .Y(_26_) );
INVX1 INVX1_106 ( .A(1'b0), .Y(_492_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_493_) );
NAND2X1 NAND2X1_146 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_494_) );
NAND3X1 NAND3X1_41 ( .A(_492_), .B(_494_), .C(_493_), .Y(_495_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_489_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_490_) );
OAI21X1 OAI21X1_146 ( .A(_489_), .B(_490_), .C(1'b0), .Y(_491_) );
NAND2X1 NAND2X1_147 ( .A(_491_), .B(_495_), .Y(_33__0_) );
OAI21X1 OAI21X1_147 ( .A(_492_), .B(_489_), .C(_494_), .Y(_35__1_) );
INVX1 INVX1_107 ( .A(_35__1_), .Y(_499_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_500_) );
NAND2X1 NAND2X1_148 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_501_) );
NAND3X1 NAND3X1_42 ( .A(_499_), .B(_501_), .C(_500_), .Y(_502_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_496_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_497_) );
OAI21X1 OAI21X1_148 ( .A(_496_), .B(_497_), .C(_35__1_), .Y(_498_) );
NAND2X1 NAND2X1_149 ( .A(_498_), .B(_502_), .Y(_33__1_) );
OAI21X1 OAI21X1_149 ( .A(_499_), .B(_496_), .C(_501_), .Y(_35__2_) );
INVX1 INVX1_108 ( .A(_35__2_), .Y(_506_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_507_) );
NAND2X1 NAND2X1_150 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_508_) );
NAND3X1 NAND3X1_43 ( .A(_506_), .B(_508_), .C(_507_), .Y(_509_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_503_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_504_) );
OAI21X1 OAI21X1_150 ( .A(_503_), .B(_504_), .C(_35__2_), .Y(_505_) );
NAND2X1 NAND2X1_151 ( .A(_505_), .B(_509_), .Y(_33__2_) );
OAI21X1 OAI21X1_151 ( .A(_506_), .B(_503_), .C(_508_), .Y(_35__3_) );
INVX1 INVX1_109 ( .A(_35__3_), .Y(_513_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_514_) );
NAND2X1 NAND2X1_152 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_515_) );
NAND3X1 NAND3X1_44 ( .A(_513_), .B(_515_), .C(_514_), .Y(_516_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_510_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_511_) );
OAI21X1 OAI21X1_152 ( .A(_510_), .B(_511_), .C(_35__3_), .Y(_512_) );
NAND2X1 NAND2X1_153 ( .A(_512_), .B(_516_), .Y(_33__3_) );
OAI21X1 OAI21X1_153 ( .A(_513_), .B(_510_), .C(_515_), .Y(_31_) );
INVX1 INVX1_110 ( .A(1'b1), .Y(_520_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_521_) );
NAND2X1 NAND2X1_154 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_522_) );
NAND3X1 NAND3X1_45 ( .A(_520_), .B(_522_), .C(_521_), .Y(_523_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_517_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_518_) );
OAI21X1 OAI21X1_154 ( .A(_517_), .B(_518_), .C(1'b1), .Y(_519_) );
NAND2X1 NAND2X1_155 ( .A(_519_), .B(_523_), .Y(_34__0_) );
OAI21X1 OAI21X1_155 ( .A(_520_), .B(_517_), .C(_522_), .Y(_36__1_) );
INVX1 INVX1_111 ( .A(_36__1_), .Y(_527_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_528_) );
NAND2X1 NAND2X1_156 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_529_) );
NAND3X1 NAND3X1_46 ( .A(_527_), .B(_529_), .C(_528_), .Y(_530_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_524_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_525_) );
OAI21X1 OAI21X1_156 ( .A(_524_), .B(_525_), .C(_36__1_), .Y(_526_) );
NAND2X1 NAND2X1_157 ( .A(_526_), .B(_530_), .Y(_34__1_) );
OAI21X1 OAI21X1_157 ( .A(_527_), .B(_524_), .C(_529_), .Y(_36__2_) );
INVX1 INVX1_112 ( .A(_36__2_), .Y(_534_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_535_) );
NAND2X1 NAND2X1_158 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_536_) );
NAND3X1 NAND3X1_47 ( .A(_534_), .B(_536_), .C(_535_), .Y(_537_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_531_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_532_) );
OAI21X1 OAI21X1_158 ( .A(_531_), .B(_532_), .C(_36__2_), .Y(_533_) );
NAND2X1 NAND2X1_159 ( .A(_533_), .B(_537_), .Y(_34__2_) );
OAI21X1 OAI21X1_159 ( .A(_534_), .B(_531_), .C(_536_), .Y(_36__3_) );
INVX1 INVX1_113 ( .A(_36__3_), .Y(_541_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_542_) );
NAND2X1 NAND2X1_160 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_543_) );
NAND3X1 NAND3X1_48 ( .A(_541_), .B(_543_), .C(_542_), .Y(_544_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_538_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_539_) );
OAI21X1 OAI21X1_160 ( .A(_538_), .B(_539_), .C(_36__3_), .Y(_540_) );
NAND2X1 NAND2X1_161 ( .A(_540_), .B(_544_), .Y(_34__3_) );
OAI21X1 OAI21X1_161 ( .A(_541_), .B(_538_), .C(_543_), .Y(_32_) );
INVX1 INVX1_114 ( .A(1'b0), .Y(_548_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_549_) );
NAND2X1 NAND2X1_162 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_550_) );
NAND3X1 NAND3X1_49 ( .A(_548_), .B(_550_), .C(_549_), .Y(_551_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_545_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_546_) );
OAI21X1 OAI21X1_162 ( .A(_545_), .B(_546_), .C(1'b0), .Y(_547_) );
NAND2X1 NAND2X1_163 ( .A(_547_), .B(_551_), .Y(_39__0_) );
OAI21X1 OAI21X1_163 ( .A(_548_), .B(_545_), .C(_550_), .Y(_41__1_) );
INVX1 INVX1_115 ( .A(_41__1_), .Y(_555_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_556_) );
NAND2X1 NAND2X1_164 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_557_) );
NAND3X1 NAND3X1_50 ( .A(_555_), .B(_557_), .C(_556_), .Y(_558_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_552_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_553_) );
OAI21X1 OAI21X1_164 ( .A(_552_), .B(_553_), .C(_41__1_), .Y(_554_) );
NAND2X1 NAND2X1_165 ( .A(_554_), .B(_558_), .Y(_39__1_) );
OAI21X1 OAI21X1_165 ( .A(_555_), .B(_552_), .C(_557_), .Y(_41__2_) );
INVX1 INVX1_116 ( .A(_41__2_), .Y(_562_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_563_) );
NAND2X1 NAND2X1_166 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_564_) );
NAND3X1 NAND3X1_51 ( .A(_562_), .B(_564_), .C(_563_), .Y(_565_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_559_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_560_) );
OAI21X1 OAI21X1_166 ( .A(_559_), .B(_560_), .C(_41__2_), .Y(_561_) );
NAND2X1 NAND2X1_167 ( .A(_561_), .B(_565_), .Y(_39__2_) );
OAI21X1 OAI21X1_167 ( .A(_562_), .B(_559_), .C(_564_), .Y(_41__3_) );
INVX1 INVX1_117 ( .A(_41__3_), .Y(_569_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_570_) );
NAND2X1 NAND2X1_168 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_571_) );
NAND3X1 NAND3X1_52 ( .A(_569_), .B(_571_), .C(_570_), .Y(_572_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_566_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_567_) );
OAI21X1 OAI21X1_168 ( .A(_566_), .B(_567_), .C(_41__3_), .Y(_568_) );
NAND2X1 NAND2X1_169 ( .A(_568_), .B(_572_), .Y(_39__3_) );
OAI21X1 OAI21X1_169 ( .A(_569_), .B(_566_), .C(_571_), .Y(_37_) );
INVX1 INVX1_118 ( .A(1'b1), .Y(_576_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_577_) );
NAND2X1 NAND2X1_170 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_578_) );
NAND3X1 NAND3X1_53 ( .A(_576_), .B(_578_), .C(_577_), .Y(_579_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_573_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_574_) );
OAI21X1 OAI21X1_170 ( .A(_573_), .B(_574_), .C(1'b1), .Y(_575_) );
NAND2X1 NAND2X1_171 ( .A(_575_), .B(_579_), .Y(_40__0_) );
OAI21X1 OAI21X1_171 ( .A(_576_), .B(_573_), .C(_578_), .Y(_42__1_) );
INVX1 INVX1_119 ( .A(_42__1_), .Y(_583_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_584_) );
NAND2X1 NAND2X1_172 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_585_) );
NAND3X1 NAND3X1_54 ( .A(_583_), .B(_585_), .C(_584_), .Y(_586_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_580_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_581_) );
OAI21X1 OAI21X1_172 ( .A(_580_), .B(_581_), .C(_42__1_), .Y(_582_) );
NAND2X1 NAND2X1_173 ( .A(_582_), .B(_586_), .Y(_40__1_) );
OAI21X1 OAI21X1_173 ( .A(_583_), .B(_580_), .C(_585_), .Y(_42__2_) );
INVX1 INVX1_120 ( .A(_42__2_), .Y(_590_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_591_) );
NAND2X1 NAND2X1_174 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_592_) );
NAND3X1 NAND3X1_55 ( .A(_590_), .B(_592_), .C(_591_), .Y(_593_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_587_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_588_) );
OAI21X1 OAI21X1_174 ( .A(_587_), .B(_588_), .C(_42__2_), .Y(_589_) );
NAND2X1 NAND2X1_175 ( .A(_589_), .B(_593_), .Y(_40__2_) );
OAI21X1 OAI21X1_175 ( .A(_590_), .B(_587_), .C(_592_), .Y(_42__3_) );
INVX1 INVX1_121 ( .A(_42__3_), .Y(_597_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_598_) );
NAND2X1 NAND2X1_176 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_599_) );
NAND3X1 NAND3X1_56 ( .A(_597_), .B(_599_), .C(_598_), .Y(_600_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_594_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_595_) );
OAI21X1 OAI21X1_176 ( .A(_594_), .B(_595_), .C(_42__3_), .Y(_596_) );
NAND2X1 NAND2X1_177 ( .A(_596_), .B(_600_), .Y(_40__3_) );
OAI21X1 OAI21X1_177 ( .A(_597_), .B(_594_), .C(_599_), .Y(_38_) );
INVX1 INVX1_122 ( .A(1'b0), .Y(_604_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_605_) );
NAND2X1 NAND2X1_178 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_606_) );
NAND3X1 NAND3X1_57 ( .A(_604_), .B(_606_), .C(_605_), .Y(_607_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_601_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_602_) );
OAI21X1 OAI21X1_178 ( .A(_601_), .B(_602_), .C(1'b0), .Y(_603_) );
NAND2X1 NAND2X1_179 ( .A(_603_), .B(_607_), .Y(_45__0_) );
OAI21X1 OAI21X1_179 ( .A(_604_), .B(_601_), .C(_606_), .Y(_47__1_) );
INVX1 INVX1_123 ( .A(_47__1_), .Y(_611_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_612_) );
NAND2X1 NAND2X1_180 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_613_) );
NAND3X1 NAND3X1_58 ( .A(_611_), .B(_613_), .C(_612_), .Y(_614_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_608_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_609_) );
OAI21X1 OAI21X1_180 ( .A(_608_), .B(_609_), .C(_47__1_), .Y(_610_) );
NAND2X1 NAND2X1_181 ( .A(_610_), .B(_614_), .Y(_45__1_) );
OAI21X1 OAI21X1_181 ( .A(_611_), .B(_608_), .C(_613_), .Y(_47__2_) );
INVX1 INVX1_124 ( .A(_47__2_), .Y(_618_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_619_) );
NAND2X1 NAND2X1_182 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_620_) );
NAND3X1 NAND3X1_59 ( .A(_618_), .B(_620_), .C(_619_), .Y(_621_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_615_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_616_) );
OAI21X1 OAI21X1_182 ( .A(_615_), .B(_616_), .C(_47__2_), .Y(_617_) );
NAND2X1 NAND2X1_183 ( .A(_617_), .B(_621_), .Y(_45__2_) );
OAI21X1 OAI21X1_183 ( .A(_618_), .B(_615_), .C(_620_), .Y(_47__3_) );
INVX1 INVX1_125 ( .A(_47__3_), .Y(_625_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_626_) );
NAND2X1 NAND2X1_184 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_627_) );
NAND3X1 NAND3X1_60 ( .A(_625_), .B(_627_), .C(_626_), .Y(_628_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_622_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_623_) );
OAI21X1 OAI21X1_184 ( .A(_622_), .B(_623_), .C(_47__3_), .Y(_624_) );
NAND2X1 NAND2X1_185 ( .A(_624_), .B(_628_), .Y(_45__3_) );
OAI21X1 OAI21X1_185 ( .A(_625_), .B(_622_), .C(_627_), .Y(_43_) );
INVX1 INVX1_126 ( .A(1'b1), .Y(_632_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_633_) );
NAND2X1 NAND2X1_186 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_634_) );
NAND3X1 NAND3X1_61 ( .A(_632_), .B(_634_), .C(_633_), .Y(_635_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_629_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_630_) );
OAI21X1 OAI21X1_186 ( .A(_629_), .B(_630_), .C(1'b1), .Y(_631_) );
NAND2X1 NAND2X1_187 ( .A(_631_), .B(_635_), .Y(_46__0_) );
OAI21X1 OAI21X1_187 ( .A(_632_), .B(_629_), .C(_634_), .Y(_48__1_) );
INVX1 INVX1_127 ( .A(_48__1_), .Y(_639_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_640_) );
NAND2X1 NAND2X1_188 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_641_) );
NAND3X1 NAND3X1_62 ( .A(_639_), .B(_641_), .C(_640_), .Y(_642_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_636_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_637_) );
OAI21X1 OAI21X1_188 ( .A(_636_), .B(_637_), .C(_48__1_), .Y(_638_) );
NAND2X1 NAND2X1_189 ( .A(_638_), .B(_642_), .Y(_46__1_) );
OAI21X1 OAI21X1_189 ( .A(_639_), .B(_636_), .C(_641_), .Y(_48__2_) );
INVX1 INVX1_128 ( .A(_48__2_), .Y(_646_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_647_) );
NAND2X1 NAND2X1_190 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_648_) );
NAND3X1 NAND3X1_63 ( .A(_646_), .B(_648_), .C(_647_), .Y(_649_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_643_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_644_) );
OAI21X1 OAI21X1_190 ( .A(_643_), .B(_644_), .C(_48__2_), .Y(_645_) );
NAND2X1 NAND2X1_191 ( .A(_645_), .B(_649_), .Y(_46__2_) );
OAI21X1 OAI21X1_191 ( .A(_646_), .B(_643_), .C(_648_), .Y(_48__3_) );
INVX1 INVX1_129 ( .A(_48__3_), .Y(_653_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_654_) );
NAND2X1 NAND2X1_192 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_655_) );
NAND3X1 NAND3X1_64 ( .A(_653_), .B(_655_), .C(_654_), .Y(_656_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_650_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_651_) );
OAI21X1 OAI21X1_192 ( .A(_650_), .B(_651_), .C(_48__3_), .Y(_652_) );
NAND2X1 NAND2X1_193 ( .A(_652_), .B(_656_), .Y(_46__3_) );
OAI21X1 OAI21X1_193 ( .A(_653_), .B(_650_), .C(_655_), .Y(_44_) );
INVX1 INVX1_130 ( .A(1'b0), .Y(_660_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_661_) );
NAND2X1 NAND2X1_194 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_662_) );
NAND3X1 NAND3X1_65 ( .A(_660_), .B(_662_), .C(_661_), .Y(_663_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_657_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_658_) );
OAI21X1 OAI21X1_194 ( .A(_657_), .B(_658_), .C(1'b0), .Y(_659_) );
NAND2X1 NAND2X1_195 ( .A(_659_), .B(_663_), .Y(_51__0_) );
OAI21X1 OAI21X1_195 ( .A(_660_), .B(_657_), .C(_662_), .Y(_53__1_) );
INVX1 INVX1_131 ( .A(_53__1_), .Y(_667_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_668_) );
NAND2X1 NAND2X1_196 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_669_) );
NAND3X1 NAND3X1_66 ( .A(_667_), .B(_669_), .C(_668_), .Y(_670_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_664_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_665_) );
OAI21X1 OAI21X1_196 ( .A(_664_), .B(_665_), .C(_53__1_), .Y(_666_) );
NAND2X1 NAND2X1_197 ( .A(_666_), .B(_670_), .Y(_51__1_) );
OAI21X1 OAI21X1_197 ( .A(_667_), .B(_664_), .C(_669_), .Y(_53__2_) );
INVX1 INVX1_132 ( .A(_53__2_), .Y(_674_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_675_) );
NAND2X1 NAND2X1_198 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_676_) );
NAND3X1 NAND3X1_67 ( .A(_674_), .B(_676_), .C(_675_), .Y(_677_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_671_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_672_) );
OAI21X1 OAI21X1_198 ( .A(_671_), .B(_672_), .C(_53__2_), .Y(_673_) );
NAND2X1 NAND2X1_199 ( .A(_673_), .B(_677_), .Y(_51__2_) );
OAI21X1 OAI21X1_199 ( .A(_674_), .B(_671_), .C(_676_), .Y(_53__3_) );
INVX1 INVX1_133 ( .A(_53__3_), .Y(_681_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_682_) );
NAND2X1 NAND2X1_200 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_683_) );
NAND3X1 NAND3X1_68 ( .A(_681_), .B(_683_), .C(_682_), .Y(_684_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_678_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_679_) );
OAI21X1 OAI21X1_200 ( .A(_678_), .B(_679_), .C(_53__3_), .Y(_680_) );
NAND2X1 NAND2X1_201 ( .A(_680_), .B(_684_), .Y(_51__3_) );
OAI21X1 OAI21X1_201 ( .A(_681_), .B(_678_), .C(_683_), .Y(_49_) );
INVX1 INVX1_134 ( .A(1'b1), .Y(_688_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_689_) );
NAND2X1 NAND2X1_202 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_690_) );
NAND3X1 NAND3X1_69 ( .A(_688_), .B(_690_), .C(_689_), .Y(_691_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_685_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_686_) );
OAI21X1 OAI21X1_202 ( .A(_685_), .B(_686_), .C(1'b1), .Y(_687_) );
NAND2X1 NAND2X1_203 ( .A(_687_), .B(_691_), .Y(_52__0_) );
OAI21X1 OAI21X1_203 ( .A(_688_), .B(_685_), .C(_690_), .Y(_54__1_) );
INVX1 INVX1_135 ( .A(_54__1_), .Y(_695_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_696_) );
NAND2X1 NAND2X1_204 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_697_) );
NAND3X1 NAND3X1_70 ( .A(_695_), .B(_697_), .C(_696_), .Y(_698_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_692_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_693_) );
OAI21X1 OAI21X1_204 ( .A(_692_), .B(_693_), .C(_54__1_), .Y(_694_) );
NAND2X1 NAND2X1_205 ( .A(_694_), .B(_698_), .Y(_52__1_) );
OAI21X1 OAI21X1_205 ( .A(_695_), .B(_692_), .C(_697_), .Y(_54__2_) );
INVX1 INVX1_136 ( .A(_54__2_), .Y(_702_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_703_) );
NAND2X1 NAND2X1_206 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_704_) );
NAND3X1 NAND3X1_71 ( .A(_702_), .B(_704_), .C(_703_), .Y(_705_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_699_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_700_) );
OAI21X1 OAI21X1_206 ( .A(_699_), .B(_700_), .C(_54__2_), .Y(_701_) );
NAND2X1 NAND2X1_207 ( .A(_701_), .B(_705_), .Y(_52__2_) );
OAI21X1 OAI21X1_207 ( .A(_702_), .B(_699_), .C(_704_), .Y(_54__3_) );
INVX1 INVX1_137 ( .A(_54__3_), .Y(_709_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_710_) );
NAND2X1 NAND2X1_208 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_711_) );
NAND3X1 NAND3X1_72 ( .A(_709_), .B(_711_), .C(_710_), .Y(_712_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_706_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_707_) );
OAI21X1 OAI21X1_208 ( .A(_706_), .B(_707_), .C(_54__3_), .Y(_708_) );
NAND2X1 NAND2X1_209 ( .A(_708_), .B(_712_), .Y(_52__3_) );
OAI21X1 OAI21X1_209 ( .A(_709_), .B(_706_), .C(_711_), .Y(_50_) );
INVX1 INVX1_138 ( .A(1'b0), .Y(_716_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_717_) );
NAND2X1 NAND2X1_210 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_718_) );
NAND3X1 NAND3X1_73 ( .A(_716_), .B(_718_), .C(_717_), .Y(_719_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_713_) );
AND2X2 AND2X2_73 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_714_) );
OAI21X1 OAI21X1_210 ( .A(_713_), .B(_714_), .C(1'b0), .Y(_715_) );
NAND2X1 NAND2X1_211 ( .A(_715_), .B(_719_), .Y(_57__0_) );
OAI21X1 OAI21X1_211 ( .A(_716_), .B(_713_), .C(_718_), .Y(_59__1_) );
INVX1 INVX1_139 ( .A(_59__1_), .Y(_723_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_724_) );
NAND2X1 NAND2X1_212 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_725_) );
NAND3X1 NAND3X1_74 ( .A(_723_), .B(_725_), .C(_724_), .Y(_726_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_720_) );
AND2X2 AND2X2_74 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_721_) );
OAI21X1 OAI21X1_212 ( .A(_720_), .B(_721_), .C(_59__1_), .Y(_722_) );
NAND2X1 NAND2X1_213 ( .A(_722_), .B(_726_), .Y(_57__1_) );
OAI21X1 OAI21X1_213 ( .A(_723_), .B(_720_), .C(_725_), .Y(_59__2_) );
INVX1 INVX1_140 ( .A(_59__2_), .Y(_730_) );
OR2X2 OR2X2_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_731_) );
NAND2X1 NAND2X1_214 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_732_) );
NAND3X1 NAND3X1_75 ( .A(_730_), .B(_732_), .C(_731_), .Y(_733_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_727_) );
AND2X2 AND2X2_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_728_) );
OAI21X1 OAI21X1_214 ( .A(_727_), .B(_728_), .C(_59__2_), .Y(_729_) );
NAND2X1 NAND2X1_215 ( .A(_729_), .B(_733_), .Y(_57__2_) );
OAI21X1 OAI21X1_215 ( .A(_730_), .B(_727_), .C(_732_), .Y(_59__3_) );
INVX1 INVX1_141 ( .A(_59__3_), .Y(_737_) );
OR2X2 OR2X2_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_738_) );
NAND2X1 NAND2X1_216 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_739_) );
NAND3X1 NAND3X1_76 ( .A(_737_), .B(_739_), .C(_738_), .Y(_740_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_734_) );
AND2X2 AND2X2_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_735_) );
OAI21X1 OAI21X1_216 ( .A(_734_), .B(_735_), .C(_59__3_), .Y(_736_) );
NAND2X1 NAND2X1_217 ( .A(_736_), .B(_740_), .Y(_57__3_) );
OAI21X1 OAI21X1_217 ( .A(_737_), .B(_734_), .C(_739_), .Y(_55_) );
INVX1 INVX1_142 ( .A(1'b1), .Y(_744_) );
OR2X2 OR2X2_77 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_745_) );
NAND2X1 NAND2X1_218 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_746_) );
NAND3X1 NAND3X1_77 ( .A(_744_), .B(_746_), .C(_745_), .Y(_747_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_741_) );
AND2X2 AND2X2_77 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_742_) );
OAI21X1 OAI21X1_218 ( .A(_741_), .B(_742_), .C(1'b1), .Y(_743_) );
NAND2X1 NAND2X1_219 ( .A(_743_), .B(_747_), .Y(_58__0_) );
OAI21X1 OAI21X1_219 ( .A(_744_), .B(_741_), .C(_746_), .Y(_60__1_) );
INVX1 INVX1_143 ( .A(_60__1_), .Y(_751_) );
OR2X2 OR2X2_78 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_752_) );
NAND2X1 NAND2X1_220 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_753_) );
NAND3X1 NAND3X1_78 ( .A(_751_), .B(_753_), .C(_752_), .Y(_754_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_748_) );
AND2X2 AND2X2_78 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_749_) );
OAI21X1 OAI21X1_220 ( .A(_748_), .B(_749_), .C(_60__1_), .Y(_750_) );
NAND2X1 NAND2X1_221 ( .A(_750_), .B(_754_), .Y(_58__1_) );
OAI21X1 OAI21X1_221 ( .A(_751_), .B(_748_), .C(_753_), .Y(_60__2_) );
INVX1 INVX1_144 ( .A(_60__2_), .Y(_758_) );
OR2X2 OR2X2_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_759_) );
NAND2X1 NAND2X1_222 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_760_) );
NAND3X1 NAND3X1_79 ( .A(_758_), .B(_760_), .C(_759_), .Y(_761_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_755_) );
AND2X2 AND2X2_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_756_) );
OAI21X1 OAI21X1_222 ( .A(_755_), .B(_756_), .C(_60__2_), .Y(_757_) );
NAND2X1 NAND2X1_223 ( .A(_757_), .B(_761_), .Y(_58__2_) );
OAI21X1 OAI21X1_223 ( .A(_758_), .B(_755_), .C(_760_), .Y(_60__3_) );
INVX1 INVX1_145 ( .A(_60__3_), .Y(_765_) );
OR2X2 OR2X2_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_766_) );
NAND2X1 NAND2X1_224 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_767_) );
NAND3X1 NAND3X1_80 ( .A(_765_), .B(_767_), .C(_766_), .Y(_768_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_762_) );
AND2X2 AND2X2_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_763_) );
OAI21X1 OAI21X1_224 ( .A(_762_), .B(_763_), .C(_60__3_), .Y(_764_) );
NAND2X1 NAND2X1_225 ( .A(_764_), .B(_768_), .Y(_58__3_) );
OAI21X1 OAI21X1_225 ( .A(_765_), .B(_762_), .C(_767_), .Y(_56_) );
INVX1 INVX1_146 ( .A(1'b0), .Y(_772_) );
OR2X2 OR2X2_81 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_773_) );
NAND2X1 NAND2X1_226 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_774_) );
NAND3X1 NAND3X1_81 ( .A(_772_), .B(_774_), .C(_773_), .Y(_775_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_769_) );
AND2X2 AND2X2_81 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_770_) );
OAI21X1 OAI21X1_226 ( .A(_769_), .B(_770_), .C(1'b0), .Y(_771_) );
NAND2X1 NAND2X1_227 ( .A(_771_), .B(_775_), .Y(_63__0_) );
OAI21X1 OAI21X1_227 ( .A(_772_), .B(_769_), .C(_774_), .Y(_65__1_) );
INVX1 INVX1_147 ( .A(_65__1_), .Y(_779_) );
OR2X2 OR2X2_82 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_780_) );
NAND2X1 NAND2X1_228 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_781_) );
NAND3X1 NAND3X1_82 ( .A(_779_), .B(_781_), .C(_780_), .Y(_782_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_776_) );
AND2X2 AND2X2_82 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_777_) );
OAI21X1 OAI21X1_228 ( .A(_776_), .B(_777_), .C(_65__1_), .Y(_778_) );
NAND2X1 NAND2X1_229 ( .A(_778_), .B(_782_), .Y(_63__1_) );
OAI21X1 OAI21X1_229 ( .A(_779_), .B(_776_), .C(_781_), .Y(_65__2_) );
INVX1 INVX1_148 ( .A(_65__2_), .Y(_786_) );
OR2X2 OR2X2_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_787_) );
NAND2X1 NAND2X1_230 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_788_) );
NAND3X1 NAND3X1_83 ( .A(_786_), .B(_788_), .C(_787_), .Y(_789_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_783_) );
AND2X2 AND2X2_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_784_) );
OAI21X1 OAI21X1_230 ( .A(_783_), .B(_784_), .C(_65__2_), .Y(_785_) );
NAND2X1 NAND2X1_231 ( .A(_785_), .B(_789_), .Y(_63__2_) );
OAI21X1 OAI21X1_231 ( .A(_786_), .B(_783_), .C(_788_), .Y(_65__3_) );
INVX1 INVX1_149 ( .A(_65__3_), .Y(_793_) );
OR2X2 OR2X2_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_794_) );
NAND2X1 NAND2X1_232 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_795_) );
NAND3X1 NAND3X1_84 ( .A(_793_), .B(_795_), .C(_794_), .Y(_796_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_790_) );
AND2X2 AND2X2_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_791_) );
OAI21X1 OAI21X1_232 ( .A(_790_), .B(_791_), .C(_65__3_), .Y(_792_) );
NAND2X1 NAND2X1_233 ( .A(_792_), .B(_796_), .Y(_63__3_) );
OAI21X1 OAI21X1_233 ( .A(_793_), .B(_790_), .C(_795_), .Y(_61_) );
INVX1 INVX1_150 ( .A(1'b1), .Y(_800_) );
OR2X2 OR2X2_85 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_801_) );
NAND2X1 NAND2X1_234 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_802_) );
NAND3X1 NAND3X1_85 ( .A(_800_), .B(_802_), .C(_801_), .Y(_803_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_797_) );
AND2X2 AND2X2_85 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_798_) );
OAI21X1 OAI21X1_234 ( .A(_797_), .B(_798_), .C(1'b1), .Y(_799_) );
NAND2X1 NAND2X1_235 ( .A(_799_), .B(_803_), .Y(_64__0_) );
OAI21X1 OAI21X1_235 ( .A(_800_), .B(_797_), .C(_802_), .Y(_66__1_) );
INVX1 INVX1_151 ( .A(_66__1_), .Y(_807_) );
OR2X2 OR2X2_86 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_808_) );
NAND2X1 NAND2X1_236 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_809_) );
NAND3X1 NAND3X1_86 ( .A(_807_), .B(_809_), .C(_808_), .Y(_810_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_804_) );
AND2X2 AND2X2_86 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_805_) );
OAI21X1 OAI21X1_236 ( .A(_804_), .B(_805_), .C(_66__1_), .Y(_806_) );
NAND2X1 NAND2X1_237 ( .A(_806_), .B(_810_), .Y(_64__1_) );
OAI21X1 OAI21X1_237 ( .A(_807_), .B(_804_), .C(_809_), .Y(_66__2_) );
INVX1 INVX1_152 ( .A(_66__2_), .Y(_814_) );
OR2X2 OR2X2_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_815_) );
NAND2X1 NAND2X1_238 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_816_) );
NAND3X1 NAND3X1_87 ( .A(_814_), .B(_816_), .C(_815_), .Y(_817_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_811_) );
AND2X2 AND2X2_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_812_) );
OAI21X1 OAI21X1_238 ( .A(_811_), .B(_812_), .C(_66__2_), .Y(_813_) );
NAND2X1 NAND2X1_239 ( .A(_813_), .B(_817_), .Y(_64__2_) );
OAI21X1 OAI21X1_239 ( .A(_814_), .B(_811_), .C(_816_), .Y(_66__3_) );
INVX1 INVX1_153 ( .A(_66__3_), .Y(_821_) );
OR2X2 OR2X2_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_822_) );
NAND2X1 NAND2X1_240 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_823_) );
NAND3X1 NAND3X1_88 ( .A(_821_), .B(_823_), .C(_822_), .Y(_824_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_818_) );
AND2X2 AND2X2_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_819_) );
OAI21X1 OAI21X1_240 ( .A(_818_), .B(_819_), .C(_66__3_), .Y(_820_) );
NAND2X1 NAND2X1_241 ( .A(_820_), .B(_824_), .Y(_64__3_) );
OAI21X1 OAI21X1_241 ( .A(_821_), .B(_818_), .C(_823_), .Y(_62_) );
INVX1 INVX1_154 ( .A(1'b0), .Y(_828_) );
OR2X2 OR2X2_89 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_829_) );
NAND2X1 NAND2X1_242 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_830_) );
NAND3X1 NAND3X1_89 ( .A(_828_), .B(_830_), .C(_829_), .Y(_831_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_825_) );
AND2X2 AND2X2_89 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_826_) );
OAI21X1 OAI21X1_242 ( .A(_825_), .B(_826_), .C(1'b0), .Y(_827_) );
NAND2X1 NAND2X1_243 ( .A(_827_), .B(_831_), .Y(_69__0_) );
OAI21X1 OAI21X1_243 ( .A(_828_), .B(_825_), .C(_830_), .Y(_71__1_) );
INVX1 INVX1_155 ( .A(_71__1_), .Y(_835_) );
OR2X2 OR2X2_90 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_836_) );
NAND2X1 NAND2X1_244 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_837_) );
NAND3X1 NAND3X1_90 ( .A(_835_), .B(_837_), .C(_836_), .Y(_838_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_832_) );
AND2X2 AND2X2_90 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_833_) );
OAI21X1 OAI21X1_244 ( .A(_832_), .B(_833_), .C(_71__1_), .Y(_834_) );
NAND2X1 NAND2X1_245 ( .A(_834_), .B(_838_), .Y(_69__1_) );
OAI21X1 OAI21X1_245 ( .A(_835_), .B(_832_), .C(_837_), .Y(_71__2_) );
INVX1 INVX1_156 ( .A(_71__2_), .Y(_842_) );
OR2X2 OR2X2_91 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_843_) );
NAND2X1 NAND2X1_246 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_844_) );
NAND3X1 NAND3X1_91 ( .A(_842_), .B(_844_), .C(_843_), .Y(_845_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_839_) );
AND2X2 AND2X2_91 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_840_) );
OAI21X1 OAI21X1_246 ( .A(_839_), .B(_840_), .C(_71__2_), .Y(_841_) );
NAND2X1 NAND2X1_247 ( .A(_841_), .B(_845_), .Y(_69__2_) );
OAI21X1 OAI21X1_247 ( .A(_842_), .B(_839_), .C(_844_), .Y(_71__3_) );
INVX1 INVX1_157 ( .A(_71__3_), .Y(_849_) );
OR2X2 OR2X2_92 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_850_) );
NAND2X1 NAND2X1_248 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_851_) );
NAND3X1 NAND3X1_92 ( .A(_849_), .B(_851_), .C(_850_), .Y(_852_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_846_) );
AND2X2 AND2X2_92 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_847_) );
OAI21X1 OAI21X1_248 ( .A(_846_), .B(_847_), .C(_71__3_), .Y(_848_) );
NAND2X1 NAND2X1_249 ( .A(_848_), .B(_852_), .Y(_69__3_) );
OAI21X1 OAI21X1_249 ( .A(_849_), .B(_846_), .C(_851_), .Y(_67_) );
INVX1 INVX1_158 ( .A(1'b1), .Y(_856_) );
OR2X2 OR2X2_93 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_857_) );
NAND2X1 NAND2X1_250 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_858_) );
NAND3X1 NAND3X1_93 ( .A(_856_), .B(_858_), .C(_857_), .Y(_859_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_853_) );
AND2X2 AND2X2_93 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_854_) );
OAI21X1 OAI21X1_250 ( .A(_853_), .B(_854_), .C(1'b1), .Y(_855_) );
NAND2X1 NAND2X1_251 ( .A(_855_), .B(_859_), .Y(_70__0_) );
OAI21X1 OAI21X1_251 ( .A(_856_), .B(_853_), .C(_858_), .Y(_72__1_) );
INVX1 INVX1_159 ( .A(_72__1_), .Y(_863_) );
OR2X2 OR2X2_94 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_864_) );
NAND2X1 NAND2X1_252 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_865_) );
NAND3X1 NAND3X1_94 ( .A(_863_), .B(_865_), .C(_864_), .Y(_866_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_860_) );
AND2X2 AND2X2_94 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_861_) );
OAI21X1 OAI21X1_252 ( .A(_860_), .B(_861_), .C(_72__1_), .Y(_862_) );
NAND2X1 NAND2X1_253 ( .A(_862_), .B(_866_), .Y(_70__1_) );
OAI21X1 OAI21X1_253 ( .A(_863_), .B(_860_), .C(_865_), .Y(_72__2_) );
INVX1 INVX1_160 ( .A(_72__2_), .Y(_870_) );
OR2X2 OR2X2_95 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_871_) );
NAND2X1 NAND2X1_254 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_872_) );
NAND3X1 NAND3X1_95 ( .A(_870_), .B(_872_), .C(_871_), .Y(_873_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_867_) );
AND2X2 AND2X2_95 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_868_) );
OAI21X1 OAI21X1_254 ( .A(_867_), .B(_868_), .C(_72__2_), .Y(_869_) );
NAND2X1 NAND2X1_255 ( .A(_869_), .B(_873_), .Y(_70__2_) );
OAI21X1 OAI21X1_255 ( .A(_870_), .B(_867_), .C(_872_), .Y(_72__3_) );
INVX1 INVX1_161 ( .A(_72__3_), .Y(_877_) );
OR2X2 OR2X2_96 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_878_) );
NAND2X1 NAND2X1_256 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_879_) );
NAND3X1 NAND3X1_96 ( .A(_877_), .B(_879_), .C(_878_), .Y(_880_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_874_) );
AND2X2 AND2X2_96 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_875_) );
OAI21X1 OAI21X1_256 ( .A(_874_), .B(_875_), .C(_72__3_), .Y(_876_) );
NAND2X1 NAND2X1_257 ( .A(_876_), .B(_880_), .Y(_70__3_) );
OAI21X1 OAI21X1_257 ( .A(_877_), .B(_874_), .C(_879_), .Y(_68_) );
INVX1 INVX1_162 ( .A(1'b0), .Y(_884_) );
OR2X2 OR2X2_97 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_885_) );
NAND2X1 NAND2X1_258 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_886_) );
NAND3X1 NAND3X1_97 ( .A(_884_), .B(_886_), .C(_885_), .Y(_887_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_881_) );
AND2X2 AND2X2_97 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_882_) );
OAI21X1 OAI21X1_258 ( .A(_881_), .B(_882_), .C(1'b0), .Y(_883_) );
NAND2X1 NAND2X1_259 ( .A(_883_), .B(_887_), .Y(_75__0_) );
OAI21X1 OAI21X1_259 ( .A(_884_), .B(_881_), .C(_886_), .Y(_77__1_) );
INVX1 INVX1_163 ( .A(_77__1_), .Y(_891_) );
OR2X2 OR2X2_98 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_892_) );
NAND2X1 NAND2X1_260 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_893_) );
NAND3X1 NAND3X1_98 ( .A(_891_), .B(_893_), .C(_892_), .Y(_894_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_888_) );
AND2X2 AND2X2_98 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_889_) );
OAI21X1 OAI21X1_260 ( .A(_888_), .B(_889_), .C(_77__1_), .Y(_890_) );
NAND2X1 NAND2X1_261 ( .A(_890_), .B(_894_), .Y(_75__1_) );
OAI21X1 OAI21X1_261 ( .A(_891_), .B(_888_), .C(_893_), .Y(_77__2_) );
INVX1 INVX1_164 ( .A(_77__2_), .Y(_898_) );
OR2X2 OR2X2_99 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_899_) );
NAND2X1 NAND2X1_262 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_900_) );
NAND3X1 NAND3X1_99 ( .A(_898_), .B(_900_), .C(_899_), .Y(_901_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_895_) );
AND2X2 AND2X2_99 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_896_) );
OAI21X1 OAI21X1_262 ( .A(_895_), .B(_896_), .C(_77__2_), .Y(_897_) );
NAND2X1 NAND2X1_263 ( .A(_897_), .B(_901_), .Y(_75__2_) );
OAI21X1 OAI21X1_263 ( .A(_898_), .B(_895_), .C(_900_), .Y(_77__3_) );
INVX1 INVX1_165 ( .A(_77__3_), .Y(_905_) );
OR2X2 OR2X2_100 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_906_) );
NAND2X1 NAND2X1_264 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_907_) );
NAND3X1 NAND3X1_100 ( .A(_905_), .B(_907_), .C(_906_), .Y(_908_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_902_) );
AND2X2 AND2X2_100 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_903_) );
OAI21X1 OAI21X1_264 ( .A(_902_), .B(_903_), .C(_77__3_), .Y(_904_) );
NAND2X1 NAND2X1_265 ( .A(_904_), .B(_908_), .Y(_75__3_) );
OAI21X1 OAI21X1_265 ( .A(_905_), .B(_902_), .C(_907_), .Y(_73_) );
INVX1 INVX1_166 ( .A(1'b1), .Y(_912_) );
OR2X2 OR2X2_101 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_913_) );
NAND2X1 NAND2X1_266 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_914_) );
NAND3X1 NAND3X1_101 ( .A(_912_), .B(_914_), .C(_913_), .Y(_915_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_909_) );
AND2X2 AND2X2_101 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_910_) );
OAI21X1 OAI21X1_266 ( .A(_909_), .B(_910_), .C(1'b1), .Y(_911_) );
NAND2X1 NAND2X1_267 ( .A(_911_), .B(_915_), .Y(_76__0_) );
OAI21X1 OAI21X1_267 ( .A(_912_), .B(_909_), .C(_914_), .Y(_78__1_) );
INVX1 INVX1_167 ( .A(_78__1_), .Y(_919_) );
OR2X2 OR2X2_102 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_920_) );
NAND2X1 NAND2X1_268 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_921_) );
NAND3X1 NAND3X1_102 ( .A(_919_), .B(_921_), .C(_920_), .Y(_922_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_916_) );
AND2X2 AND2X2_102 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_917_) );
OAI21X1 OAI21X1_268 ( .A(_916_), .B(_917_), .C(_78__1_), .Y(_918_) );
NAND2X1 NAND2X1_269 ( .A(_918_), .B(_922_), .Y(_76__1_) );
OAI21X1 OAI21X1_269 ( .A(_919_), .B(_916_), .C(_921_), .Y(_78__2_) );
INVX1 INVX1_168 ( .A(_78__2_), .Y(_926_) );
OR2X2 OR2X2_103 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_927_) );
NAND2X1 NAND2X1_270 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_928_) );
NAND3X1 NAND3X1_103 ( .A(_926_), .B(_928_), .C(_927_), .Y(_929_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_923_) );
AND2X2 AND2X2_103 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_924_) );
OAI21X1 OAI21X1_270 ( .A(_923_), .B(_924_), .C(_78__2_), .Y(_925_) );
NAND2X1 NAND2X1_271 ( .A(_925_), .B(_929_), .Y(_76__2_) );
OAI21X1 OAI21X1_271 ( .A(_926_), .B(_923_), .C(_928_), .Y(_78__3_) );
INVX1 INVX1_169 ( .A(_78__3_), .Y(_933_) );
OR2X2 OR2X2_104 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_934_) );
NAND2X1 NAND2X1_272 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_935_) );
NAND3X1 NAND3X1_104 ( .A(_933_), .B(_935_), .C(_934_), .Y(_936_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_930_) );
AND2X2 AND2X2_104 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_931_) );
OAI21X1 OAI21X1_272 ( .A(_930_), .B(_931_), .C(_78__3_), .Y(_932_) );
NAND2X1 NAND2X1_273 ( .A(_932_), .B(_936_), .Y(_76__3_) );
OAI21X1 OAI21X1_273 ( .A(_933_), .B(_930_), .C(_935_), .Y(_74_) );
INVX1 INVX1_170 ( .A(1'b0), .Y(_940_) );
OR2X2 OR2X2_105 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_941_) );
NAND2X1 NAND2X1_274 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_942_) );
NAND3X1 NAND3X1_105 ( .A(_940_), .B(_942_), .C(_941_), .Y(_943_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_937_) );
AND2X2 AND2X2_105 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_938_) );
OAI21X1 OAI21X1_274 ( .A(_937_), .B(_938_), .C(1'b0), .Y(_939_) );
NAND2X1 NAND2X1_275 ( .A(_939_), .B(_943_), .Y(_0__0_) );
OAI21X1 OAI21X1_275 ( .A(_940_), .B(_937_), .C(_942_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_171 ( .A(rca_inst_w_CARRY_1_), .Y(_947_) );
OR2X2 OR2X2_106 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_948_) );
NAND2X1 NAND2X1_276 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_949_) );
NAND3X1 NAND3X1_106 ( .A(_947_), .B(_949_), .C(_948_), .Y(_950_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_944_) );
AND2X2 AND2X2_106 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_945_) );
OAI21X1 OAI21X1_276 ( .A(_944_), .B(_945_), .C(rca_inst_w_CARRY_1_), .Y(_946_) );
NAND2X1 NAND2X1_277 ( .A(_946_), .B(_950_), .Y(_0__1_) );
OAI21X1 OAI21X1_277 ( .A(_947_), .B(_944_), .C(_949_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_172 ( .A(rca_inst_w_CARRY_2_), .Y(_954_) );
OR2X2 OR2X2_107 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_955_) );
NAND2X1 NAND2X1_278 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_956_) );
NAND3X1 NAND3X1_107 ( .A(_954_), .B(_956_), .C(_955_), .Y(_957_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_951_) );
AND2X2 AND2X2_107 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_952_) );
OAI21X1 OAI21X1_278 ( .A(_951_), .B(_952_), .C(rca_inst_w_CARRY_2_), .Y(_953_) );
NAND2X1 NAND2X1_279 ( .A(_953_), .B(_957_), .Y(_0__2_) );
BUFX2 BUFX2_15 ( .A(w_cout_13_), .Y(cout) );
BUFX2 BUFX2_16 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_17 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_18 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_19 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_20 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_21 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_22 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_23 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_24 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_25 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_26 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_27 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_28 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_29 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_30 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_31 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_32 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_33 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_34 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_35 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_36 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_37 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_38 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_39 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_40 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_41 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_42 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_43 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_44 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_45 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_46 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_47 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_48 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_49 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_50 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_51 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_52 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_53 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_54 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_55 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_56 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_57 ( .A(1'b0), .Y(_5__0_) );
BUFX2 BUFX2_58 ( .A(_1_), .Y(_5__4_) );
BUFX2 BUFX2_59 ( .A(1'b1), .Y(_6__0_) );
BUFX2 BUFX2_60 ( .A(_2_), .Y(_6__4_) );
BUFX2 BUFX2_61 ( .A(1'b0), .Y(_11__0_) );
BUFX2 BUFX2_62 ( .A(_7_), .Y(_11__4_) );
BUFX2 BUFX2_63 ( .A(1'b1), .Y(_12__0_) );
BUFX2 BUFX2_64 ( .A(_8_), .Y(_12__4_) );
BUFX2 BUFX2_65 ( .A(1'b0), .Y(_17__0_) );
BUFX2 BUFX2_66 ( .A(_13_), .Y(_17__4_) );
BUFX2 BUFX2_67 ( .A(1'b1), .Y(_18__0_) );
BUFX2 BUFX2_68 ( .A(_14_), .Y(_18__4_) );
BUFX2 BUFX2_69 ( .A(1'b0), .Y(_23__0_) );
BUFX2 BUFX2_70 ( .A(_19_), .Y(_23__4_) );
BUFX2 BUFX2_71 ( .A(1'b1), .Y(_24__0_) );
BUFX2 BUFX2_72 ( .A(_20_), .Y(_24__4_) );
BUFX2 BUFX2_73 ( .A(1'b0), .Y(_29__0_) );
BUFX2 BUFX2_74 ( .A(_25_), .Y(_29__4_) );
BUFX2 BUFX2_75 ( .A(1'b1), .Y(_30__0_) );
BUFX2 BUFX2_76 ( .A(_26_), .Y(_30__4_) );
BUFX2 BUFX2_77 ( .A(1'b0), .Y(_35__0_) );
BUFX2 BUFX2_78 ( .A(_31_), .Y(_35__4_) );
BUFX2 BUFX2_79 ( .A(1'b1), .Y(_36__0_) );
BUFX2 BUFX2_80 ( .A(_32_), .Y(_36__4_) );
BUFX2 BUFX2_81 ( .A(1'b0), .Y(_41__0_) );
BUFX2 BUFX2_82 ( .A(_37_), .Y(_41__4_) );
BUFX2 BUFX2_83 ( .A(1'b1), .Y(_42__0_) );
BUFX2 BUFX2_84 ( .A(_38_), .Y(_42__4_) );
BUFX2 BUFX2_85 ( .A(1'b0), .Y(_47__0_) );
BUFX2 BUFX2_86 ( .A(_43_), .Y(_47__4_) );
BUFX2 BUFX2_87 ( .A(1'b1), .Y(_48__0_) );
BUFX2 BUFX2_88 ( .A(_44_), .Y(_48__4_) );
BUFX2 BUFX2_89 ( .A(1'b0), .Y(_53__0_) );
BUFX2 BUFX2_90 ( .A(_49_), .Y(_53__4_) );
BUFX2 BUFX2_91 ( .A(1'b1), .Y(_54__0_) );
BUFX2 BUFX2_92 ( .A(_50_), .Y(_54__4_) );
BUFX2 BUFX2_93 ( .A(1'b0), .Y(_59__0_) );
BUFX2 BUFX2_94 ( .A(_55_), .Y(_59__4_) );
BUFX2 BUFX2_95 ( .A(1'b1), .Y(_60__0_) );
BUFX2 BUFX2_96 ( .A(_56_), .Y(_60__4_) );
BUFX2 BUFX2_97 ( .A(1'b0), .Y(_65__0_) );
BUFX2 BUFX2_98 ( .A(_61_), .Y(_65__4_) );
BUFX2 BUFX2_99 ( .A(1'b1), .Y(_66__0_) );
BUFX2 BUFX2_100 ( .A(_62_), .Y(_66__4_) );
BUFX2 BUFX2_101 ( .A(1'b0), .Y(_71__0_) );
BUFX2 BUFX2_102 ( .A(_67_), .Y(_71__4_) );
BUFX2 BUFX2_103 ( .A(1'b1), .Y(_72__0_) );
BUFX2 BUFX2_104 ( .A(_68_), .Y(_72__4_) );
BUFX2 BUFX2_105 ( .A(1'b0), .Y(_77__0_) );
BUFX2 BUFX2_106 ( .A(_73_), .Y(_77__4_) );
BUFX2 BUFX2_107 ( .A(1'b1), .Y(_78__0_) );
BUFX2 BUFX2_108 ( .A(_74_), .Y(_78__4_) );
BUFX2 BUFX2_109 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_110 ( .A(1'b0), .Y(w_cout_0_) );
endmodule
