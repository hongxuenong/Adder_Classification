module CSkipA_42bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output cout;

NAND3X1 NAND3X1_1 ( .A(_407_), .B(_409_), .C(_408_), .Y(_410_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_404_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_405_) );
OAI21X1 OAI21X1_1 ( .A(_404_), .B(_405_), .C(_26__2_), .Y(_406_) );
NAND2X1 NAND2X1_1 ( .A(_406_), .B(_410_), .Y(_0__34_) );
OAI21X1 OAI21X1_2 ( .A(_407_), .B(_404_), .C(_409_), .Y(_26__3_) );
INVX1 INVX1_1 ( .A(i_add_term1[32]), .Y(_411_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[32]), .B(_411_), .Y(_412_) );
INVX1 INVX1_2 ( .A(i_add_term2[32]), .Y(_413_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term1[32]), .B(_413_), .Y(_414_) );
INVX1 INVX1_3 ( .A(i_add_term1[33]), .Y(_415_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[33]), .B(_415_), .Y(_416_) );
INVX1 INVX1_4 ( .A(i_add_term2[33]), .Y(_417_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term1[33]), .B(_417_), .Y(_418_) );
OAI22X1 OAI22X1_1 ( .A(_412_), .B(_414_), .C(_416_), .D(_418_), .Y(_419_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_420_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_421_) );
NOR2X1 NOR2X1_7 ( .A(_420_), .B(_421_), .Y(_422_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_423_) );
NAND2X1 NAND2X1_2 ( .A(_422_), .B(_423_), .Y(_424_) );
NOR2X1 NOR2X1_8 ( .A(_419_), .B(_424_), .Y(_27_) );
INVX1 INVX1_5 ( .A(_25_), .Y(_425_) );
NAND2X1 NAND2X1_3 ( .A(1'b0), .B(_27_), .Y(_426_) );
OAI21X1 OAI21X1_3 ( .A(_27_), .B(_425_), .C(_426_), .Y(w_cout_9_) );
INVX1 INVX1_6 ( .A(w_cout_9_), .Y(_430_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_431_) );
NAND2X1 NAND2X1_4 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_432_) );
NAND3X1 NAND3X1_2 ( .A(_430_), .B(_432_), .C(_431_), .Y(_433_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_427_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_428_) );
OAI21X1 OAI21X1_4 ( .A(_427_), .B(_428_), .C(w_cout_9_), .Y(_429_) );
NAND2X1 NAND2X1_5 ( .A(_429_), .B(_433_), .Y(_0__36_) );
OAI21X1 OAI21X1_5 ( .A(_430_), .B(_427_), .C(_432_), .Y(_29__1_) );
INVX1 INVX1_7 ( .A(_29__3_), .Y(_437_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_438_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_439_) );
NAND3X1 NAND3X1_3 ( .A(_437_), .B(_439_), .C(_438_), .Y(_440_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_434_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_435_) );
OAI21X1 OAI21X1_6 ( .A(_434_), .B(_435_), .C(_29__3_), .Y(_436_) );
NAND2X1 NAND2X1_7 ( .A(_436_), .B(_440_), .Y(_0__39_) );
OAI21X1 OAI21X1_7 ( .A(_437_), .B(_434_), .C(_439_), .Y(_28_) );
INVX1 INVX1_8 ( .A(_29__1_), .Y(_444_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_445_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_446_) );
NAND3X1 NAND3X1_4 ( .A(_444_), .B(_446_), .C(_445_), .Y(_447_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_441_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_442_) );
OAI21X1 OAI21X1_8 ( .A(_441_), .B(_442_), .C(_29__1_), .Y(_443_) );
NAND2X1 NAND2X1_9 ( .A(_443_), .B(_447_), .Y(_0__37_) );
OAI21X1 OAI21X1_9 ( .A(_444_), .B(_441_), .C(_446_), .Y(_29__2_) );
INVX1 INVX1_9 ( .A(_29__2_), .Y(_451_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_452_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_453_) );
NAND3X1 NAND3X1_5 ( .A(_451_), .B(_453_), .C(_452_), .Y(_454_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_448_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_449_) );
OAI21X1 OAI21X1_10 ( .A(_448_), .B(_449_), .C(_29__2_), .Y(_450_) );
NAND2X1 NAND2X1_11 ( .A(_450_), .B(_454_), .Y(_0__38_) );
OAI21X1 OAI21X1_11 ( .A(_451_), .B(_448_), .C(_453_), .Y(_29__3_) );
INVX1 INVX1_10 ( .A(i_add_term1[36]), .Y(_455_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[36]), .B(_455_), .Y(_456_) );
INVX1 INVX1_11 ( .A(i_add_term2[36]), .Y(_457_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term1[36]), .B(_457_), .Y(_458_) );
INVX1 INVX1_12 ( .A(i_add_term1[37]), .Y(_459_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[37]), .B(_459_), .Y(_460_) );
INVX1 INVX1_13 ( .A(i_add_term2[37]), .Y(_461_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term1[37]), .B(_461_), .Y(_462_) );
OAI22X1 OAI22X1_2 ( .A(_456_), .B(_458_), .C(_460_), .D(_462_), .Y(_463_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_464_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_465_) );
NOR2X1 NOR2X1_18 ( .A(_464_), .B(_465_), .Y(_466_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_467_) );
NAND2X1 NAND2X1_12 ( .A(_466_), .B(_467_), .Y(_468_) );
NOR2X1 NOR2X1_19 ( .A(_463_), .B(_468_), .Y(_30_) );
INVX1 INVX1_14 ( .A(_28_), .Y(_469_) );
NAND2X1 NAND2X1_13 ( .A(1'b0), .B(_30_), .Y(_470_) );
OAI21X1 OAI21X1_12 ( .A(_30_), .B(_469_), .C(_470_), .Y(cskip2_inst_cin) );
INVX1 INVX1_15 ( .A(cskip2_inst_cin), .Y(_474_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_475_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_476_) );
NAND3X1 NAND3X1_6 ( .A(_474_), .B(_476_), .C(_475_), .Y(_477_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_471_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_472_) );
OAI21X1 OAI21X1_13 ( .A(_471_), .B(_472_), .C(cskip2_inst_cin), .Y(_473_) );
NAND2X1 NAND2X1_15 ( .A(_473_), .B(_477_), .Y(cskip2_inst_rca0_fa0_o_sum) );
OAI21X1 OAI21X1_14 ( .A(_474_), .B(_471_), .C(_476_), .Y(cskip2_inst_rca0_c) );
INVX1 INVX1_16 ( .A(cskip2_inst_rca0_c), .Y(_481_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_482_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_483_) );
NAND3X1 NAND3X1_7 ( .A(_481_), .B(_483_), .C(_482_), .Y(_484_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_478_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_479_) );
OAI21X1 OAI21X1_15 ( .A(_478_), .B(_479_), .C(cskip2_inst_rca0_c), .Y(_480_) );
NAND2X1 NAND2X1_17 ( .A(_480_), .B(_484_), .Y(cskip2_inst_rca0_fa31_o_sum) );
OAI21X1 OAI21X1_16 ( .A(_481_), .B(_478_), .C(_483_), .Y(cskip2_inst_cout0) );
INVX1 INVX1_17 ( .A(i_add_term1[41]), .Y(_489_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[41]), .B(_489_), .Y(_490_) );
INVX1 INVX1_18 ( .A(i_add_term2[41]), .Y(_491_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term1[41]), .B(_491_), .Y(_492_) );
INVX1 INVX1_19 ( .A(i_add_term1[40]), .Y(_485_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[40]), .B(_485_), .Y(_486_) );
INVX1 INVX1_20 ( .A(i_add_term2[40]), .Y(_487_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term1[40]), .B(_487_), .Y(_488_) );
AOI22X1 AOI22X1_1 ( .A(_490_), .B(_492_), .C(_486_), .D(_488_), .Y(cskip2_inst_skip0_P) );
INVX1 INVX1_21 ( .A(cskip2_inst_cout0), .Y(_493_) );
NAND2X1 NAND2X1_22 ( .A(1'b0), .B(cskip2_inst_skip0_P), .Y(_494_) );
OAI21X1 OAI21X1_17 ( .A(cskip2_inst_skip0_P), .B(_493_), .C(_494_), .Y(w_cout_11_) );
BUFX2 BUFX2_1 ( .A(w_cout_11_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(cskip2_inst_rca0_fa0_o_sum), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(cskip2_inst_rca0_fa31_o_sum), .Y(sum[41]) );
INVX1 INVX1_22 ( .A(1'b0), .Y(_34_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_35_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_36_) );
NAND3X1 NAND3X1_8 ( .A(_34_), .B(_36_), .C(_35_), .Y(_37_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_31_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_32_) );
OAI21X1 OAI21X1_18 ( .A(_31_), .B(_32_), .C(1'b0), .Y(_33_) );
NAND2X1 NAND2X1_24 ( .A(_33_), .B(_37_), .Y(_0__0_) );
OAI21X1 OAI21X1_19 ( .A(_34_), .B(_31_), .C(_36_), .Y(_2__1_) );
INVX1 INVX1_23 ( .A(_2__3_), .Y(_41_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_42_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_43_) );
NAND3X1 NAND3X1_9 ( .A(_41_), .B(_43_), .C(_42_), .Y(_44_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_38_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_39_) );
OAI21X1 OAI21X1_20 ( .A(_38_), .B(_39_), .C(_2__3_), .Y(_40_) );
NAND2X1 NAND2X1_26 ( .A(_40_), .B(_44_), .Y(_0__3_) );
OAI21X1 OAI21X1_21 ( .A(_41_), .B(_38_), .C(_43_), .Y(_1_) );
INVX1 INVX1_24 ( .A(_2__1_), .Y(_48_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_49_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_50_) );
NAND3X1 NAND3X1_10 ( .A(_48_), .B(_50_), .C(_49_), .Y(_51_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_45_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_46_) );
OAI21X1 OAI21X1_22 ( .A(_45_), .B(_46_), .C(_2__1_), .Y(_47_) );
NAND2X1 NAND2X1_28 ( .A(_47_), .B(_51_), .Y(_0__1_) );
OAI21X1 OAI21X1_23 ( .A(_48_), .B(_45_), .C(_50_), .Y(_2__2_) );
INVX1 INVX1_25 ( .A(_2__2_), .Y(_55_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_56_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_57_) );
NAND3X1 NAND3X1_11 ( .A(_55_), .B(_57_), .C(_56_), .Y(_58_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_52_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_53_) );
OAI21X1 OAI21X1_24 ( .A(_52_), .B(_53_), .C(_2__2_), .Y(_54_) );
NAND2X1 NAND2X1_30 ( .A(_54_), .B(_58_), .Y(_0__2_) );
OAI21X1 OAI21X1_25 ( .A(_55_), .B(_52_), .C(_57_), .Y(_2__3_) );
INVX1 INVX1_26 ( .A(i_add_term1[0]), .Y(_59_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[0]), .B(_59_), .Y(_60_) );
INVX1 INVX1_27 ( .A(i_add_term2[0]), .Y(_61_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term1[0]), .B(_61_), .Y(_62_) );
INVX1 INVX1_28 ( .A(i_add_term1[1]), .Y(_63_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[1]), .B(_63_), .Y(_64_) );
INVX1 INVX1_29 ( .A(i_add_term2[1]), .Y(_65_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term1[1]), .B(_65_), .Y(_66_) );
OAI22X1 OAI22X1_3 ( .A(_60_), .B(_62_), .C(_64_), .D(_66_), .Y(_67_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_68_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_69_) );
NOR2X1 NOR2X1_31 ( .A(_68_), .B(_69_), .Y(_70_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_71_) );
NAND2X1 NAND2X1_31 ( .A(_70_), .B(_71_), .Y(_72_) );
NOR2X1 NOR2X1_32 ( .A(_67_), .B(_72_), .Y(_3_) );
INVX1 INVX1_30 ( .A(_1_), .Y(_73_) );
NAND2X1 NAND2X1_32 ( .A(1'b0), .B(_3_), .Y(_74_) );
OAI21X1 OAI21X1_26 ( .A(_3_), .B(_73_), .C(_74_), .Y(w_cout_1_) );
INVX1 INVX1_31 ( .A(w_cout_1_), .Y(_78_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_79_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_80_) );
NAND3X1 NAND3X1_12 ( .A(_78_), .B(_80_), .C(_79_), .Y(_81_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_75_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_76_) );
OAI21X1 OAI21X1_27 ( .A(_75_), .B(_76_), .C(w_cout_1_), .Y(_77_) );
NAND2X1 NAND2X1_34 ( .A(_77_), .B(_81_), .Y(_0__4_) );
OAI21X1 OAI21X1_28 ( .A(_78_), .B(_75_), .C(_80_), .Y(_5__1_) );
INVX1 INVX1_32 ( .A(_5__3_), .Y(_85_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_86_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_87_) );
NAND3X1 NAND3X1_13 ( .A(_85_), .B(_87_), .C(_86_), .Y(_88_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_82_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_83_) );
OAI21X1 OAI21X1_29 ( .A(_82_), .B(_83_), .C(_5__3_), .Y(_84_) );
NAND2X1 NAND2X1_36 ( .A(_84_), .B(_88_), .Y(_0__7_) );
OAI21X1 OAI21X1_30 ( .A(_85_), .B(_82_), .C(_87_), .Y(_4_) );
INVX1 INVX1_33 ( .A(_5__1_), .Y(_92_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_93_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_94_) );
NAND3X1 NAND3X1_14 ( .A(_92_), .B(_94_), .C(_93_), .Y(_95_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_89_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_90_) );
OAI21X1 OAI21X1_31 ( .A(_89_), .B(_90_), .C(_5__1_), .Y(_91_) );
NAND2X1 NAND2X1_38 ( .A(_91_), .B(_95_), .Y(_0__5_) );
OAI21X1 OAI21X1_32 ( .A(_92_), .B(_89_), .C(_94_), .Y(_5__2_) );
INVX1 INVX1_34 ( .A(_5__2_), .Y(_99_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_100_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_101_) );
NAND3X1 NAND3X1_15 ( .A(_99_), .B(_101_), .C(_100_), .Y(_102_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_96_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_97_) );
OAI21X1 OAI21X1_33 ( .A(_96_), .B(_97_), .C(_5__2_), .Y(_98_) );
NAND2X1 NAND2X1_40 ( .A(_98_), .B(_102_), .Y(_0__6_) );
OAI21X1 OAI21X1_34 ( .A(_99_), .B(_96_), .C(_101_), .Y(_5__3_) );
INVX1 INVX1_35 ( .A(i_add_term1[4]), .Y(_103_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[4]), .B(_103_), .Y(_104_) );
INVX1 INVX1_36 ( .A(i_add_term2[4]), .Y(_105_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term1[4]), .B(_105_), .Y(_106_) );
INVX1 INVX1_37 ( .A(i_add_term1[5]), .Y(_107_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[5]), .B(_107_), .Y(_108_) );
INVX1 INVX1_38 ( .A(i_add_term2[5]), .Y(_109_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term1[5]), .B(_109_), .Y(_110_) );
OAI22X1 OAI22X1_4 ( .A(_104_), .B(_106_), .C(_108_), .D(_110_), .Y(_111_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_112_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_113_) );
NOR2X1 NOR2X1_42 ( .A(_112_), .B(_113_), .Y(_114_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_115_) );
NAND2X1 NAND2X1_41 ( .A(_114_), .B(_115_), .Y(_116_) );
NOR2X1 NOR2X1_43 ( .A(_111_), .B(_116_), .Y(_6_) );
INVX1 INVX1_39 ( .A(_4_), .Y(_117_) );
NAND2X1 NAND2X1_42 ( .A(1'b0), .B(_6_), .Y(_118_) );
OAI21X1 OAI21X1_35 ( .A(_6_), .B(_117_), .C(_118_), .Y(w_cout_2_) );
INVX1 INVX1_40 ( .A(w_cout_2_), .Y(_122_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_123_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_124_) );
NAND3X1 NAND3X1_16 ( .A(_122_), .B(_124_), .C(_123_), .Y(_125_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_119_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_120_) );
OAI21X1 OAI21X1_36 ( .A(_119_), .B(_120_), .C(w_cout_2_), .Y(_121_) );
NAND2X1 NAND2X1_44 ( .A(_121_), .B(_125_), .Y(_0__8_) );
OAI21X1 OAI21X1_37 ( .A(_122_), .B(_119_), .C(_124_), .Y(_8__1_) );
INVX1 INVX1_41 ( .A(_8__3_), .Y(_129_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_130_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_131_) );
NAND3X1 NAND3X1_17 ( .A(_129_), .B(_131_), .C(_130_), .Y(_132_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_126_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_127_) );
OAI21X1 OAI21X1_38 ( .A(_126_), .B(_127_), .C(_8__3_), .Y(_128_) );
NAND2X1 NAND2X1_46 ( .A(_128_), .B(_132_), .Y(_0__11_) );
OAI21X1 OAI21X1_39 ( .A(_129_), .B(_126_), .C(_131_), .Y(_7_) );
INVX1 INVX1_42 ( .A(_8__1_), .Y(_136_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_137_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_138_) );
NAND3X1 NAND3X1_18 ( .A(_136_), .B(_138_), .C(_137_), .Y(_139_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_133_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_134_) );
OAI21X1 OAI21X1_40 ( .A(_133_), .B(_134_), .C(_8__1_), .Y(_135_) );
NAND2X1 NAND2X1_48 ( .A(_135_), .B(_139_), .Y(_0__9_) );
OAI21X1 OAI21X1_41 ( .A(_136_), .B(_133_), .C(_138_), .Y(_8__2_) );
INVX1 INVX1_43 ( .A(_8__2_), .Y(_143_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_144_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_145_) );
NAND3X1 NAND3X1_19 ( .A(_143_), .B(_145_), .C(_144_), .Y(_146_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_140_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_141_) );
OAI21X1 OAI21X1_42 ( .A(_140_), .B(_141_), .C(_8__2_), .Y(_142_) );
NAND2X1 NAND2X1_50 ( .A(_142_), .B(_146_), .Y(_0__10_) );
OAI21X1 OAI21X1_43 ( .A(_143_), .B(_140_), .C(_145_), .Y(_8__3_) );
INVX1 INVX1_44 ( .A(i_add_term1[8]), .Y(_147_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[8]), .B(_147_), .Y(_148_) );
INVX1 INVX1_45 ( .A(i_add_term2[8]), .Y(_149_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term1[8]), .B(_149_), .Y(_150_) );
INVX1 INVX1_46 ( .A(i_add_term1[9]), .Y(_151_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[9]), .B(_151_), .Y(_152_) );
INVX1 INVX1_47 ( .A(i_add_term2[9]), .Y(_153_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term1[9]), .B(_153_), .Y(_154_) );
OAI22X1 OAI22X1_5 ( .A(_148_), .B(_150_), .C(_152_), .D(_154_), .Y(_155_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_156_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_157_) );
NOR2X1 NOR2X1_53 ( .A(_156_), .B(_157_), .Y(_158_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_159_) );
NAND2X1 NAND2X1_51 ( .A(_158_), .B(_159_), .Y(_160_) );
NOR2X1 NOR2X1_54 ( .A(_155_), .B(_160_), .Y(_9_) );
INVX1 INVX1_48 ( .A(_7_), .Y(_161_) );
NAND2X1 NAND2X1_52 ( .A(1'b0), .B(_9_), .Y(_162_) );
OAI21X1 OAI21X1_44 ( .A(_9_), .B(_161_), .C(_162_), .Y(w_cout_3_) );
INVX1 INVX1_49 ( .A(w_cout_3_), .Y(_166_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_167_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_168_) );
NAND3X1 NAND3X1_20 ( .A(_166_), .B(_168_), .C(_167_), .Y(_169_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_163_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_164_) );
OAI21X1 OAI21X1_45 ( .A(_163_), .B(_164_), .C(w_cout_3_), .Y(_165_) );
NAND2X1 NAND2X1_54 ( .A(_165_), .B(_169_), .Y(_0__12_) );
OAI21X1 OAI21X1_46 ( .A(_166_), .B(_163_), .C(_168_), .Y(_11__1_) );
INVX1 INVX1_50 ( .A(_11__3_), .Y(_173_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_174_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_175_) );
NAND3X1 NAND3X1_21 ( .A(_173_), .B(_175_), .C(_174_), .Y(_176_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_170_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_171_) );
OAI21X1 OAI21X1_47 ( .A(_170_), .B(_171_), .C(_11__3_), .Y(_172_) );
NAND2X1 NAND2X1_56 ( .A(_172_), .B(_176_), .Y(_0__15_) );
OAI21X1 OAI21X1_48 ( .A(_173_), .B(_170_), .C(_175_), .Y(_10_) );
INVX1 INVX1_51 ( .A(_11__1_), .Y(_180_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_181_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_182_) );
NAND3X1 NAND3X1_22 ( .A(_180_), .B(_182_), .C(_181_), .Y(_183_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_177_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_178_) );
OAI21X1 OAI21X1_49 ( .A(_177_), .B(_178_), .C(_11__1_), .Y(_179_) );
NAND2X1 NAND2X1_58 ( .A(_179_), .B(_183_), .Y(_0__13_) );
OAI21X1 OAI21X1_50 ( .A(_180_), .B(_177_), .C(_182_), .Y(_11__2_) );
INVX1 INVX1_52 ( .A(_11__2_), .Y(_187_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_188_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_189_) );
NAND3X1 NAND3X1_23 ( .A(_187_), .B(_189_), .C(_188_), .Y(_190_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_184_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_185_) );
OAI21X1 OAI21X1_51 ( .A(_184_), .B(_185_), .C(_11__2_), .Y(_186_) );
NAND2X1 NAND2X1_60 ( .A(_186_), .B(_190_), .Y(_0__14_) );
OAI21X1 OAI21X1_52 ( .A(_187_), .B(_184_), .C(_189_), .Y(_11__3_) );
INVX1 INVX1_53 ( .A(i_add_term1[12]), .Y(_191_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[12]), .B(_191_), .Y(_192_) );
INVX1 INVX1_54 ( .A(i_add_term2[12]), .Y(_193_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term1[12]), .B(_193_), .Y(_194_) );
INVX1 INVX1_55 ( .A(i_add_term1[13]), .Y(_195_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[13]), .B(_195_), .Y(_196_) );
INVX1 INVX1_56 ( .A(i_add_term2[13]), .Y(_197_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term1[13]), .B(_197_), .Y(_198_) );
OAI22X1 OAI22X1_6 ( .A(_192_), .B(_194_), .C(_196_), .D(_198_), .Y(_199_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_200_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_201_) );
NOR2X1 NOR2X1_64 ( .A(_200_), .B(_201_), .Y(_202_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_203_) );
NAND2X1 NAND2X1_61 ( .A(_202_), .B(_203_), .Y(_204_) );
NOR2X1 NOR2X1_65 ( .A(_199_), .B(_204_), .Y(_12_) );
INVX1 INVX1_57 ( .A(_10_), .Y(_205_) );
NAND2X1 NAND2X1_62 ( .A(1'b0), .B(_12_), .Y(_206_) );
OAI21X1 OAI21X1_53 ( .A(_12_), .B(_205_), .C(_206_), .Y(w_cout_4_) );
INVX1 INVX1_58 ( .A(w_cout_4_), .Y(_210_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_211_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_212_) );
NAND3X1 NAND3X1_24 ( .A(_210_), .B(_212_), .C(_211_), .Y(_213_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_207_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_208_) );
OAI21X1 OAI21X1_54 ( .A(_207_), .B(_208_), .C(w_cout_4_), .Y(_209_) );
NAND2X1 NAND2X1_64 ( .A(_209_), .B(_213_), .Y(_0__16_) );
OAI21X1 OAI21X1_55 ( .A(_210_), .B(_207_), .C(_212_), .Y(_14__1_) );
INVX1 INVX1_59 ( .A(_14__3_), .Y(_217_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_218_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_219_) );
NAND3X1 NAND3X1_25 ( .A(_217_), .B(_219_), .C(_218_), .Y(_220_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_214_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_215_) );
OAI21X1 OAI21X1_56 ( .A(_214_), .B(_215_), .C(_14__3_), .Y(_216_) );
NAND2X1 NAND2X1_66 ( .A(_216_), .B(_220_), .Y(_0__19_) );
OAI21X1 OAI21X1_57 ( .A(_217_), .B(_214_), .C(_219_), .Y(_13_) );
INVX1 INVX1_60 ( .A(_14__1_), .Y(_224_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_225_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_226_) );
NAND3X1 NAND3X1_26 ( .A(_224_), .B(_226_), .C(_225_), .Y(_227_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_221_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_222_) );
OAI21X1 OAI21X1_58 ( .A(_221_), .B(_222_), .C(_14__1_), .Y(_223_) );
NAND2X1 NAND2X1_68 ( .A(_223_), .B(_227_), .Y(_0__17_) );
OAI21X1 OAI21X1_59 ( .A(_224_), .B(_221_), .C(_226_), .Y(_14__2_) );
INVX1 INVX1_61 ( .A(_14__2_), .Y(_231_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_232_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_233_) );
NAND3X1 NAND3X1_27 ( .A(_231_), .B(_233_), .C(_232_), .Y(_234_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_228_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_229_) );
OAI21X1 OAI21X1_60 ( .A(_228_), .B(_229_), .C(_14__2_), .Y(_230_) );
NAND2X1 NAND2X1_70 ( .A(_230_), .B(_234_), .Y(_0__18_) );
OAI21X1 OAI21X1_61 ( .A(_231_), .B(_228_), .C(_233_), .Y(_14__3_) );
INVX1 INVX1_62 ( .A(i_add_term1[16]), .Y(_235_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[16]), .B(_235_), .Y(_236_) );
INVX1 INVX1_63 ( .A(i_add_term2[16]), .Y(_237_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term1[16]), .B(_237_), .Y(_238_) );
INVX1 INVX1_64 ( .A(i_add_term1[17]), .Y(_239_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[17]), .B(_239_), .Y(_240_) );
INVX1 INVX1_65 ( .A(i_add_term2[17]), .Y(_241_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term1[17]), .B(_241_), .Y(_242_) );
OAI22X1 OAI22X1_7 ( .A(_236_), .B(_238_), .C(_240_), .D(_242_), .Y(_243_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_244_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_245_) );
NOR2X1 NOR2X1_75 ( .A(_244_), .B(_245_), .Y(_246_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_247_) );
NAND2X1 NAND2X1_71 ( .A(_246_), .B(_247_), .Y(_248_) );
NOR2X1 NOR2X1_76 ( .A(_243_), .B(_248_), .Y(_15_) );
INVX1 INVX1_66 ( .A(_13_), .Y(_249_) );
NAND2X1 NAND2X1_72 ( .A(1'b0), .B(_15_), .Y(_250_) );
OAI21X1 OAI21X1_62 ( .A(_15_), .B(_249_), .C(_250_), .Y(w_cout_5_) );
INVX1 INVX1_67 ( .A(w_cout_5_), .Y(_254_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_255_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_256_) );
NAND3X1 NAND3X1_28 ( .A(_254_), .B(_256_), .C(_255_), .Y(_257_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_251_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_252_) );
OAI21X1 OAI21X1_63 ( .A(_251_), .B(_252_), .C(w_cout_5_), .Y(_253_) );
NAND2X1 NAND2X1_74 ( .A(_253_), .B(_257_), .Y(_0__20_) );
OAI21X1 OAI21X1_64 ( .A(_254_), .B(_251_), .C(_256_), .Y(_17__1_) );
INVX1 INVX1_68 ( .A(_17__3_), .Y(_261_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_262_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_263_) );
NAND3X1 NAND3X1_29 ( .A(_261_), .B(_263_), .C(_262_), .Y(_264_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_258_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_259_) );
OAI21X1 OAI21X1_65 ( .A(_258_), .B(_259_), .C(_17__3_), .Y(_260_) );
NAND2X1 NAND2X1_76 ( .A(_260_), .B(_264_), .Y(_0__23_) );
OAI21X1 OAI21X1_66 ( .A(_261_), .B(_258_), .C(_263_), .Y(_16_) );
INVX1 INVX1_69 ( .A(_17__1_), .Y(_268_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_269_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_270_) );
NAND3X1 NAND3X1_30 ( .A(_268_), .B(_270_), .C(_269_), .Y(_271_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_265_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_266_) );
OAI21X1 OAI21X1_67 ( .A(_265_), .B(_266_), .C(_17__1_), .Y(_267_) );
NAND2X1 NAND2X1_78 ( .A(_267_), .B(_271_), .Y(_0__21_) );
OAI21X1 OAI21X1_68 ( .A(_268_), .B(_265_), .C(_270_), .Y(_17__2_) );
INVX1 INVX1_70 ( .A(_17__2_), .Y(_275_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_276_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_277_) );
NAND3X1 NAND3X1_31 ( .A(_275_), .B(_277_), .C(_276_), .Y(_278_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_272_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_273_) );
OAI21X1 OAI21X1_69 ( .A(_272_), .B(_273_), .C(_17__2_), .Y(_274_) );
NAND2X1 NAND2X1_80 ( .A(_274_), .B(_278_), .Y(_0__22_) );
OAI21X1 OAI21X1_70 ( .A(_275_), .B(_272_), .C(_277_), .Y(_17__3_) );
INVX1 INVX1_71 ( .A(i_add_term1[20]), .Y(_279_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[20]), .B(_279_), .Y(_280_) );
INVX1 INVX1_72 ( .A(i_add_term2[20]), .Y(_281_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term1[20]), .B(_281_), .Y(_282_) );
INVX1 INVX1_73 ( .A(i_add_term1[21]), .Y(_283_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[21]), .B(_283_), .Y(_284_) );
INVX1 INVX1_74 ( .A(i_add_term2[21]), .Y(_285_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term1[21]), .B(_285_), .Y(_286_) );
OAI22X1 OAI22X1_8 ( .A(_280_), .B(_282_), .C(_284_), .D(_286_), .Y(_287_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_288_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_289_) );
NOR2X1 NOR2X1_86 ( .A(_288_), .B(_289_), .Y(_290_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_291_) );
NAND2X1 NAND2X1_81 ( .A(_290_), .B(_291_), .Y(_292_) );
NOR2X1 NOR2X1_87 ( .A(_287_), .B(_292_), .Y(_18_) );
INVX1 INVX1_75 ( .A(_16_), .Y(_293_) );
NAND2X1 NAND2X1_82 ( .A(1'b0), .B(_18_), .Y(_294_) );
OAI21X1 OAI21X1_71 ( .A(_18_), .B(_293_), .C(_294_), .Y(w_cout_6_) );
INVX1 INVX1_76 ( .A(w_cout_6_), .Y(_298_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_299_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_300_) );
NAND3X1 NAND3X1_32 ( .A(_298_), .B(_300_), .C(_299_), .Y(_301_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_295_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_296_) );
OAI21X1 OAI21X1_72 ( .A(_295_), .B(_296_), .C(w_cout_6_), .Y(_297_) );
NAND2X1 NAND2X1_84 ( .A(_297_), .B(_301_), .Y(_0__24_) );
OAI21X1 OAI21X1_73 ( .A(_298_), .B(_295_), .C(_300_), .Y(_20__1_) );
INVX1 INVX1_77 ( .A(_20__3_), .Y(_305_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_306_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_307_) );
NAND3X1 NAND3X1_33 ( .A(_305_), .B(_307_), .C(_306_), .Y(_308_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_302_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_303_) );
OAI21X1 OAI21X1_74 ( .A(_302_), .B(_303_), .C(_20__3_), .Y(_304_) );
NAND2X1 NAND2X1_86 ( .A(_304_), .B(_308_), .Y(_0__27_) );
OAI21X1 OAI21X1_75 ( .A(_305_), .B(_302_), .C(_307_), .Y(_19_) );
INVX1 INVX1_78 ( .A(_20__1_), .Y(_312_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_313_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_314_) );
NAND3X1 NAND3X1_34 ( .A(_312_), .B(_314_), .C(_313_), .Y(_315_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_309_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_310_) );
OAI21X1 OAI21X1_76 ( .A(_309_), .B(_310_), .C(_20__1_), .Y(_311_) );
NAND2X1 NAND2X1_88 ( .A(_311_), .B(_315_), .Y(_0__25_) );
OAI21X1 OAI21X1_77 ( .A(_312_), .B(_309_), .C(_314_), .Y(_20__2_) );
INVX1 INVX1_79 ( .A(_20__2_), .Y(_319_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_320_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_321_) );
NAND3X1 NAND3X1_35 ( .A(_319_), .B(_321_), .C(_320_), .Y(_322_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_316_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_317_) );
OAI21X1 OAI21X1_78 ( .A(_316_), .B(_317_), .C(_20__2_), .Y(_318_) );
NAND2X1 NAND2X1_90 ( .A(_318_), .B(_322_), .Y(_0__26_) );
OAI21X1 OAI21X1_79 ( .A(_319_), .B(_316_), .C(_321_), .Y(_20__3_) );
INVX1 INVX1_80 ( .A(i_add_term1[24]), .Y(_323_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[24]), .B(_323_), .Y(_324_) );
INVX1 INVX1_81 ( .A(i_add_term2[24]), .Y(_325_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term1[24]), .B(_325_), .Y(_326_) );
INVX1 INVX1_82 ( .A(i_add_term1[25]), .Y(_327_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[25]), .B(_327_), .Y(_328_) );
INVX1 INVX1_83 ( .A(i_add_term2[25]), .Y(_329_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term1[25]), .B(_329_), .Y(_330_) );
OAI22X1 OAI22X1_9 ( .A(_324_), .B(_326_), .C(_328_), .D(_330_), .Y(_331_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_332_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_333_) );
NOR2X1 NOR2X1_97 ( .A(_332_), .B(_333_), .Y(_334_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_335_) );
NAND2X1 NAND2X1_91 ( .A(_334_), .B(_335_), .Y(_336_) );
NOR2X1 NOR2X1_98 ( .A(_331_), .B(_336_), .Y(_21_) );
INVX1 INVX1_84 ( .A(_19_), .Y(_337_) );
NAND2X1 NAND2X1_92 ( .A(1'b0), .B(_21_), .Y(_338_) );
OAI21X1 OAI21X1_80 ( .A(_21_), .B(_337_), .C(_338_), .Y(w_cout_7_) );
INVX1 INVX1_85 ( .A(w_cout_7_), .Y(_342_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_343_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_344_) );
NAND3X1 NAND3X1_36 ( .A(_342_), .B(_344_), .C(_343_), .Y(_345_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_339_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_340_) );
OAI21X1 OAI21X1_81 ( .A(_339_), .B(_340_), .C(w_cout_7_), .Y(_341_) );
NAND2X1 NAND2X1_94 ( .A(_341_), .B(_345_), .Y(_0__28_) );
OAI21X1 OAI21X1_82 ( .A(_342_), .B(_339_), .C(_344_), .Y(_23__1_) );
INVX1 INVX1_86 ( .A(_23__3_), .Y(_349_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_350_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_351_) );
NAND3X1 NAND3X1_37 ( .A(_349_), .B(_351_), .C(_350_), .Y(_352_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_346_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_347_) );
OAI21X1 OAI21X1_83 ( .A(_346_), .B(_347_), .C(_23__3_), .Y(_348_) );
NAND2X1 NAND2X1_96 ( .A(_348_), .B(_352_), .Y(_0__31_) );
OAI21X1 OAI21X1_84 ( .A(_349_), .B(_346_), .C(_351_), .Y(_22_) );
INVX1 INVX1_87 ( .A(_23__1_), .Y(_356_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_357_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_358_) );
NAND3X1 NAND3X1_38 ( .A(_356_), .B(_358_), .C(_357_), .Y(_359_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_353_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_354_) );
OAI21X1 OAI21X1_85 ( .A(_353_), .B(_354_), .C(_23__1_), .Y(_355_) );
NAND2X1 NAND2X1_98 ( .A(_355_), .B(_359_), .Y(_0__29_) );
OAI21X1 OAI21X1_86 ( .A(_356_), .B(_353_), .C(_358_), .Y(_23__2_) );
INVX1 INVX1_88 ( .A(_23__2_), .Y(_363_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_364_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_365_) );
NAND3X1 NAND3X1_39 ( .A(_363_), .B(_365_), .C(_364_), .Y(_366_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_360_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_361_) );
OAI21X1 OAI21X1_87 ( .A(_360_), .B(_361_), .C(_23__2_), .Y(_362_) );
NAND2X1 NAND2X1_100 ( .A(_362_), .B(_366_), .Y(_0__30_) );
OAI21X1 OAI21X1_88 ( .A(_363_), .B(_360_), .C(_365_), .Y(_23__3_) );
INVX1 INVX1_89 ( .A(i_add_term1[28]), .Y(_367_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[28]), .B(_367_), .Y(_368_) );
INVX1 INVX1_90 ( .A(i_add_term2[28]), .Y(_369_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term1[28]), .B(_369_), .Y(_370_) );
INVX1 INVX1_91 ( .A(i_add_term1[29]), .Y(_371_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[29]), .B(_371_), .Y(_372_) );
INVX1 INVX1_92 ( .A(i_add_term2[29]), .Y(_373_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term1[29]), .B(_373_), .Y(_374_) );
OAI22X1 OAI22X1_10 ( .A(_368_), .B(_370_), .C(_372_), .D(_374_), .Y(_375_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_376_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_377_) );
NOR2X1 NOR2X1_108 ( .A(_376_), .B(_377_), .Y(_378_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_379_) );
NAND2X1 NAND2X1_101 ( .A(_378_), .B(_379_), .Y(_380_) );
NOR2X1 NOR2X1_109 ( .A(_375_), .B(_380_), .Y(_24_) );
INVX1 INVX1_93 ( .A(_22_), .Y(_381_) );
NAND2X1 NAND2X1_102 ( .A(1'b0), .B(_24_), .Y(_382_) );
OAI21X1 OAI21X1_89 ( .A(_24_), .B(_381_), .C(_382_), .Y(w_cout_8_) );
INVX1 INVX1_94 ( .A(w_cout_8_), .Y(_386_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_387_) );
NAND2X1 NAND2X1_103 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_388_) );
NAND3X1 NAND3X1_40 ( .A(_386_), .B(_388_), .C(_387_), .Y(_389_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_383_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_384_) );
OAI21X1 OAI21X1_90 ( .A(_383_), .B(_384_), .C(w_cout_8_), .Y(_385_) );
NAND2X1 NAND2X1_104 ( .A(_385_), .B(_389_), .Y(_0__32_) );
OAI21X1 OAI21X1_91 ( .A(_386_), .B(_383_), .C(_388_), .Y(_26__1_) );
INVX1 INVX1_95 ( .A(_26__3_), .Y(_393_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_394_) );
NAND2X1 NAND2X1_105 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_395_) );
NAND3X1 NAND3X1_41 ( .A(_393_), .B(_395_), .C(_394_), .Y(_396_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_390_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_391_) );
OAI21X1 OAI21X1_92 ( .A(_390_), .B(_391_), .C(_26__3_), .Y(_392_) );
NAND2X1 NAND2X1_106 ( .A(_392_), .B(_396_), .Y(_0__35_) );
OAI21X1 OAI21X1_93 ( .A(_393_), .B(_390_), .C(_395_), .Y(_25_) );
INVX1 INVX1_96 ( .A(_26__1_), .Y(_400_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_401_) );
NAND2X1 NAND2X1_107 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_402_) );
NAND3X1 NAND3X1_42 ( .A(_400_), .B(_402_), .C(_401_), .Y(_403_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_397_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_398_) );
OAI21X1 OAI21X1_94 ( .A(_397_), .B(_398_), .C(_26__1_), .Y(_399_) );
NAND2X1 NAND2X1_108 ( .A(_399_), .B(_403_), .Y(_0__33_) );
OAI21X1 OAI21X1_95 ( .A(_400_), .B(_397_), .C(_402_), .Y(_26__2_) );
INVX1 INVX1_97 ( .A(_26__2_), .Y(_407_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_408_) );
NAND2X1 NAND2X1_109 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_409_) );
BUFX2 BUFX2_44 ( .A(cskip2_inst_rca0_fa0_o_sum), .Y(_0__40_) );
BUFX2 BUFX2_45 ( .A(cskip2_inst_rca0_fa31_o_sum), .Y(_0__41_) );
BUFX2 BUFX2_46 ( .A(1'b0), .Y(w_cout_0_) );
BUFX2 BUFX2_47 ( .A(cskip2_inst_cin), .Y(w_cout_10_) );
endmodule
