module cla_5bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [4:0] i_add1;
input [4:0] i_add2;
output [5:0] o_result;

OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_40_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_41_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_41_), .C(_40_), .Y(_42_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_36_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_37_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_37_), .C(w_C_2_), .Y(_38_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_42_), .Y(_14__2_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_46_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_47_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_48_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_48_), .C(_47_), .Y(_49_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_43_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_44_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_44_), .C(w_C_3_), .Y(_45_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_49_), .Y(_14__3_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_1_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_2_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_3_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_4_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_4_), .Y(_5_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(_3_), .C(_5_), .Y(_6_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_6_), .Y(w_C_3_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_7_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_8_), .C(_6_), .Y(_9_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_7_), .Y(w_C_4_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_10_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_11_), .C(_9_), .Y(_12_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_12_), .Y(w_C_5_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .C(_5_), .Y(_13_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(w_C_2_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_14__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_14__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_14__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_14__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_14__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(o_result[5]) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_18_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_19_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_20_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_20_), .C(_19_), .Y(_21_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_15_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_16_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_16_), .C(w_C_4_), .Y(_17_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_21_), .Y(_14__4_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_25_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_26_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_27_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_27_), .C(_26_), .Y(_28_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_22_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_23_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_23_), .C(gnd), .Y(_24_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_28_), .Y(_14__0_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_32_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_33_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_34_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_34_), .C(_33_), .Y(_35_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_29_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_30_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_30_), .C(w_C_1_), .Y(_31_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_35_), .Y(_14__1_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_39_) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_14__5_) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
