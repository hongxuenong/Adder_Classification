module cla_36bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add1[19], i_add1[20], i_add1[21], i_add1[22], i_add1[23], i_add1[24], i_add1[25], i_add1[26], i_add1[27], i_add1[28], i_add1[29], i_add1[30], i_add1[31], i_add1[32], i_add1[33], i_add1[34], i_add1[35], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], i_add2[19], i_add2[20], i_add2[21], i_add2[22], i_add2[23], i_add2[24], i_add2[25], i_add2[26], i_add2[27], i_add2[28], i_add2[29], i_add2[30], i_add2[31], i_add2[32], i_add2[33], i_add2[34], i_add2[35], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21], o_result[22], o_result[23], o_result[24], o_result[25], o_result[26], o_result[27], o_result[28], o_result[29], o_result[30], o_result[31], o_result[32], o_result[33], o_result[34], o_result[35], o_result[36]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add1[19];
input i_add1[20];
input i_add1[21];
input i_add1[22];
input i_add1[23];
input i_add1[24];
input i_add1[25];
input i_add1[26];
input i_add1[27];
input i_add1[28];
input i_add1[29];
input i_add1[30];
input i_add1[31];
input i_add1[32];
input i_add1[33];
input i_add1[34];
input i_add1[35];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
input i_add2[19];
input i_add2[20];
input i_add2[21];
input i_add2[22];
input i_add2[23];
input i_add2[24];
input i_add2[25];
input i_add2[26];
input i_add2[27];
input i_add2[28];
input i_add2[29];
input i_add2[30];
input i_add2[31];
input i_add2[32];
input i_add2[33];
input i_add2[34];
input i_add2[35];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];
output o_result[22];
output o_result[23];
output o_result[24];
output o_result[25];
output o_result[26];
output o_result[27];
output o_result[28];
output o_result[29];
output o_result[30];
output o_result[31];
output o_result[32];
output o_result[33];
output o_result[34];
output o_result[35];
output o_result[36];

INVX1 INVX1_1 ( .A(w_C_3_), .Y(_446_) );
OR2X2 OR2X2_1 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_447_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_448_) );
NAND3X1 NAND3X1_1 ( .A(_446_), .B(_448_), .C(_447_), .Y(_449_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_443_) );
AND2X2 AND2X2_1 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_444_) );
OAI21X1 OAI21X1_1 ( .A(_443_), .B(_444_), .C(w_C_3_), .Y(_445_) );
NAND2X1 NAND2X1_2 ( .A(_445_), .B(_449_), .Y(_197__3_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_2 ( .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_3 ( .A(_1_), .B(_2_), .Y(w_C_2_) );
INVX1 INVX1_3 ( .A(i_add2[2]), .Y(_3_) );
INVX1 INVX1_4 ( .A(i_add1[2]), .Y(_4_) );
NAND2X1 NAND2X1_4 ( .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
OAI21X1 OAI21X1_2 ( .A(_1_), .B(_2_), .C(_6_), .Y(_7_) );
AND2X2 AND2X2_2 ( .A(_7_), .B(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
OR2X2 OR2X2_2 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_2 ( .A(_5_), .B(_9_), .C(_7_), .Y(_10_) );
NAND2X1 NAND2X1_7 ( .A(_8_), .B(_10_), .Y(w_C_4_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
INVX1 INVX1_5 ( .A(_11_), .Y(_12_) );
NAND2X1 NAND2X1_8 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
NAND3X1 NAND3X1_3 ( .A(_8_), .B(_13_), .C(_10_), .Y(_14_) );
AND2X2 AND2X2_3 ( .A(_14_), .B(_12_), .Y(w_C_5_) );
AND2X2 AND2X2_4 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_15_) );
INVX1 INVX1_6 ( .A(_15_), .Y(_16_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_17_) );
INVX1 INVX1_7 ( .A(_17_), .Y(_18_) );
NAND3X1 NAND3X1_4 ( .A(_12_), .B(_18_), .C(_14_), .Y(_19_) );
AND2X2 AND2X2_5 ( .A(_19_), .B(_16_), .Y(_20_) );
INVX1 INVX1_8 ( .A(_20_), .Y(w_C_6_) );
AND2X2 AND2X2_6 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_21_) );
INVX1 INVX1_9 ( .A(_21_), .Y(_22_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_23_) );
OAI21X1 OAI21X1_3 ( .A(_23_), .B(_20_), .C(_22_), .Y(w_C_7_) );
AND2X2 AND2X2_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_24_) );
INVX1 INVX1_10 ( .A(_24_), .Y(_25_) );
INVX1 INVX1_11 ( .A(_23_), .Y(_26_) );
NAND3X1 NAND3X1_5 ( .A(_16_), .B(_22_), .C(_19_), .Y(_27_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_28_) );
INVX1 INVX1_12 ( .A(_28_), .Y(_29_) );
NAND3X1 NAND3X1_6 ( .A(_26_), .B(_29_), .C(_27_), .Y(_30_) );
AND2X2 AND2X2_8 ( .A(_30_), .B(_25_), .Y(_31_) );
INVX1 INVX1_13 ( .A(_31_), .Y(w_C_8_) );
AND2X2 AND2X2_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_32_) );
INVX1 INVX1_14 ( .A(_32_), .Y(_33_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_34_) );
OAI21X1 OAI21X1_4 ( .A(_34_), .B(_31_), .C(_33_), .Y(w_C_9_) );
INVX1 INVX1_15 ( .A(i_add2[9]), .Y(_35_) );
INVX1 INVX1_16 ( .A(i_add1[9]), .Y(_36_) );
INVX1 INVX1_17 ( .A(_34_), .Y(_37_) );
NAND3X1 NAND3X1_7 ( .A(_25_), .B(_33_), .C(_30_), .Y(_38_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_39_) );
INVX1 INVX1_18 ( .A(_39_), .Y(_40_) );
NAND3X1 NAND3X1_8 ( .A(_37_), .B(_40_), .C(_38_), .Y(_41_) );
OAI21X1 OAI21X1_5 ( .A(_35_), .B(_36_), .C(_41_), .Y(w_C_10_) );
NOR2X1 NOR2X1_10 ( .A(_35_), .B(_36_), .Y(_42_) );
INVX1 INVX1_19 ( .A(_42_), .Y(_43_) );
AND2X2 AND2X2_10 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_44_) );
INVX1 INVX1_20 ( .A(_44_), .Y(_45_) );
NAND3X1 NAND3X1_9 ( .A(_43_), .B(_45_), .C(_41_), .Y(_46_) );
OAI21X1 OAI21X1_6 ( .A(i_add2[10]), .B(i_add1[10]), .C(_46_), .Y(_47_) );
INVX1 INVX1_21 ( .A(_47_), .Y(w_C_11_) );
INVX1 INVX1_22 ( .A(i_add2[11]), .Y(_48_) );
INVX1 INVX1_23 ( .A(i_add1[11]), .Y(_49_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_50_) );
INVX1 INVX1_24 ( .A(_50_), .Y(_51_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_52_) );
INVX1 INVX1_25 ( .A(_52_), .Y(_53_) );
NAND3X1 NAND3X1_10 ( .A(_51_), .B(_53_), .C(_46_), .Y(_54_) );
OAI21X1 OAI21X1_7 ( .A(_48_), .B(_49_), .C(_54_), .Y(w_C_12_) );
NOR2X1 NOR2X1_13 ( .A(_48_), .B(_49_), .Y(_55_) );
INVX1 INVX1_26 ( .A(_55_), .Y(_56_) );
AND2X2 AND2X2_11 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_57_) );
INVX1 INVX1_27 ( .A(_57_), .Y(_58_) );
NAND3X1 NAND3X1_11 ( .A(_56_), .B(_58_), .C(_54_), .Y(_59_) );
OAI21X1 OAI21X1_8 ( .A(i_add2[12]), .B(i_add1[12]), .C(_59_), .Y(_60_) );
INVX1 INVX1_28 ( .A(_60_), .Y(w_C_13_) );
INVX1 INVX1_29 ( .A(i_add2[13]), .Y(_61_) );
INVX1 INVX1_30 ( .A(i_add1[13]), .Y(_62_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_63_) );
INVX1 INVX1_31 ( .A(_63_), .Y(_64_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_65_) );
INVX1 INVX1_32 ( .A(_65_), .Y(_66_) );
NAND3X1 NAND3X1_12 ( .A(_64_), .B(_66_), .C(_59_), .Y(_67_) );
OAI21X1 OAI21X1_9 ( .A(_61_), .B(_62_), .C(_67_), .Y(w_C_14_) );
NOR2X1 NOR2X1_16 ( .A(_61_), .B(_62_), .Y(_68_) );
INVX1 INVX1_33 ( .A(_68_), .Y(_69_) );
AND2X2 AND2X2_12 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_70_) );
INVX1 INVX1_34 ( .A(_70_), .Y(_71_) );
NAND3X1 NAND3X1_13 ( .A(_69_), .B(_71_), .C(_67_), .Y(_72_) );
OAI21X1 OAI21X1_10 ( .A(i_add2[14]), .B(i_add1[14]), .C(_72_), .Y(_73_) );
INVX1 INVX1_35 ( .A(_73_), .Y(w_C_15_) );
INVX1 INVX1_36 ( .A(i_add2[15]), .Y(_74_) );
INVX1 INVX1_37 ( .A(i_add1[15]), .Y(_75_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_76_) );
INVX1 INVX1_38 ( .A(_76_), .Y(_77_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_78_) );
INVX1 INVX1_39 ( .A(_78_), .Y(_79_) );
NAND3X1 NAND3X1_14 ( .A(_77_), .B(_79_), .C(_72_), .Y(_80_) );
OAI21X1 OAI21X1_11 ( .A(_74_), .B(_75_), .C(_80_), .Y(w_C_16_) );
NOR2X1 NOR2X1_19 ( .A(_74_), .B(_75_), .Y(_81_) );
INVX1 INVX1_40 ( .A(_81_), .Y(_82_) );
AND2X2 AND2X2_13 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_83_) );
INVX1 INVX1_41 ( .A(_83_), .Y(_84_) );
NAND3X1 NAND3X1_15 ( .A(_82_), .B(_84_), .C(_80_), .Y(_85_) );
OAI21X1 OAI21X1_12 ( .A(i_add2[16]), .B(i_add1[16]), .C(_85_), .Y(_86_) );
INVX1 INVX1_42 ( .A(_86_), .Y(w_C_17_) );
INVX1 INVX1_43 ( .A(i_add2[17]), .Y(_87_) );
INVX1 INVX1_44 ( .A(i_add1[17]), .Y(_88_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_89_) );
INVX1 INVX1_45 ( .A(_89_), .Y(_90_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_91_) );
INVX1 INVX1_46 ( .A(_91_), .Y(_92_) );
NAND3X1 NAND3X1_16 ( .A(_90_), .B(_92_), .C(_85_), .Y(_93_) );
OAI21X1 OAI21X1_13 ( .A(_87_), .B(_88_), .C(_93_), .Y(w_C_18_) );
NOR2X1 NOR2X1_22 ( .A(_87_), .B(_88_), .Y(_94_) );
INVX1 INVX1_47 ( .A(_94_), .Y(_95_) );
AND2X2 AND2X2_14 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_96_) );
INVX1 INVX1_48 ( .A(_96_), .Y(_97_) );
NAND3X1 NAND3X1_17 ( .A(_95_), .B(_97_), .C(_93_), .Y(_98_) );
OAI21X1 OAI21X1_14 ( .A(i_add2[18]), .B(i_add1[18]), .C(_98_), .Y(_99_) );
INVX1 INVX1_49 ( .A(_99_), .Y(w_C_19_) );
INVX1 INVX1_50 ( .A(i_add2[19]), .Y(_100_) );
INVX1 INVX1_51 ( .A(i_add1[19]), .Y(_101_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_102_) );
INVX1 INVX1_52 ( .A(_102_), .Y(_103_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_104_) );
INVX1 INVX1_53 ( .A(_104_), .Y(_105_) );
NAND3X1 NAND3X1_18 ( .A(_103_), .B(_105_), .C(_98_), .Y(_106_) );
OAI21X1 OAI21X1_15 ( .A(_100_), .B(_101_), .C(_106_), .Y(w_C_20_) );
NOR2X1 NOR2X1_25 ( .A(_100_), .B(_101_), .Y(_107_) );
INVX1 INVX1_54 ( .A(_107_), .Y(_108_) );
AND2X2 AND2X2_15 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_109_) );
INVX1 INVX1_55 ( .A(_109_), .Y(_110_) );
NAND3X1 NAND3X1_19 ( .A(_108_), .B(_110_), .C(_106_), .Y(_111_) );
OAI21X1 OAI21X1_16 ( .A(i_add2[20]), .B(i_add1[20]), .C(_111_), .Y(_112_) );
INVX1 INVX1_56 ( .A(_112_), .Y(w_C_21_) );
INVX1 INVX1_57 ( .A(i_add2[21]), .Y(_113_) );
INVX1 INVX1_58 ( .A(i_add1[21]), .Y(_114_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_115_) );
INVX1 INVX1_59 ( .A(_115_), .Y(_116_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_117_) );
INVX1 INVX1_60 ( .A(_117_), .Y(_118_) );
NAND3X1 NAND3X1_20 ( .A(_116_), .B(_118_), .C(_111_), .Y(_119_) );
OAI21X1 OAI21X1_17 ( .A(_113_), .B(_114_), .C(_119_), .Y(w_C_22_) );
NOR2X1 NOR2X1_28 ( .A(_113_), .B(_114_), .Y(_120_) );
INVX1 INVX1_61 ( .A(_120_), .Y(_121_) );
AND2X2 AND2X2_16 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_122_) );
INVX1 INVX1_62 ( .A(_122_), .Y(_123_) );
NAND3X1 NAND3X1_21 ( .A(_121_), .B(_123_), .C(_119_), .Y(_124_) );
OAI21X1 OAI21X1_18 ( .A(i_add2[22]), .B(i_add1[22]), .C(_124_), .Y(_125_) );
INVX1 INVX1_63 ( .A(_125_), .Y(w_C_23_) );
INVX1 INVX1_64 ( .A(i_add2[23]), .Y(_126_) );
INVX1 INVX1_65 ( .A(i_add1[23]), .Y(_127_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_128_) );
INVX1 INVX1_66 ( .A(_128_), .Y(_129_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_130_) );
INVX1 INVX1_67 ( .A(_130_), .Y(_131_) );
NAND3X1 NAND3X1_22 ( .A(_129_), .B(_131_), .C(_124_), .Y(_132_) );
OAI21X1 OAI21X1_19 ( .A(_126_), .B(_127_), .C(_132_), .Y(w_C_24_) );
NOR2X1 NOR2X1_31 ( .A(_126_), .B(_127_), .Y(_133_) );
INVX1 INVX1_68 ( .A(_133_), .Y(_134_) );
AND2X2 AND2X2_17 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_135_) );
INVX1 INVX1_69 ( .A(_135_), .Y(_136_) );
NAND3X1 NAND3X1_23 ( .A(_134_), .B(_136_), .C(_132_), .Y(_137_) );
OAI21X1 OAI21X1_20 ( .A(i_add2[24]), .B(i_add1[24]), .C(_137_), .Y(_138_) );
INVX1 INVX1_70 ( .A(_138_), .Y(w_C_25_) );
INVX1 INVX1_71 ( .A(i_add2[25]), .Y(_139_) );
INVX1 INVX1_72 ( .A(i_add1[25]), .Y(_140_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_141_) );
INVX1 INVX1_73 ( .A(_141_), .Y(_142_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_143_) );
INVX1 INVX1_74 ( .A(_143_), .Y(_144_) );
NAND3X1 NAND3X1_24 ( .A(_142_), .B(_144_), .C(_137_), .Y(_145_) );
OAI21X1 OAI21X1_21 ( .A(_139_), .B(_140_), .C(_145_), .Y(w_C_26_) );
NOR2X1 NOR2X1_34 ( .A(_139_), .B(_140_), .Y(_146_) );
INVX1 INVX1_75 ( .A(_146_), .Y(_147_) );
AND2X2 AND2X2_18 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_148_) );
INVX1 INVX1_76 ( .A(_148_), .Y(_149_) );
NAND3X1 NAND3X1_25 ( .A(_147_), .B(_149_), .C(_145_), .Y(_150_) );
OAI21X1 OAI21X1_22 ( .A(i_add2[26]), .B(i_add1[26]), .C(_150_), .Y(_151_) );
INVX1 INVX1_77 ( .A(_151_), .Y(w_C_27_) );
INVX1 INVX1_78 ( .A(i_add2[27]), .Y(_152_) );
INVX1 INVX1_79 ( .A(i_add1[27]), .Y(_153_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_154_) );
INVX1 INVX1_80 ( .A(_154_), .Y(_155_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_156_) );
INVX1 INVX1_81 ( .A(_156_), .Y(_157_) );
NAND3X1 NAND3X1_26 ( .A(_155_), .B(_157_), .C(_150_), .Y(_158_) );
OAI21X1 OAI21X1_23 ( .A(_152_), .B(_153_), .C(_158_), .Y(w_C_28_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_159_) );
INVX1 INVX1_82 ( .A(_159_), .Y(_160_) );
NOR2X1 NOR2X1_38 ( .A(_152_), .B(_153_), .Y(_161_) );
INVX1 INVX1_83 ( .A(_161_), .Y(_162_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_163_) );
NAND3X1 NAND3X1_27 ( .A(_162_), .B(_163_), .C(_158_), .Y(_164_) );
AND2X2 AND2X2_19 ( .A(_164_), .B(_160_), .Y(w_C_29_) );
INVX1 INVX1_84 ( .A(i_add2[29]), .Y(_165_) );
INVX1 INVX1_85 ( .A(i_add1[29]), .Y(_166_) );
NAND2X1 NAND2X1_10 ( .A(_165_), .B(_166_), .Y(_167_) );
NAND3X1 NAND3X1_28 ( .A(_160_), .B(_167_), .C(_164_), .Y(_168_) );
OAI21X1 OAI21X1_24 ( .A(_165_), .B(_166_), .C(_168_), .Y(w_C_30_) );
INVX1 INVX1_86 ( .A(i_add2[30]), .Y(_169_) );
INVX1 INVX1_87 ( .A(i_add1[30]), .Y(_170_) );
NAND2X1 NAND2X1_11 ( .A(_169_), .B(_170_), .Y(_171_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_172_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_173_) );
NAND3X1 NAND3X1_29 ( .A(_172_), .B(_173_), .C(_168_), .Y(_174_) );
AND2X2 AND2X2_20 ( .A(_174_), .B(_171_), .Y(w_C_31_) );
INVX1 INVX1_88 ( .A(i_add2[31]), .Y(_175_) );
INVX1 INVX1_89 ( .A(i_add1[31]), .Y(_176_) );
NAND2X1 NAND2X1_14 ( .A(_175_), .B(_176_), .Y(_177_) );
NAND3X1 NAND3X1_30 ( .A(_171_), .B(_177_), .C(_174_), .Y(_178_) );
OAI21X1 OAI21X1_25 ( .A(_175_), .B(_176_), .C(_178_), .Y(w_C_32_) );
NOR2X1 NOR2X1_39 ( .A(_175_), .B(_176_), .Y(_179_) );
INVX1 INVX1_90 ( .A(_179_), .Y(_180_) );
AND2X2 AND2X2_21 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_181_) );
INVX1 INVX1_91 ( .A(_181_), .Y(_182_) );
NAND3X1 NAND3X1_31 ( .A(_180_), .B(_182_), .C(_178_), .Y(_183_) );
OAI21X1 OAI21X1_26 ( .A(i_add2[32]), .B(i_add1[32]), .C(_183_), .Y(_184_) );
INVX1 INVX1_92 ( .A(_184_), .Y(w_C_33_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_185_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_186_) );
OAI21X1 OAI21X1_27 ( .A(_186_), .B(_184_), .C(_185_), .Y(w_C_34_) );
OR2X2 OR2X2_3 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_187_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_188_) );
INVX1 INVX1_93 ( .A(_188_), .Y(_189_) );
INVX1 INVX1_94 ( .A(_186_), .Y(_190_) );
NAND3X1 NAND3X1_32 ( .A(_189_), .B(_190_), .C(_183_), .Y(_191_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_192_) );
NAND3X1 NAND3X1_33 ( .A(_185_), .B(_192_), .C(_191_), .Y(_193_) );
AND2X2 AND2X2_22 ( .A(_193_), .B(_187_), .Y(w_C_35_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_194_) );
OR2X2 OR2X2_4 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_195_) );
NAND3X1 NAND3X1_34 ( .A(_187_), .B(_195_), .C(_193_), .Y(_196_) );
NAND2X1 NAND2X1_18 ( .A(_194_), .B(_196_), .Y(w_C_36_) );
BUFX2 BUFX2_1 ( .A(_197__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_197__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_197__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_197__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_197__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_197__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_197__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_197__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_197__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_197__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_197__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_197__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_197__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_197__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_197__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_197__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_197__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_197__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_197__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_197__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_197__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_197__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_197__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_197__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_197__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_197__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_197__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_197__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_197__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_197__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_197__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_197__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_197__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_197__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_197__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_197__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(w_C_36_), .Y(o_result[36]) );
INVX1 INVX1_95 ( .A(w_C_4_), .Y(_201_) );
OR2X2 OR2X2_5 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_202_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_203_) );
NAND3X1 NAND3X1_35 ( .A(_201_), .B(_203_), .C(_202_), .Y(_204_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_198_) );
AND2X2 AND2X2_23 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_199_) );
OAI21X1 OAI21X1_28 ( .A(_198_), .B(_199_), .C(w_C_4_), .Y(_200_) );
NAND2X1 NAND2X1_20 ( .A(_200_), .B(_204_), .Y(_197__4_) );
INVX1 INVX1_96 ( .A(w_C_5_), .Y(_208_) );
OR2X2 OR2X2_6 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_209_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_210_) );
NAND3X1 NAND3X1_36 ( .A(_208_), .B(_210_), .C(_209_), .Y(_211_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_205_) );
AND2X2 AND2X2_24 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_206_) );
OAI21X1 OAI21X1_29 ( .A(_205_), .B(_206_), .C(w_C_5_), .Y(_207_) );
NAND2X1 NAND2X1_22 ( .A(_207_), .B(_211_), .Y(_197__5_) );
INVX1 INVX1_97 ( .A(w_C_6_), .Y(_215_) );
OR2X2 OR2X2_7 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_216_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_217_) );
NAND3X1 NAND3X1_37 ( .A(_215_), .B(_217_), .C(_216_), .Y(_218_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_212_) );
AND2X2 AND2X2_25 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_213_) );
OAI21X1 OAI21X1_30 ( .A(_212_), .B(_213_), .C(w_C_6_), .Y(_214_) );
NAND2X1 NAND2X1_24 ( .A(_214_), .B(_218_), .Y(_197__6_) );
INVX1 INVX1_98 ( .A(w_C_7_), .Y(_222_) );
OR2X2 OR2X2_8 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_223_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_224_) );
NAND3X1 NAND3X1_38 ( .A(_222_), .B(_224_), .C(_223_), .Y(_225_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_219_) );
AND2X2 AND2X2_26 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_220_) );
OAI21X1 OAI21X1_31 ( .A(_219_), .B(_220_), .C(w_C_7_), .Y(_221_) );
NAND2X1 NAND2X1_26 ( .A(_221_), .B(_225_), .Y(_197__7_) );
INVX1 INVX1_99 ( .A(w_C_8_), .Y(_229_) );
OR2X2 OR2X2_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_230_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_231_) );
NAND3X1 NAND3X1_39 ( .A(_229_), .B(_231_), .C(_230_), .Y(_232_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_226_) );
AND2X2 AND2X2_27 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_227_) );
OAI21X1 OAI21X1_32 ( .A(_226_), .B(_227_), .C(w_C_8_), .Y(_228_) );
NAND2X1 NAND2X1_28 ( .A(_228_), .B(_232_), .Y(_197__8_) );
INVX1 INVX1_100 ( .A(w_C_9_), .Y(_236_) );
OR2X2 OR2X2_10 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_237_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_238_) );
NAND3X1 NAND3X1_40 ( .A(_236_), .B(_238_), .C(_237_), .Y(_239_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_233_) );
AND2X2 AND2X2_28 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_234_) );
OAI21X1 OAI21X1_33 ( .A(_233_), .B(_234_), .C(w_C_9_), .Y(_235_) );
NAND2X1 NAND2X1_30 ( .A(_235_), .B(_239_), .Y(_197__9_) );
INVX1 INVX1_101 ( .A(w_C_10_), .Y(_243_) );
OR2X2 OR2X2_11 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_244_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_245_) );
NAND3X1 NAND3X1_41 ( .A(_243_), .B(_245_), .C(_244_), .Y(_246_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_240_) );
AND2X2 AND2X2_29 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_241_) );
OAI21X1 OAI21X1_34 ( .A(_240_), .B(_241_), .C(w_C_10_), .Y(_242_) );
NAND2X1 NAND2X1_32 ( .A(_242_), .B(_246_), .Y(_197__10_) );
INVX1 INVX1_102 ( .A(w_C_11_), .Y(_250_) );
OR2X2 OR2X2_12 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_251_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_252_) );
NAND3X1 NAND3X1_42 ( .A(_250_), .B(_252_), .C(_251_), .Y(_253_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_247_) );
AND2X2 AND2X2_30 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_248_) );
OAI21X1 OAI21X1_35 ( .A(_247_), .B(_248_), .C(w_C_11_), .Y(_249_) );
NAND2X1 NAND2X1_34 ( .A(_249_), .B(_253_), .Y(_197__11_) );
INVX1 INVX1_103 ( .A(w_C_12_), .Y(_257_) );
OR2X2 OR2X2_13 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_258_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_259_) );
NAND3X1 NAND3X1_43 ( .A(_257_), .B(_259_), .C(_258_), .Y(_260_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_254_) );
AND2X2 AND2X2_31 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_255_) );
OAI21X1 OAI21X1_36 ( .A(_254_), .B(_255_), .C(w_C_12_), .Y(_256_) );
NAND2X1 NAND2X1_36 ( .A(_256_), .B(_260_), .Y(_197__12_) );
INVX1 INVX1_104 ( .A(w_C_13_), .Y(_264_) );
OR2X2 OR2X2_14 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_265_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_266_) );
NAND3X1 NAND3X1_44 ( .A(_264_), .B(_266_), .C(_265_), .Y(_267_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_261_) );
AND2X2 AND2X2_32 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_262_) );
OAI21X1 OAI21X1_37 ( .A(_261_), .B(_262_), .C(w_C_13_), .Y(_263_) );
NAND2X1 NAND2X1_38 ( .A(_263_), .B(_267_), .Y(_197__13_) );
INVX1 INVX1_105 ( .A(w_C_14_), .Y(_271_) );
OR2X2 OR2X2_15 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_272_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_273_) );
NAND3X1 NAND3X1_45 ( .A(_271_), .B(_273_), .C(_272_), .Y(_274_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_268_) );
AND2X2 AND2X2_33 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_269_) );
OAI21X1 OAI21X1_38 ( .A(_268_), .B(_269_), .C(w_C_14_), .Y(_270_) );
NAND2X1 NAND2X1_40 ( .A(_270_), .B(_274_), .Y(_197__14_) );
INVX1 INVX1_106 ( .A(w_C_15_), .Y(_278_) );
OR2X2 OR2X2_16 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_279_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_280_) );
NAND3X1 NAND3X1_46 ( .A(_278_), .B(_280_), .C(_279_), .Y(_281_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_275_) );
AND2X2 AND2X2_34 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_276_) );
OAI21X1 OAI21X1_39 ( .A(_275_), .B(_276_), .C(w_C_15_), .Y(_277_) );
NAND2X1 NAND2X1_42 ( .A(_277_), .B(_281_), .Y(_197__15_) );
INVX1 INVX1_107 ( .A(w_C_16_), .Y(_285_) );
OR2X2 OR2X2_17 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_286_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_287_) );
NAND3X1 NAND3X1_47 ( .A(_285_), .B(_287_), .C(_286_), .Y(_288_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_282_) );
AND2X2 AND2X2_35 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_283_) );
OAI21X1 OAI21X1_40 ( .A(_282_), .B(_283_), .C(w_C_16_), .Y(_284_) );
NAND2X1 NAND2X1_44 ( .A(_284_), .B(_288_), .Y(_197__16_) );
INVX1 INVX1_108 ( .A(w_C_17_), .Y(_292_) );
OR2X2 OR2X2_18 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_293_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_294_) );
NAND3X1 NAND3X1_48 ( .A(_292_), .B(_294_), .C(_293_), .Y(_295_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_289_) );
AND2X2 AND2X2_36 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_290_) );
OAI21X1 OAI21X1_41 ( .A(_289_), .B(_290_), .C(w_C_17_), .Y(_291_) );
NAND2X1 NAND2X1_46 ( .A(_291_), .B(_295_), .Y(_197__17_) );
INVX1 INVX1_109 ( .A(w_C_18_), .Y(_299_) );
OR2X2 OR2X2_19 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_300_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_301_) );
NAND3X1 NAND3X1_49 ( .A(_299_), .B(_301_), .C(_300_), .Y(_302_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_296_) );
AND2X2 AND2X2_37 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_297_) );
OAI21X1 OAI21X1_42 ( .A(_296_), .B(_297_), .C(w_C_18_), .Y(_298_) );
NAND2X1 NAND2X1_48 ( .A(_298_), .B(_302_), .Y(_197__18_) );
INVX1 INVX1_110 ( .A(w_C_19_), .Y(_306_) );
OR2X2 OR2X2_20 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_307_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_308_) );
NAND3X1 NAND3X1_50 ( .A(_306_), .B(_308_), .C(_307_), .Y(_309_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_303_) );
AND2X2 AND2X2_38 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_304_) );
OAI21X1 OAI21X1_43 ( .A(_303_), .B(_304_), .C(w_C_19_), .Y(_305_) );
NAND2X1 NAND2X1_50 ( .A(_305_), .B(_309_), .Y(_197__19_) );
INVX1 INVX1_111 ( .A(w_C_20_), .Y(_313_) );
OR2X2 OR2X2_21 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_314_) );
NAND2X1 NAND2X1_51 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_315_) );
NAND3X1 NAND3X1_51 ( .A(_313_), .B(_315_), .C(_314_), .Y(_316_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_310_) );
AND2X2 AND2X2_39 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_311_) );
OAI21X1 OAI21X1_44 ( .A(_310_), .B(_311_), .C(w_C_20_), .Y(_312_) );
NAND2X1 NAND2X1_52 ( .A(_312_), .B(_316_), .Y(_197__20_) );
INVX1 INVX1_112 ( .A(w_C_21_), .Y(_320_) );
OR2X2 OR2X2_22 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_321_) );
NAND2X1 NAND2X1_53 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_322_) );
NAND3X1 NAND3X1_52 ( .A(_320_), .B(_322_), .C(_321_), .Y(_323_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_317_) );
AND2X2 AND2X2_40 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_318_) );
OAI21X1 OAI21X1_45 ( .A(_317_), .B(_318_), .C(w_C_21_), .Y(_319_) );
NAND2X1 NAND2X1_54 ( .A(_319_), .B(_323_), .Y(_197__21_) );
INVX1 INVX1_113 ( .A(w_C_22_), .Y(_327_) );
OR2X2 OR2X2_23 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_328_) );
NAND2X1 NAND2X1_55 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_329_) );
NAND3X1 NAND3X1_53 ( .A(_327_), .B(_329_), .C(_328_), .Y(_330_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_324_) );
AND2X2 AND2X2_41 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_325_) );
OAI21X1 OAI21X1_46 ( .A(_324_), .B(_325_), .C(w_C_22_), .Y(_326_) );
NAND2X1 NAND2X1_56 ( .A(_326_), .B(_330_), .Y(_197__22_) );
INVX1 INVX1_114 ( .A(w_C_23_), .Y(_334_) );
OR2X2 OR2X2_24 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_335_) );
NAND2X1 NAND2X1_57 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_336_) );
NAND3X1 NAND3X1_54 ( .A(_334_), .B(_336_), .C(_335_), .Y(_337_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_331_) );
AND2X2 AND2X2_42 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_332_) );
OAI21X1 OAI21X1_47 ( .A(_331_), .B(_332_), .C(w_C_23_), .Y(_333_) );
NAND2X1 NAND2X1_58 ( .A(_333_), .B(_337_), .Y(_197__23_) );
INVX1 INVX1_115 ( .A(w_C_24_), .Y(_341_) );
OR2X2 OR2X2_25 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_342_) );
NAND2X1 NAND2X1_59 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_343_) );
NAND3X1 NAND3X1_55 ( .A(_341_), .B(_343_), .C(_342_), .Y(_344_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_338_) );
AND2X2 AND2X2_43 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_339_) );
OAI21X1 OAI21X1_48 ( .A(_338_), .B(_339_), .C(w_C_24_), .Y(_340_) );
NAND2X1 NAND2X1_60 ( .A(_340_), .B(_344_), .Y(_197__24_) );
INVX1 INVX1_116 ( .A(w_C_25_), .Y(_348_) );
OR2X2 OR2X2_26 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_349_) );
NAND2X1 NAND2X1_61 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_350_) );
NAND3X1 NAND3X1_56 ( .A(_348_), .B(_350_), .C(_349_), .Y(_351_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_345_) );
AND2X2 AND2X2_44 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_346_) );
OAI21X1 OAI21X1_49 ( .A(_345_), .B(_346_), .C(w_C_25_), .Y(_347_) );
NAND2X1 NAND2X1_62 ( .A(_347_), .B(_351_), .Y(_197__25_) );
INVX1 INVX1_117 ( .A(w_C_26_), .Y(_355_) );
OR2X2 OR2X2_27 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_356_) );
NAND2X1 NAND2X1_63 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_357_) );
NAND3X1 NAND3X1_57 ( .A(_355_), .B(_357_), .C(_356_), .Y(_358_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_352_) );
AND2X2 AND2X2_45 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_353_) );
OAI21X1 OAI21X1_50 ( .A(_352_), .B(_353_), .C(w_C_26_), .Y(_354_) );
NAND2X1 NAND2X1_64 ( .A(_354_), .B(_358_), .Y(_197__26_) );
INVX1 INVX1_118 ( .A(w_C_27_), .Y(_362_) );
OR2X2 OR2X2_28 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_363_) );
NAND2X1 NAND2X1_65 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_364_) );
NAND3X1 NAND3X1_58 ( .A(_362_), .B(_364_), .C(_363_), .Y(_365_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_359_) );
AND2X2 AND2X2_46 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_360_) );
OAI21X1 OAI21X1_51 ( .A(_359_), .B(_360_), .C(w_C_27_), .Y(_361_) );
NAND2X1 NAND2X1_66 ( .A(_361_), .B(_365_), .Y(_197__27_) );
INVX1 INVX1_119 ( .A(w_C_28_), .Y(_369_) );
OR2X2 OR2X2_29 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_370_) );
NAND2X1 NAND2X1_67 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_371_) );
NAND3X1 NAND3X1_59 ( .A(_369_), .B(_371_), .C(_370_), .Y(_372_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_366_) );
AND2X2 AND2X2_47 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_367_) );
OAI21X1 OAI21X1_52 ( .A(_366_), .B(_367_), .C(w_C_28_), .Y(_368_) );
NAND2X1 NAND2X1_68 ( .A(_368_), .B(_372_), .Y(_197__28_) );
INVX1 INVX1_120 ( .A(w_C_29_), .Y(_376_) );
OR2X2 OR2X2_30 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_377_) );
NAND2X1 NAND2X1_69 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_378_) );
NAND3X1 NAND3X1_60 ( .A(_376_), .B(_378_), .C(_377_), .Y(_379_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_373_) );
AND2X2 AND2X2_48 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_374_) );
OAI21X1 OAI21X1_53 ( .A(_373_), .B(_374_), .C(w_C_29_), .Y(_375_) );
NAND2X1 NAND2X1_70 ( .A(_375_), .B(_379_), .Y(_197__29_) );
INVX1 INVX1_121 ( .A(w_C_30_), .Y(_383_) );
OR2X2 OR2X2_31 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_384_) );
NAND2X1 NAND2X1_71 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_385_) );
NAND3X1 NAND3X1_61 ( .A(_383_), .B(_385_), .C(_384_), .Y(_386_) );
NOR2X1 NOR2X1_68 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_380_) );
AND2X2 AND2X2_49 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_381_) );
OAI21X1 OAI21X1_54 ( .A(_380_), .B(_381_), .C(w_C_30_), .Y(_382_) );
NAND2X1 NAND2X1_72 ( .A(_382_), .B(_386_), .Y(_197__30_) );
INVX1 INVX1_122 ( .A(w_C_31_), .Y(_390_) );
OR2X2 OR2X2_32 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_391_) );
NAND2X1 NAND2X1_73 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_392_) );
NAND3X1 NAND3X1_62 ( .A(_390_), .B(_392_), .C(_391_), .Y(_393_) );
NOR2X1 NOR2X1_69 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_387_) );
AND2X2 AND2X2_50 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_388_) );
OAI21X1 OAI21X1_55 ( .A(_387_), .B(_388_), .C(w_C_31_), .Y(_389_) );
NAND2X1 NAND2X1_74 ( .A(_389_), .B(_393_), .Y(_197__31_) );
INVX1 INVX1_123 ( .A(w_C_32_), .Y(_397_) );
OR2X2 OR2X2_33 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_398_) );
NAND2X1 NAND2X1_75 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_399_) );
NAND3X1 NAND3X1_63 ( .A(_397_), .B(_399_), .C(_398_), .Y(_400_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_394_) );
AND2X2 AND2X2_51 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_395_) );
OAI21X1 OAI21X1_56 ( .A(_394_), .B(_395_), .C(w_C_32_), .Y(_396_) );
NAND2X1 NAND2X1_76 ( .A(_396_), .B(_400_), .Y(_197__32_) );
INVX1 INVX1_124 ( .A(w_C_33_), .Y(_404_) );
OR2X2 OR2X2_34 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_405_) );
NAND2X1 NAND2X1_77 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_406_) );
NAND3X1 NAND3X1_64 ( .A(_404_), .B(_406_), .C(_405_), .Y(_407_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_401_) );
AND2X2 AND2X2_52 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_402_) );
OAI21X1 OAI21X1_57 ( .A(_401_), .B(_402_), .C(w_C_33_), .Y(_403_) );
NAND2X1 NAND2X1_78 ( .A(_403_), .B(_407_), .Y(_197__33_) );
INVX1 INVX1_125 ( .A(w_C_34_), .Y(_411_) );
OR2X2 OR2X2_35 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_412_) );
NAND2X1 NAND2X1_79 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_413_) );
NAND3X1 NAND3X1_65 ( .A(_411_), .B(_413_), .C(_412_), .Y(_414_) );
NOR2X1 NOR2X1_72 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_408_) );
AND2X2 AND2X2_53 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_409_) );
OAI21X1 OAI21X1_58 ( .A(_408_), .B(_409_), .C(w_C_34_), .Y(_410_) );
NAND2X1 NAND2X1_80 ( .A(_410_), .B(_414_), .Y(_197__34_) );
INVX1 INVX1_126 ( .A(w_C_35_), .Y(_418_) );
OR2X2 OR2X2_36 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_419_) );
NAND2X1 NAND2X1_81 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_420_) );
NAND3X1 NAND3X1_66 ( .A(_418_), .B(_420_), .C(_419_), .Y(_421_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_415_) );
AND2X2 AND2X2_54 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_416_) );
OAI21X1 OAI21X1_59 ( .A(_415_), .B(_416_), .C(w_C_35_), .Y(_417_) );
NAND2X1 NAND2X1_82 ( .A(_417_), .B(_421_), .Y(_197__35_) );
INVX1 INVX1_127 ( .A(1'b0), .Y(_425_) );
OR2X2 OR2X2_37 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_426_) );
NAND2X1 NAND2X1_83 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_427_) );
NAND3X1 NAND3X1_67 ( .A(_425_), .B(_427_), .C(_426_), .Y(_428_) );
NOR2X1 NOR2X1_74 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_422_) );
AND2X2 AND2X2_55 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_423_) );
OAI21X1 OAI21X1_60 ( .A(_422_), .B(_423_), .C(1'b0), .Y(_424_) );
NAND2X1 NAND2X1_84 ( .A(_424_), .B(_428_), .Y(_197__0_) );
INVX1 INVX1_128 ( .A(w_C_1_), .Y(_432_) );
OR2X2 OR2X2_38 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_433_) );
NAND2X1 NAND2X1_85 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_434_) );
NAND3X1 NAND3X1_68 ( .A(_432_), .B(_434_), .C(_433_), .Y(_435_) );
NOR2X1 NOR2X1_75 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_429_) );
AND2X2 AND2X2_56 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_430_) );
OAI21X1 OAI21X1_61 ( .A(_429_), .B(_430_), .C(w_C_1_), .Y(_431_) );
NAND2X1 NAND2X1_86 ( .A(_431_), .B(_435_), .Y(_197__1_) );
INVX1 INVX1_129 ( .A(w_C_2_), .Y(_439_) );
OR2X2 OR2X2_39 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_440_) );
NAND2X1 NAND2X1_87 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_441_) );
NAND3X1 NAND3X1_69 ( .A(_439_), .B(_441_), .C(_440_), .Y(_442_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_436_) );
AND2X2 AND2X2_57 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_437_) );
OAI21X1 OAI21X1_62 ( .A(_436_), .B(_437_), .C(w_C_2_), .Y(_438_) );
NAND2X1 NAND2X1_88 ( .A(_438_), .B(_442_), .Y(_197__2_) );
BUFX2 BUFX2_38 ( .A(w_C_36_), .Y(_197__36_) );
BUFX2 BUFX2_39 ( .A(1'b0), .Y(w_C_0_) );
endmodule
