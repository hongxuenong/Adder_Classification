module CSkipA_59bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [58:0] i_add_term1;
input [58:0] i_add_term2;
output [58:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

NOR2X1 NOR2X1_1 ( .A(i_add_term2[16]), .B(_247_), .Y(_248_) );
INVX1 INVX1_1 ( .A(i_add_term2[16]), .Y(_249_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term1[16]), .B(_249_), .Y(_250_) );
INVX1 INVX1_2 ( .A(i_add_term1[17]), .Y(_251_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[17]), .B(_251_), .Y(_252_) );
INVX1 INVX1_3 ( .A(i_add_term2[17]), .Y(_253_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term1[17]), .B(_253_), .Y(_254_) );
OAI22X1 OAI22X1_1 ( .A(_248_), .B(_250_), .C(_252_), .D(_254_), .Y(_255_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_256_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_257_) );
NOR2X1 NOR2X1_6 ( .A(_256_), .B(_257_), .Y(_258_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_259_) );
NAND2X1 NAND2X1_1 ( .A(_258_), .B(_259_), .Y(_260_) );
NOR2X1 NOR2X1_7 ( .A(_255_), .B(_260_), .Y(_15_) );
INVX1 INVX1_4 ( .A(_13_), .Y(_261_) );
NAND2X1 NAND2X1_2 ( .A(gnd), .B(_15_), .Y(_262_) );
OAI21X1 OAI21X1_1 ( .A(_15_), .B(_261_), .C(_262_), .Y(w_cout_5_) );
INVX1 INVX1_5 ( .A(w_cout_5_), .Y(_266_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_267_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_268_) );
NAND3X1 NAND3X1_1 ( .A(_266_), .B(_268_), .C(_267_), .Y(_269_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_263_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_264_) );
OAI21X1 OAI21X1_2 ( .A(_263_), .B(_264_), .C(w_cout_5_), .Y(_265_) );
NAND2X1 NAND2X1_4 ( .A(_265_), .B(_269_), .Y(_0__20_) );
OAI21X1 OAI21X1_3 ( .A(_266_), .B(_263_), .C(_268_), .Y(_17__1_) );
INVX1 INVX1_6 ( .A(_17__3_), .Y(_273_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_274_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_275_) );
NAND3X1 NAND3X1_2 ( .A(_273_), .B(_275_), .C(_274_), .Y(_276_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_270_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_271_) );
OAI21X1 OAI21X1_4 ( .A(_270_), .B(_271_), .C(_17__3_), .Y(_272_) );
NAND2X1 NAND2X1_6 ( .A(_272_), .B(_276_), .Y(_0__23_) );
OAI21X1 OAI21X1_5 ( .A(_273_), .B(_270_), .C(_275_), .Y(_16_) );
INVX1 INVX1_7 ( .A(_17__1_), .Y(_280_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_281_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_282_) );
NAND3X1 NAND3X1_3 ( .A(_280_), .B(_282_), .C(_281_), .Y(_283_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_277_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_278_) );
OAI21X1 OAI21X1_6 ( .A(_277_), .B(_278_), .C(_17__1_), .Y(_279_) );
NAND2X1 NAND2X1_8 ( .A(_279_), .B(_283_), .Y(_0__21_) );
OAI21X1 OAI21X1_7 ( .A(_280_), .B(_277_), .C(_282_), .Y(_17__2_) );
INVX1 INVX1_8 ( .A(_17__2_), .Y(_287_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_288_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_289_) );
NAND3X1 NAND3X1_4 ( .A(_287_), .B(_289_), .C(_288_), .Y(_290_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_284_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_285_) );
OAI21X1 OAI21X1_8 ( .A(_284_), .B(_285_), .C(_17__2_), .Y(_286_) );
NAND2X1 NAND2X1_10 ( .A(_286_), .B(_290_), .Y(_0__22_) );
OAI21X1 OAI21X1_9 ( .A(_287_), .B(_284_), .C(_289_), .Y(_17__3_) );
INVX1 INVX1_9 ( .A(i_add_term1[20]), .Y(_291_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[20]), .B(_291_), .Y(_292_) );
INVX1 INVX1_10 ( .A(i_add_term2[20]), .Y(_293_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term1[20]), .B(_293_), .Y(_294_) );
INVX1 INVX1_11 ( .A(i_add_term1[21]), .Y(_295_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[21]), .B(_295_), .Y(_296_) );
INVX1 INVX1_12 ( .A(i_add_term2[21]), .Y(_297_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term1[21]), .B(_297_), .Y(_298_) );
OAI22X1 OAI22X1_2 ( .A(_292_), .B(_294_), .C(_296_), .D(_298_), .Y(_299_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_300_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_301_) );
NOR2X1 NOR2X1_17 ( .A(_300_), .B(_301_), .Y(_302_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_303_) );
NAND2X1 NAND2X1_11 ( .A(_302_), .B(_303_), .Y(_304_) );
NOR2X1 NOR2X1_18 ( .A(_299_), .B(_304_), .Y(_18_) );
INVX1 INVX1_13 ( .A(_16_), .Y(_305_) );
NAND2X1 NAND2X1_12 ( .A(gnd), .B(_18_), .Y(_306_) );
OAI21X1 OAI21X1_10 ( .A(_18_), .B(_305_), .C(_306_), .Y(w_cout_6_) );
INVX1 INVX1_14 ( .A(w_cout_6_), .Y(_310_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_311_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_312_) );
NAND3X1 NAND3X1_5 ( .A(_310_), .B(_312_), .C(_311_), .Y(_313_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_307_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_308_) );
OAI21X1 OAI21X1_11 ( .A(_307_), .B(_308_), .C(w_cout_6_), .Y(_309_) );
NAND2X1 NAND2X1_14 ( .A(_309_), .B(_313_), .Y(_0__24_) );
OAI21X1 OAI21X1_12 ( .A(_310_), .B(_307_), .C(_312_), .Y(_20__1_) );
INVX1 INVX1_15 ( .A(_20__3_), .Y(_317_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_318_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_319_) );
NAND3X1 NAND3X1_6 ( .A(_317_), .B(_319_), .C(_318_), .Y(_320_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_314_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_315_) );
OAI21X1 OAI21X1_13 ( .A(_314_), .B(_315_), .C(_20__3_), .Y(_316_) );
NAND2X1 NAND2X1_16 ( .A(_316_), .B(_320_), .Y(_0__27_) );
OAI21X1 OAI21X1_14 ( .A(_317_), .B(_314_), .C(_319_), .Y(_19_) );
INVX1 INVX1_16 ( .A(_20__1_), .Y(_324_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_325_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_326_) );
NAND3X1 NAND3X1_7 ( .A(_324_), .B(_326_), .C(_325_), .Y(_327_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_321_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_322_) );
OAI21X1 OAI21X1_15 ( .A(_321_), .B(_322_), .C(_20__1_), .Y(_323_) );
NAND2X1 NAND2X1_18 ( .A(_323_), .B(_327_), .Y(_0__25_) );
OAI21X1 OAI21X1_16 ( .A(_324_), .B(_321_), .C(_326_), .Y(_20__2_) );
INVX1 INVX1_17 ( .A(_20__2_), .Y(_331_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_332_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_333_) );
NAND3X1 NAND3X1_8 ( .A(_331_), .B(_333_), .C(_332_), .Y(_334_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_328_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_329_) );
OAI21X1 OAI21X1_17 ( .A(_328_), .B(_329_), .C(_20__2_), .Y(_330_) );
NAND2X1 NAND2X1_20 ( .A(_330_), .B(_334_), .Y(_0__26_) );
OAI21X1 OAI21X1_18 ( .A(_331_), .B(_328_), .C(_333_), .Y(_20__3_) );
INVX1 INVX1_18 ( .A(i_add_term1[24]), .Y(_335_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[24]), .B(_335_), .Y(_336_) );
INVX1 INVX1_19 ( .A(i_add_term2[24]), .Y(_337_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term1[24]), .B(_337_), .Y(_338_) );
INVX1 INVX1_20 ( .A(i_add_term1[25]), .Y(_339_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[25]), .B(_339_), .Y(_340_) );
INVX1 INVX1_21 ( .A(i_add_term2[25]), .Y(_341_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term1[25]), .B(_341_), .Y(_342_) );
OAI22X1 OAI22X1_3 ( .A(_336_), .B(_338_), .C(_340_), .D(_342_), .Y(_343_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_344_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_345_) );
NOR2X1 NOR2X1_28 ( .A(_344_), .B(_345_), .Y(_346_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_347_) );
NAND2X1 NAND2X1_21 ( .A(_346_), .B(_347_), .Y(_348_) );
NOR2X1 NOR2X1_29 ( .A(_343_), .B(_348_), .Y(_21_) );
INVX1 INVX1_22 ( .A(_19_), .Y(_349_) );
NAND2X1 NAND2X1_22 ( .A(gnd), .B(_21_), .Y(_350_) );
OAI21X1 OAI21X1_19 ( .A(_21_), .B(_349_), .C(_350_), .Y(w_cout_7_) );
INVX1 INVX1_23 ( .A(w_cout_7_), .Y(_354_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_355_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_356_) );
NAND3X1 NAND3X1_9 ( .A(_354_), .B(_356_), .C(_355_), .Y(_357_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_351_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_352_) );
OAI21X1 OAI21X1_20 ( .A(_351_), .B(_352_), .C(w_cout_7_), .Y(_353_) );
NAND2X1 NAND2X1_24 ( .A(_353_), .B(_357_), .Y(_0__28_) );
OAI21X1 OAI21X1_21 ( .A(_354_), .B(_351_), .C(_356_), .Y(_23__1_) );
INVX1 INVX1_24 ( .A(_23__3_), .Y(_361_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_362_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_363_) );
NAND3X1 NAND3X1_10 ( .A(_361_), .B(_363_), .C(_362_), .Y(_364_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_358_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_359_) );
OAI21X1 OAI21X1_22 ( .A(_358_), .B(_359_), .C(_23__3_), .Y(_360_) );
NAND2X1 NAND2X1_26 ( .A(_360_), .B(_364_), .Y(_0__31_) );
OAI21X1 OAI21X1_23 ( .A(_361_), .B(_358_), .C(_363_), .Y(_22_) );
INVX1 INVX1_25 ( .A(_23__1_), .Y(_368_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_369_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_370_) );
NAND3X1 NAND3X1_11 ( .A(_368_), .B(_370_), .C(_369_), .Y(_371_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_365_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_366_) );
OAI21X1 OAI21X1_24 ( .A(_365_), .B(_366_), .C(_23__1_), .Y(_367_) );
NAND2X1 NAND2X1_28 ( .A(_367_), .B(_371_), .Y(_0__29_) );
OAI21X1 OAI21X1_25 ( .A(_368_), .B(_365_), .C(_370_), .Y(_23__2_) );
INVX1 INVX1_26 ( .A(_23__2_), .Y(_375_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_376_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_377_) );
NAND3X1 NAND3X1_12 ( .A(_375_), .B(_377_), .C(_376_), .Y(_378_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_372_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_373_) );
OAI21X1 OAI21X1_26 ( .A(_372_), .B(_373_), .C(_23__2_), .Y(_374_) );
NAND2X1 NAND2X1_30 ( .A(_374_), .B(_378_), .Y(_0__30_) );
OAI21X1 OAI21X1_27 ( .A(_375_), .B(_372_), .C(_377_), .Y(_23__3_) );
INVX1 INVX1_27 ( .A(i_add_term1[28]), .Y(_379_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[28]), .B(_379_), .Y(_380_) );
INVX1 INVX1_28 ( .A(i_add_term2[28]), .Y(_381_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term1[28]), .B(_381_), .Y(_382_) );
INVX1 INVX1_29 ( .A(i_add_term1[29]), .Y(_383_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[29]), .B(_383_), .Y(_384_) );
INVX1 INVX1_30 ( .A(i_add_term2[29]), .Y(_385_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term1[29]), .B(_385_), .Y(_386_) );
OAI22X1 OAI22X1_4 ( .A(_380_), .B(_382_), .C(_384_), .D(_386_), .Y(_387_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_388_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_389_) );
NOR2X1 NOR2X1_39 ( .A(_388_), .B(_389_), .Y(_390_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_391_) );
NAND2X1 NAND2X1_31 ( .A(_390_), .B(_391_), .Y(_392_) );
NOR2X1 NOR2X1_40 ( .A(_387_), .B(_392_), .Y(_24_) );
INVX1 INVX1_31 ( .A(_22_), .Y(_393_) );
NAND2X1 NAND2X1_32 ( .A(gnd), .B(_24_), .Y(_394_) );
OAI21X1 OAI21X1_28 ( .A(_24_), .B(_393_), .C(_394_), .Y(w_cout_8_) );
INVX1 INVX1_32 ( .A(w_cout_8_), .Y(_398_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_399_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_400_) );
NAND3X1 NAND3X1_13 ( .A(_398_), .B(_400_), .C(_399_), .Y(_401_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_395_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_396_) );
OAI21X1 OAI21X1_29 ( .A(_395_), .B(_396_), .C(w_cout_8_), .Y(_397_) );
NAND2X1 NAND2X1_34 ( .A(_397_), .B(_401_), .Y(_0__32_) );
OAI21X1 OAI21X1_30 ( .A(_398_), .B(_395_), .C(_400_), .Y(_26__1_) );
INVX1 INVX1_33 ( .A(_26__3_), .Y(_405_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_406_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_407_) );
NAND3X1 NAND3X1_14 ( .A(_405_), .B(_407_), .C(_406_), .Y(_408_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_402_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_403_) );
OAI21X1 OAI21X1_31 ( .A(_402_), .B(_403_), .C(_26__3_), .Y(_404_) );
NAND2X1 NAND2X1_36 ( .A(_404_), .B(_408_), .Y(_0__35_) );
OAI21X1 OAI21X1_32 ( .A(_405_), .B(_402_), .C(_407_), .Y(_25_) );
INVX1 INVX1_34 ( .A(_26__1_), .Y(_412_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_413_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_414_) );
NAND3X1 NAND3X1_15 ( .A(_412_), .B(_414_), .C(_413_), .Y(_415_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_409_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_410_) );
OAI21X1 OAI21X1_33 ( .A(_409_), .B(_410_), .C(_26__1_), .Y(_411_) );
NAND2X1 NAND2X1_38 ( .A(_411_), .B(_415_), .Y(_0__33_) );
OAI21X1 OAI21X1_34 ( .A(_412_), .B(_409_), .C(_414_), .Y(_26__2_) );
INVX1 INVX1_35 ( .A(_26__2_), .Y(_419_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_420_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_421_) );
NAND3X1 NAND3X1_16 ( .A(_419_), .B(_421_), .C(_420_), .Y(_422_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_416_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_417_) );
OAI21X1 OAI21X1_35 ( .A(_416_), .B(_417_), .C(_26__2_), .Y(_418_) );
NAND2X1 NAND2X1_40 ( .A(_418_), .B(_422_), .Y(_0__34_) );
OAI21X1 OAI21X1_36 ( .A(_419_), .B(_416_), .C(_421_), .Y(_26__3_) );
INVX1 INVX1_36 ( .A(i_add_term1[32]), .Y(_423_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[32]), .B(_423_), .Y(_424_) );
INVX1 INVX1_37 ( .A(i_add_term2[32]), .Y(_425_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term1[32]), .B(_425_), .Y(_426_) );
INVX1 INVX1_38 ( .A(i_add_term1[33]), .Y(_427_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[33]), .B(_427_), .Y(_428_) );
INVX1 INVX1_39 ( .A(i_add_term2[33]), .Y(_429_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term1[33]), .B(_429_), .Y(_430_) );
OAI22X1 OAI22X1_5 ( .A(_424_), .B(_426_), .C(_428_), .D(_430_), .Y(_431_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_432_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_433_) );
NOR2X1 NOR2X1_50 ( .A(_432_), .B(_433_), .Y(_434_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_435_) );
NAND2X1 NAND2X1_41 ( .A(_434_), .B(_435_), .Y(_436_) );
NOR2X1 NOR2X1_51 ( .A(_431_), .B(_436_), .Y(_27_) );
INVX1 INVX1_40 ( .A(_25_), .Y(_437_) );
NAND2X1 NAND2X1_42 ( .A(gnd), .B(_27_), .Y(_438_) );
OAI21X1 OAI21X1_37 ( .A(_27_), .B(_437_), .C(_438_), .Y(w_cout_9_) );
INVX1 INVX1_41 ( .A(w_cout_9_), .Y(_442_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_443_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_444_) );
NAND3X1 NAND3X1_17 ( .A(_442_), .B(_444_), .C(_443_), .Y(_445_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_439_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_440_) );
OAI21X1 OAI21X1_38 ( .A(_439_), .B(_440_), .C(w_cout_9_), .Y(_441_) );
NAND2X1 NAND2X1_44 ( .A(_441_), .B(_445_), .Y(_0__36_) );
OAI21X1 OAI21X1_39 ( .A(_442_), .B(_439_), .C(_444_), .Y(_29__1_) );
INVX1 INVX1_42 ( .A(_29__3_), .Y(_449_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_450_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_451_) );
NAND3X1 NAND3X1_18 ( .A(_449_), .B(_451_), .C(_450_), .Y(_452_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_446_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_447_) );
OAI21X1 OAI21X1_40 ( .A(_446_), .B(_447_), .C(_29__3_), .Y(_448_) );
NAND2X1 NAND2X1_46 ( .A(_448_), .B(_452_), .Y(_0__39_) );
OAI21X1 OAI21X1_41 ( .A(_449_), .B(_446_), .C(_451_), .Y(_28_) );
INVX1 INVX1_43 ( .A(_29__1_), .Y(_456_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_457_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_458_) );
NAND3X1 NAND3X1_19 ( .A(_456_), .B(_458_), .C(_457_), .Y(_459_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_453_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_454_) );
OAI21X1 OAI21X1_42 ( .A(_453_), .B(_454_), .C(_29__1_), .Y(_455_) );
NAND2X1 NAND2X1_48 ( .A(_455_), .B(_459_), .Y(_0__37_) );
OAI21X1 OAI21X1_43 ( .A(_456_), .B(_453_), .C(_458_), .Y(_29__2_) );
INVX1 INVX1_44 ( .A(_29__2_), .Y(_463_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_464_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_465_) );
NAND3X1 NAND3X1_20 ( .A(_463_), .B(_465_), .C(_464_), .Y(_466_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_460_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_461_) );
OAI21X1 OAI21X1_44 ( .A(_460_), .B(_461_), .C(_29__2_), .Y(_462_) );
NAND2X1 NAND2X1_50 ( .A(_462_), .B(_466_), .Y(_0__38_) );
OAI21X1 OAI21X1_45 ( .A(_463_), .B(_460_), .C(_465_), .Y(_29__3_) );
INVX1 INVX1_45 ( .A(i_add_term1[36]), .Y(_467_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[36]), .B(_467_), .Y(_468_) );
INVX1 INVX1_46 ( .A(i_add_term2[36]), .Y(_469_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term1[36]), .B(_469_), .Y(_470_) );
INVX1 INVX1_47 ( .A(i_add_term1[37]), .Y(_471_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[37]), .B(_471_), .Y(_472_) );
INVX1 INVX1_48 ( .A(i_add_term2[37]), .Y(_473_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term1[37]), .B(_473_), .Y(_474_) );
OAI22X1 OAI22X1_6 ( .A(_468_), .B(_470_), .C(_472_), .D(_474_), .Y(_475_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_476_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_477_) );
NOR2X1 NOR2X1_61 ( .A(_476_), .B(_477_), .Y(_478_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_479_) );
NAND2X1 NAND2X1_51 ( .A(_478_), .B(_479_), .Y(_480_) );
NOR2X1 NOR2X1_62 ( .A(_475_), .B(_480_), .Y(_30_) );
INVX1 INVX1_49 ( .A(_28_), .Y(_481_) );
NAND2X1 NAND2X1_52 ( .A(gnd), .B(_30_), .Y(_482_) );
OAI21X1 OAI21X1_46 ( .A(_30_), .B(_481_), .C(_482_), .Y(w_cout_10_) );
INVX1 INVX1_50 ( .A(w_cout_10_), .Y(_486_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_487_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_488_) );
NAND3X1 NAND3X1_21 ( .A(_486_), .B(_488_), .C(_487_), .Y(_489_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_483_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_484_) );
OAI21X1 OAI21X1_47 ( .A(_483_), .B(_484_), .C(w_cout_10_), .Y(_485_) );
NAND2X1 NAND2X1_54 ( .A(_485_), .B(_489_), .Y(_0__40_) );
OAI21X1 OAI21X1_48 ( .A(_486_), .B(_483_), .C(_488_), .Y(_32__1_) );
INVX1 INVX1_51 ( .A(_32__3_), .Y(_493_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_494_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_495_) );
NAND3X1 NAND3X1_22 ( .A(_493_), .B(_495_), .C(_494_), .Y(_496_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_490_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_491_) );
OAI21X1 OAI21X1_49 ( .A(_490_), .B(_491_), .C(_32__3_), .Y(_492_) );
NAND2X1 NAND2X1_56 ( .A(_492_), .B(_496_), .Y(_0__43_) );
OAI21X1 OAI21X1_50 ( .A(_493_), .B(_490_), .C(_495_), .Y(_31_) );
INVX1 INVX1_52 ( .A(_32__1_), .Y(_500_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_501_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_502_) );
NAND3X1 NAND3X1_23 ( .A(_500_), .B(_502_), .C(_501_), .Y(_503_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_497_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_498_) );
OAI21X1 OAI21X1_51 ( .A(_497_), .B(_498_), .C(_32__1_), .Y(_499_) );
NAND2X1 NAND2X1_58 ( .A(_499_), .B(_503_), .Y(_0__41_) );
OAI21X1 OAI21X1_52 ( .A(_500_), .B(_497_), .C(_502_), .Y(_32__2_) );
INVX1 INVX1_53 ( .A(_32__2_), .Y(_507_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_508_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_509_) );
NAND3X1 NAND3X1_24 ( .A(_507_), .B(_509_), .C(_508_), .Y(_510_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_504_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_505_) );
OAI21X1 OAI21X1_53 ( .A(_504_), .B(_505_), .C(_32__2_), .Y(_506_) );
NAND2X1 NAND2X1_60 ( .A(_506_), .B(_510_), .Y(_0__42_) );
OAI21X1 OAI21X1_54 ( .A(_507_), .B(_504_), .C(_509_), .Y(_32__3_) );
INVX1 INVX1_54 ( .A(i_add_term1[40]), .Y(_511_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[40]), .B(_511_), .Y(_512_) );
INVX1 INVX1_55 ( .A(i_add_term2[40]), .Y(_513_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term1[40]), .B(_513_), .Y(_514_) );
INVX1 INVX1_56 ( .A(i_add_term1[41]), .Y(_515_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[41]), .B(_515_), .Y(_516_) );
INVX1 INVX1_57 ( .A(i_add_term2[41]), .Y(_517_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term1[41]), .B(_517_), .Y(_518_) );
OAI22X1 OAI22X1_7 ( .A(_512_), .B(_514_), .C(_516_), .D(_518_), .Y(_519_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_520_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_521_) );
NOR2X1 NOR2X1_72 ( .A(_520_), .B(_521_), .Y(_522_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_523_) );
NAND2X1 NAND2X1_61 ( .A(_522_), .B(_523_), .Y(_524_) );
NOR2X1 NOR2X1_73 ( .A(_519_), .B(_524_), .Y(_33_) );
INVX1 INVX1_58 ( .A(_31_), .Y(_525_) );
NAND2X1 NAND2X1_62 ( .A(gnd), .B(_33_), .Y(_526_) );
OAI21X1 OAI21X1_55 ( .A(_33_), .B(_525_), .C(_526_), .Y(w_cout_11_) );
INVX1 INVX1_59 ( .A(w_cout_11_), .Y(_530_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_531_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_532_) );
NAND3X1 NAND3X1_25 ( .A(_530_), .B(_532_), .C(_531_), .Y(_533_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_527_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_528_) );
OAI21X1 OAI21X1_56 ( .A(_527_), .B(_528_), .C(w_cout_11_), .Y(_529_) );
NAND2X1 NAND2X1_64 ( .A(_529_), .B(_533_), .Y(_0__44_) );
OAI21X1 OAI21X1_57 ( .A(_530_), .B(_527_), .C(_532_), .Y(_35__1_) );
INVX1 INVX1_60 ( .A(_35__3_), .Y(_537_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_538_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_539_) );
NAND3X1 NAND3X1_26 ( .A(_537_), .B(_539_), .C(_538_), .Y(_540_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_534_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_535_) );
OAI21X1 OAI21X1_58 ( .A(_534_), .B(_535_), .C(_35__3_), .Y(_536_) );
NAND2X1 NAND2X1_66 ( .A(_536_), .B(_540_), .Y(_0__47_) );
OAI21X1 OAI21X1_59 ( .A(_537_), .B(_534_), .C(_539_), .Y(_34_) );
INVX1 INVX1_61 ( .A(_35__1_), .Y(_544_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_545_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_546_) );
NAND3X1 NAND3X1_27 ( .A(_544_), .B(_546_), .C(_545_), .Y(_547_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_541_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_542_) );
OAI21X1 OAI21X1_60 ( .A(_541_), .B(_542_), .C(_35__1_), .Y(_543_) );
NAND2X1 NAND2X1_68 ( .A(_543_), .B(_547_), .Y(_0__45_) );
OAI21X1 OAI21X1_61 ( .A(_544_), .B(_541_), .C(_546_), .Y(_35__2_) );
INVX1 INVX1_62 ( .A(_35__2_), .Y(_551_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_552_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_553_) );
NAND3X1 NAND3X1_28 ( .A(_551_), .B(_553_), .C(_552_), .Y(_554_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_548_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_549_) );
OAI21X1 OAI21X1_62 ( .A(_548_), .B(_549_), .C(_35__2_), .Y(_550_) );
NAND2X1 NAND2X1_70 ( .A(_550_), .B(_554_), .Y(_0__46_) );
OAI21X1 OAI21X1_63 ( .A(_551_), .B(_548_), .C(_553_), .Y(_35__3_) );
INVX1 INVX1_63 ( .A(i_add_term1[44]), .Y(_555_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[44]), .B(_555_), .Y(_556_) );
INVX1 INVX1_64 ( .A(i_add_term2[44]), .Y(_557_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term1[44]), .B(_557_), .Y(_558_) );
INVX1 INVX1_65 ( .A(i_add_term1[45]), .Y(_559_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[45]), .B(_559_), .Y(_560_) );
INVX1 INVX1_66 ( .A(i_add_term2[45]), .Y(_561_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term1[45]), .B(_561_), .Y(_562_) );
OAI22X1 OAI22X1_8 ( .A(_556_), .B(_558_), .C(_560_), .D(_562_), .Y(_563_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_564_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_565_) );
NOR2X1 NOR2X1_83 ( .A(_564_), .B(_565_), .Y(_566_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_567_) );
NAND2X1 NAND2X1_71 ( .A(_566_), .B(_567_), .Y(_568_) );
NOR2X1 NOR2X1_84 ( .A(_563_), .B(_568_), .Y(_36_) );
INVX1 INVX1_67 ( .A(_34_), .Y(_569_) );
NAND2X1 NAND2X1_72 ( .A(gnd), .B(_36_), .Y(_570_) );
OAI21X1 OAI21X1_64 ( .A(_36_), .B(_569_), .C(_570_), .Y(w_cout_12_) );
INVX1 INVX1_68 ( .A(w_cout_12_), .Y(_574_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_575_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_576_) );
NAND3X1 NAND3X1_29 ( .A(_574_), .B(_576_), .C(_575_), .Y(_577_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_571_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_572_) );
OAI21X1 OAI21X1_65 ( .A(_571_), .B(_572_), .C(w_cout_12_), .Y(_573_) );
NAND2X1 NAND2X1_74 ( .A(_573_), .B(_577_), .Y(_0__48_) );
OAI21X1 OAI21X1_66 ( .A(_574_), .B(_571_), .C(_576_), .Y(_38__1_) );
INVX1 INVX1_69 ( .A(_38__3_), .Y(_581_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_582_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_583_) );
NAND3X1 NAND3X1_30 ( .A(_581_), .B(_583_), .C(_582_), .Y(_584_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_578_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_579_) );
OAI21X1 OAI21X1_67 ( .A(_578_), .B(_579_), .C(_38__3_), .Y(_580_) );
NAND2X1 NAND2X1_76 ( .A(_580_), .B(_584_), .Y(_0__51_) );
OAI21X1 OAI21X1_68 ( .A(_581_), .B(_578_), .C(_583_), .Y(_37_) );
INVX1 INVX1_70 ( .A(_38__1_), .Y(_588_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_589_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_590_) );
NAND3X1 NAND3X1_31 ( .A(_588_), .B(_590_), .C(_589_), .Y(_591_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_585_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_586_) );
OAI21X1 OAI21X1_69 ( .A(_585_), .B(_586_), .C(_38__1_), .Y(_587_) );
NAND2X1 NAND2X1_78 ( .A(_587_), .B(_591_), .Y(_0__49_) );
OAI21X1 OAI21X1_70 ( .A(_588_), .B(_585_), .C(_590_), .Y(_38__2_) );
INVX1 INVX1_71 ( .A(_38__2_), .Y(_595_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_596_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_597_) );
NAND3X1 NAND3X1_32 ( .A(_595_), .B(_597_), .C(_596_), .Y(_598_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_592_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_593_) );
OAI21X1 OAI21X1_71 ( .A(_592_), .B(_593_), .C(_38__2_), .Y(_594_) );
NAND2X1 NAND2X1_80 ( .A(_594_), .B(_598_), .Y(_0__50_) );
OAI21X1 OAI21X1_72 ( .A(_595_), .B(_592_), .C(_597_), .Y(_38__3_) );
INVX1 INVX1_72 ( .A(i_add_term1[48]), .Y(_599_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[48]), .B(_599_), .Y(_600_) );
INVX1 INVX1_73 ( .A(i_add_term2[48]), .Y(_601_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term1[48]), .B(_601_), .Y(_602_) );
INVX1 INVX1_74 ( .A(i_add_term1[49]), .Y(_603_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[49]), .B(_603_), .Y(_604_) );
INVX1 INVX1_75 ( .A(i_add_term2[49]), .Y(_605_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term1[49]), .B(_605_), .Y(_606_) );
OAI22X1 OAI22X1_9 ( .A(_600_), .B(_602_), .C(_604_), .D(_606_), .Y(_607_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_608_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_609_) );
NOR2X1 NOR2X1_94 ( .A(_608_), .B(_609_), .Y(_610_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_611_) );
NAND2X1 NAND2X1_81 ( .A(_610_), .B(_611_), .Y(_612_) );
NOR2X1 NOR2X1_95 ( .A(_607_), .B(_612_), .Y(_39_) );
INVX1 INVX1_76 ( .A(_37_), .Y(_613_) );
NAND2X1 NAND2X1_82 ( .A(gnd), .B(_39_), .Y(_614_) );
OAI21X1 OAI21X1_73 ( .A(_39_), .B(_613_), .C(_614_), .Y(w_cout_13_) );
INVX1 INVX1_77 ( .A(w_cout_13_), .Y(_618_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_619_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_620_) );
NAND3X1 NAND3X1_33 ( .A(_618_), .B(_620_), .C(_619_), .Y(_621_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_615_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_616_) );
OAI21X1 OAI21X1_74 ( .A(_615_), .B(_616_), .C(w_cout_13_), .Y(_617_) );
NAND2X1 NAND2X1_84 ( .A(_617_), .B(_621_), .Y(_0__52_) );
OAI21X1 OAI21X1_75 ( .A(_618_), .B(_615_), .C(_620_), .Y(_41__1_) );
INVX1 INVX1_78 ( .A(_41__3_), .Y(_625_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_626_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_627_) );
NAND3X1 NAND3X1_34 ( .A(_625_), .B(_627_), .C(_626_), .Y(_628_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_622_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_623_) );
OAI21X1 OAI21X1_76 ( .A(_622_), .B(_623_), .C(_41__3_), .Y(_624_) );
NAND2X1 NAND2X1_86 ( .A(_624_), .B(_628_), .Y(_0__55_) );
OAI21X1 OAI21X1_77 ( .A(_625_), .B(_622_), .C(_627_), .Y(_40_) );
INVX1 INVX1_79 ( .A(_41__1_), .Y(_632_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_633_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_634_) );
NAND3X1 NAND3X1_35 ( .A(_632_), .B(_634_), .C(_633_), .Y(_635_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_629_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_630_) );
OAI21X1 OAI21X1_78 ( .A(_629_), .B(_630_), .C(_41__1_), .Y(_631_) );
NAND2X1 NAND2X1_88 ( .A(_631_), .B(_635_), .Y(_0__53_) );
OAI21X1 OAI21X1_79 ( .A(_632_), .B(_629_), .C(_634_), .Y(_41__2_) );
INVX1 INVX1_80 ( .A(_41__2_), .Y(_639_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_640_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_641_) );
NAND3X1 NAND3X1_36 ( .A(_639_), .B(_641_), .C(_640_), .Y(_642_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_636_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_637_) );
OAI21X1 OAI21X1_80 ( .A(_636_), .B(_637_), .C(_41__2_), .Y(_638_) );
NAND2X1 NAND2X1_90 ( .A(_638_), .B(_642_), .Y(_0__54_) );
OAI21X1 OAI21X1_81 ( .A(_639_), .B(_636_), .C(_641_), .Y(_41__3_) );
INVX1 INVX1_81 ( .A(i_add_term1[52]), .Y(_643_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[52]), .B(_643_), .Y(_644_) );
INVX1 INVX1_82 ( .A(i_add_term2[52]), .Y(_645_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term1[52]), .B(_645_), .Y(_646_) );
INVX1 INVX1_83 ( .A(i_add_term1[53]), .Y(_647_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[53]), .B(_647_), .Y(_648_) );
INVX1 INVX1_84 ( .A(i_add_term2[53]), .Y(_649_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term1[53]), .B(_649_), .Y(_650_) );
OAI22X1 OAI22X1_10 ( .A(_644_), .B(_646_), .C(_648_), .D(_650_), .Y(_651_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_652_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_653_) );
NOR2X1 NOR2X1_105 ( .A(_652_), .B(_653_), .Y(_654_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_655_) );
NAND2X1 NAND2X1_91 ( .A(_654_), .B(_655_), .Y(_656_) );
NOR2X1 NOR2X1_106 ( .A(_651_), .B(_656_), .Y(_42_) );
INVX1 INVX1_85 ( .A(_40_), .Y(_657_) );
NAND2X1 NAND2X1_92 ( .A(gnd), .B(_42_), .Y(_658_) );
OAI21X1 OAI21X1_82 ( .A(_42_), .B(_657_), .C(_658_), .Y(cskip3_inst_cin) );
INVX1 INVX1_86 ( .A(cskip3_inst_cin), .Y(_662_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_663_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_664_) );
NAND3X1 NAND3X1_37 ( .A(_662_), .B(_664_), .C(_663_), .Y(_665_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_659_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_660_) );
OAI21X1 OAI21X1_83 ( .A(_659_), .B(_660_), .C(cskip3_inst_cin), .Y(_661_) );
NAND2X1 NAND2X1_94 ( .A(_661_), .B(_665_), .Y(cskip3_inst_rca0_fa0_o_sum) );
OAI21X1 OAI21X1_84 ( .A(_662_), .B(_659_), .C(_664_), .Y(cskip3_inst_rca0_fa0_o_carry) );
INVX1 INVX1_87 ( .A(cskip3_inst_rca0_fa0_o_carry), .Y(_669_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_670_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_671_) );
NAND3X1 NAND3X1_38 ( .A(_669_), .B(_671_), .C(_670_), .Y(_672_) );
NOR2X1 NOR2X1_108 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_666_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_667_) );
OAI21X1 OAI21X1_85 ( .A(_666_), .B(_667_), .C(cskip3_inst_rca0_fa0_o_carry), .Y(_668_) );
NAND2X1 NAND2X1_96 ( .A(_668_), .B(_672_), .Y(cskip3_inst_rca0_fa1_o_sum) );
OAI21X1 OAI21X1_86 ( .A(_669_), .B(_666_), .C(_671_), .Y(cskip3_inst_rca0_fa1_o_carry) );
INVX1 INVX1_88 ( .A(cskip3_inst_rca0_fa1_o_carry), .Y(_676_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_677_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_678_) );
NAND3X1 NAND3X1_39 ( .A(_676_), .B(_678_), .C(_677_), .Y(_679_) );
NOR2X1 NOR2X1_109 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_673_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_674_) );
OAI21X1 OAI21X1_87 ( .A(_673_), .B(_674_), .C(cskip3_inst_rca0_fa1_o_carry), .Y(_675_) );
NAND2X1 NAND2X1_98 ( .A(_675_), .B(_679_), .Y(cskip3_inst_rca0_fa2_o_sum) );
OAI21X1 OAI21X1_88 ( .A(_676_), .B(_673_), .C(_678_), .Y(cskip3_inst_cout0) );
OR2X2 OR2X2_40 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_683_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_684_) );
NAND2X1 NAND2X1_100 ( .A(_684_), .B(_683_), .Y(_680_) );
XNOR2X1 XNOR2X1_1 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_681_) );
XNOR2X1 XNOR2X1_2 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_682_) );
NOR3X1 NOR3X1_1 ( .A(_680_), .B(_681_), .C(_682_), .Y(cskip3_inst_skip0_P) );
INVX1 INVX1_89 ( .A(cskip3_inst_cout0), .Y(_685_) );
NAND2X1 NAND2X1_101 ( .A(gnd), .B(cskip3_inst_skip0_P), .Y(_686_) );
OAI21X1 OAI21X1_89 ( .A(cskip3_inst_skip0_P), .B(_685_), .C(_686_), .Y(w_cout_15_) );
BUFX2 BUFX2_1 ( .A(w_cout_15_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .A(_0__54_), .Y(sum[54]) );
BUFX2 BUFX2_57 ( .A(_0__55_), .Y(sum[55]) );
BUFX2 BUFX2_58 ( .A(cskip3_inst_rca0_fa0_o_sum), .Y(sum[56]) );
BUFX2 BUFX2_59 ( .A(cskip3_inst_rca0_fa1_o_sum), .Y(sum[57]) );
BUFX2 BUFX2_60 ( .A(cskip3_inst_rca0_fa2_o_sum), .Y(sum[58]) );
INVX1 INVX1_90 ( .A(gnd), .Y(_46_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_47_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_48_) );
NAND3X1 NAND3X1_40 ( .A(_46_), .B(_48_), .C(_47_), .Y(_49_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_43_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_44_) );
OAI21X1 OAI21X1_90 ( .A(_43_), .B(_44_), .C(gnd), .Y(_45_) );
NAND2X1 NAND2X1_103 ( .A(_45_), .B(_49_), .Y(_0__0_) );
OAI21X1 OAI21X1_91 ( .A(_46_), .B(_43_), .C(_48_), .Y(_2__1_) );
INVX1 INVX1_91 ( .A(_2__3_), .Y(_53_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_54_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_55_) );
NAND3X1 NAND3X1_41 ( .A(_53_), .B(_55_), .C(_54_), .Y(_56_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_50_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_51_) );
OAI21X1 OAI21X1_92 ( .A(_50_), .B(_51_), .C(_2__3_), .Y(_52_) );
NAND2X1 NAND2X1_105 ( .A(_52_), .B(_56_), .Y(_0__3_) );
OAI21X1 OAI21X1_93 ( .A(_53_), .B(_50_), .C(_55_), .Y(_1_) );
INVX1 INVX1_92 ( .A(_2__1_), .Y(_60_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_61_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_62_) );
NAND3X1 NAND3X1_42 ( .A(_60_), .B(_62_), .C(_61_), .Y(_63_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_57_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_58_) );
OAI21X1 OAI21X1_94 ( .A(_57_), .B(_58_), .C(_2__1_), .Y(_59_) );
NAND2X1 NAND2X1_107 ( .A(_59_), .B(_63_), .Y(_0__1_) );
OAI21X1 OAI21X1_95 ( .A(_60_), .B(_57_), .C(_62_), .Y(_2__2_) );
INVX1 INVX1_93 ( .A(_2__2_), .Y(_67_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_68_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_69_) );
NAND3X1 NAND3X1_43 ( .A(_67_), .B(_69_), .C(_68_), .Y(_70_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_64_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_65_) );
OAI21X1 OAI21X1_96 ( .A(_64_), .B(_65_), .C(_2__2_), .Y(_66_) );
NAND2X1 NAND2X1_109 ( .A(_66_), .B(_70_), .Y(_0__2_) );
OAI21X1 OAI21X1_97 ( .A(_67_), .B(_64_), .C(_69_), .Y(_2__3_) );
INVX1 INVX1_94 ( .A(i_add_term1[0]), .Y(_71_) );
NOR2X1 NOR2X1_114 ( .A(i_add_term2[0]), .B(_71_), .Y(_72_) );
INVX1 INVX1_95 ( .A(i_add_term2[0]), .Y(_73_) );
NOR2X1 NOR2X1_115 ( .A(i_add_term1[0]), .B(_73_), .Y(_74_) );
INVX1 INVX1_96 ( .A(i_add_term1[1]), .Y(_75_) );
NOR2X1 NOR2X1_116 ( .A(i_add_term2[1]), .B(_75_), .Y(_76_) );
INVX1 INVX1_97 ( .A(i_add_term2[1]), .Y(_77_) );
NOR2X1 NOR2X1_117 ( .A(i_add_term1[1]), .B(_77_), .Y(_78_) );
OAI22X1 OAI22X1_11 ( .A(_72_), .B(_74_), .C(_76_), .D(_78_), .Y(_79_) );
NOR2X1 NOR2X1_118 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_80_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_81_) );
NOR2X1 NOR2X1_119 ( .A(_80_), .B(_81_), .Y(_82_) );
XOR2X1 XOR2X1_11 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_83_) );
NAND2X1 NAND2X1_110 ( .A(_82_), .B(_83_), .Y(_84_) );
NOR2X1 NOR2X1_120 ( .A(_79_), .B(_84_), .Y(_3_) );
INVX1 INVX1_98 ( .A(_1_), .Y(_85_) );
NAND2X1 NAND2X1_111 ( .A(gnd), .B(_3_), .Y(_86_) );
OAI21X1 OAI21X1_98 ( .A(_3_), .B(_85_), .C(_86_), .Y(w_cout_1_) );
INVX1 INVX1_99 ( .A(w_cout_1_), .Y(_90_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_91_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_92_) );
NAND3X1 NAND3X1_44 ( .A(_90_), .B(_92_), .C(_91_), .Y(_93_) );
NOR2X1 NOR2X1_121 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_87_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_88_) );
OAI21X1 OAI21X1_99 ( .A(_87_), .B(_88_), .C(w_cout_1_), .Y(_89_) );
NAND2X1 NAND2X1_113 ( .A(_89_), .B(_93_), .Y(_0__4_) );
OAI21X1 OAI21X1_100 ( .A(_90_), .B(_87_), .C(_92_), .Y(_5__1_) );
INVX1 INVX1_100 ( .A(_5__3_), .Y(_97_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_98_) );
NAND2X1 NAND2X1_114 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_99_) );
NAND3X1 NAND3X1_45 ( .A(_97_), .B(_99_), .C(_98_), .Y(_100_) );
NOR2X1 NOR2X1_122 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_94_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_95_) );
OAI21X1 OAI21X1_101 ( .A(_94_), .B(_95_), .C(_5__3_), .Y(_96_) );
NAND2X1 NAND2X1_115 ( .A(_96_), .B(_100_), .Y(_0__7_) );
OAI21X1 OAI21X1_102 ( .A(_97_), .B(_94_), .C(_99_), .Y(_4_) );
INVX1 INVX1_101 ( .A(_5__1_), .Y(_104_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_105_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_106_) );
NAND3X1 NAND3X1_46 ( .A(_104_), .B(_106_), .C(_105_), .Y(_107_) );
NOR2X1 NOR2X1_123 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_101_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_102_) );
OAI21X1 OAI21X1_103 ( .A(_101_), .B(_102_), .C(_5__1_), .Y(_103_) );
NAND2X1 NAND2X1_117 ( .A(_103_), .B(_107_), .Y(_0__5_) );
OAI21X1 OAI21X1_104 ( .A(_104_), .B(_101_), .C(_106_), .Y(_5__2_) );
INVX1 INVX1_102 ( .A(_5__2_), .Y(_111_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_112_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_113_) );
NAND3X1 NAND3X1_47 ( .A(_111_), .B(_113_), .C(_112_), .Y(_114_) );
NOR2X1 NOR2X1_124 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_108_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_109_) );
OAI21X1 OAI21X1_105 ( .A(_108_), .B(_109_), .C(_5__2_), .Y(_110_) );
NAND2X1 NAND2X1_119 ( .A(_110_), .B(_114_), .Y(_0__6_) );
OAI21X1 OAI21X1_106 ( .A(_111_), .B(_108_), .C(_113_), .Y(_5__3_) );
INVX1 INVX1_103 ( .A(i_add_term1[4]), .Y(_115_) );
NOR2X1 NOR2X1_125 ( .A(i_add_term2[4]), .B(_115_), .Y(_116_) );
INVX1 INVX1_104 ( .A(i_add_term2[4]), .Y(_117_) );
NOR2X1 NOR2X1_126 ( .A(i_add_term1[4]), .B(_117_), .Y(_118_) );
INVX1 INVX1_105 ( .A(i_add_term1[5]), .Y(_119_) );
NOR2X1 NOR2X1_127 ( .A(i_add_term2[5]), .B(_119_), .Y(_120_) );
INVX1 INVX1_106 ( .A(i_add_term2[5]), .Y(_121_) );
NOR2X1 NOR2X1_128 ( .A(i_add_term1[5]), .B(_121_), .Y(_122_) );
OAI22X1 OAI22X1_12 ( .A(_116_), .B(_118_), .C(_120_), .D(_122_), .Y(_123_) );
NOR2X1 NOR2X1_129 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_124_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_125_) );
NOR2X1 NOR2X1_130 ( .A(_124_), .B(_125_), .Y(_126_) );
XOR2X1 XOR2X1_12 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_127_) );
NAND2X1 NAND2X1_120 ( .A(_126_), .B(_127_), .Y(_128_) );
NOR2X1 NOR2X1_131 ( .A(_123_), .B(_128_), .Y(_6_) );
INVX1 INVX1_107 ( .A(_4_), .Y(_129_) );
NAND2X1 NAND2X1_121 ( .A(gnd), .B(_6_), .Y(_130_) );
OAI21X1 OAI21X1_107 ( .A(_6_), .B(_129_), .C(_130_), .Y(w_cout_2_) );
INVX1 INVX1_108 ( .A(w_cout_2_), .Y(_134_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_135_) );
NAND2X1 NAND2X1_122 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_136_) );
NAND3X1 NAND3X1_48 ( .A(_134_), .B(_136_), .C(_135_), .Y(_137_) );
NOR2X1 NOR2X1_132 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_131_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_132_) );
OAI21X1 OAI21X1_108 ( .A(_131_), .B(_132_), .C(w_cout_2_), .Y(_133_) );
NAND2X1 NAND2X1_123 ( .A(_133_), .B(_137_), .Y(_0__8_) );
OAI21X1 OAI21X1_109 ( .A(_134_), .B(_131_), .C(_136_), .Y(_8__1_) );
INVX1 INVX1_109 ( .A(_8__3_), .Y(_141_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_142_) );
NAND2X1 NAND2X1_124 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_143_) );
NAND3X1 NAND3X1_49 ( .A(_141_), .B(_143_), .C(_142_), .Y(_144_) );
NOR2X1 NOR2X1_133 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_138_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_139_) );
OAI21X1 OAI21X1_110 ( .A(_138_), .B(_139_), .C(_8__3_), .Y(_140_) );
NAND2X1 NAND2X1_125 ( .A(_140_), .B(_144_), .Y(_0__11_) );
OAI21X1 OAI21X1_111 ( .A(_141_), .B(_138_), .C(_143_), .Y(_7_) );
INVX1 INVX1_110 ( .A(_8__1_), .Y(_148_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_149_) );
NAND2X1 NAND2X1_126 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_150_) );
NAND3X1 NAND3X1_50 ( .A(_148_), .B(_150_), .C(_149_), .Y(_151_) );
NOR2X1 NOR2X1_134 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_145_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_146_) );
OAI21X1 OAI21X1_112 ( .A(_145_), .B(_146_), .C(_8__1_), .Y(_147_) );
NAND2X1 NAND2X1_127 ( .A(_147_), .B(_151_), .Y(_0__9_) );
OAI21X1 OAI21X1_113 ( .A(_148_), .B(_145_), .C(_150_), .Y(_8__2_) );
INVX1 INVX1_111 ( .A(_8__2_), .Y(_155_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_156_) );
NAND2X1 NAND2X1_128 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_157_) );
NAND3X1 NAND3X1_51 ( .A(_155_), .B(_157_), .C(_156_), .Y(_158_) );
NOR2X1 NOR2X1_135 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_152_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_153_) );
OAI21X1 OAI21X1_114 ( .A(_152_), .B(_153_), .C(_8__2_), .Y(_154_) );
NAND2X1 NAND2X1_129 ( .A(_154_), .B(_158_), .Y(_0__10_) );
OAI21X1 OAI21X1_115 ( .A(_155_), .B(_152_), .C(_157_), .Y(_8__3_) );
INVX1 INVX1_112 ( .A(i_add_term1[8]), .Y(_159_) );
NOR2X1 NOR2X1_136 ( .A(i_add_term2[8]), .B(_159_), .Y(_160_) );
INVX1 INVX1_113 ( .A(i_add_term2[8]), .Y(_161_) );
NOR2X1 NOR2X1_137 ( .A(i_add_term1[8]), .B(_161_), .Y(_162_) );
INVX1 INVX1_114 ( .A(i_add_term1[9]), .Y(_163_) );
NOR2X1 NOR2X1_138 ( .A(i_add_term2[9]), .B(_163_), .Y(_164_) );
INVX1 INVX1_115 ( .A(i_add_term2[9]), .Y(_165_) );
NOR2X1 NOR2X1_139 ( .A(i_add_term1[9]), .B(_165_), .Y(_166_) );
OAI22X1 OAI22X1_13 ( .A(_160_), .B(_162_), .C(_164_), .D(_166_), .Y(_167_) );
NOR2X1 NOR2X1_140 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_168_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_169_) );
NOR2X1 NOR2X1_141 ( .A(_168_), .B(_169_), .Y(_170_) );
XOR2X1 XOR2X1_13 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_171_) );
NAND2X1 NAND2X1_130 ( .A(_170_), .B(_171_), .Y(_172_) );
NOR2X1 NOR2X1_142 ( .A(_167_), .B(_172_), .Y(_9_) );
INVX1 INVX1_116 ( .A(_7_), .Y(_173_) );
NAND2X1 NAND2X1_131 ( .A(gnd), .B(_9_), .Y(_174_) );
OAI21X1 OAI21X1_116 ( .A(_9_), .B(_173_), .C(_174_), .Y(w_cout_3_) );
INVX1 INVX1_117 ( .A(w_cout_3_), .Y(_178_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_179_) );
NAND2X1 NAND2X1_132 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_180_) );
NAND3X1 NAND3X1_52 ( .A(_178_), .B(_180_), .C(_179_), .Y(_181_) );
NOR2X1 NOR2X1_143 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_175_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_176_) );
OAI21X1 OAI21X1_117 ( .A(_175_), .B(_176_), .C(w_cout_3_), .Y(_177_) );
NAND2X1 NAND2X1_133 ( .A(_177_), .B(_181_), .Y(_0__12_) );
OAI21X1 OAI21X1_118 ( .A(_178_), .B(_175_), .C(_180_), .Y(_11__1_) );
INVX1 INVX1_118 ( .A(_11__3_), .Y(_185_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_186_) );
NAND2X1 NAND2X1_134 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_187_) );
NAND3X1 NAND3X1_53 ( .A(_185_), .B(_187_), .C(_186_), .Y(_188_) );
NOR2X1 NOR2X1_144 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_182_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_183_) );
OAI21X1 OAI21X1_119 ( .A(_182_), .B(_183_), .C(_11__3_), .Y(_184_) );
NAND2X1 NAND2X1_135 ( .A(_184_), .B(_188_), .Y(_0__15_) );
OAI21X1 OAI21X1_120 ( .A(_185_), .B(_182_), .C(_187_), .Y(_10_) );
INVX1 INVX1_119 ( .A(_11__1_), .Y(_192_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_193_) );
NAND2X1 NAND2X1_136 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_194_) );
NAND3X1 NAND3X1_54 ( .A(_192_), .B(_194_), .C(_193_), .Y(_195_) );
NOR2X1 NOR2X1_145 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_189_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_190_) );
OAI21X1 OAI21X1_121 ( .A(_189_), .B(_190_), .C(_11__1_), .Y(_191_) );
NAND2X1 NAND2X1_137 ( .A(_191_), .B(_195_), .Y(_0__13_) );
OAI21X1 OAI21X1_122 ( .A(_192_), .B(_189_), .C(_194_), .Y(_11__2_) );
INVX1 INVX1_120 ( .A(_11__2_), .Y(_199_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_200_) );
NAND2X1 NAND2X1_138 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_201_) );
NAND3X1 NAND3X1_55 ( .A(_199_), .B(_201_), .C(_200_), .Y(_202_) );
NOR2X1 NOR2X1_146 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_196_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_197_) );
OAI21X1 OAI21X1_123 ( .A(_196_), .B(_197_), .C(_11__2_), .Y(_198_) );
NAND2X1 NAND2X1_139 ( .A(_198_), .B(_202_), .Y(_0__14_) );
OAI21X1 OAI21X1_124 ( .A(_199_), .B(_196_), .C(_201_), .Y(_11__3_) );
INVX1 INVX1_121 ( .A(i_add_term1[12]), .Y(_203_) );
NOR2X1 NOR2X1_147 ( .A(i_add_term2[12]), .B(_203_), .Y(_204_) );
INVX1 INVX1_122 ( .A(i_add_term2[12]), .Y(_205_) );
NOR2X1 NOR2X1_148 ( .A(i_add_term1[12]), .B(_205_), .Y(_206_) );
INVX1 INVX1_123 ( .A(i_add_term1[13]), .Y(_207_) );
NOR2X1 NOR2X1_149 ( .A(i_add_term2[13]), .B(_207_), .Y(_208_) );
INVX1 INVX1_124 ( .A(i_add_term2[13]), .Y(_209_) );
NOR2X1 NOR2X1_150 ( .A(i_add_term1[13]), .B(_209_), .Y(_210_) );
OAI22X1 OAI22X1_14 ( .A(_204_), .B(_206_), .C(_208_), .D(_210_), .Y(_211_) );
NOR2X1 NOR2X1_151 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_212_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_213_) );
NOR2X1 NOR2X1_152 ( .A(_212_), .B(_213_), .Y(_214_) );
XOR2X1 XOR2X1_14 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_215_) );
NAND2X1 NAND2X1_140 ( .A(_214_), .B(_215_), .Y(_216_) );
NOR2X1 NOR2X1_153 ( .A(_211_), .B(_216_), .Y(_12_) );
INVX1 INVX1_125 ( .A(_10_), .Y(_217_) );
NAND2X1 NAND2X1_141 ( .A(gnd), .B(_12_), .Y(_218_) );
OAI21X1 OAI21X1_125 ( .A(_12_), .B(_217_), .C(_218_), .Y(w_cout_4_) );
INVX1 INVX1_126 ( .A(w_cout_4_), .Y(_222_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_223_) );
NAND2X1 NAND2X1_142 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_224_) );
NAND3X1 NAND3X1_56 ( .A(_222_), .B(_224_), .C(_223_), .Y(_225_) );
NOR2X1 NOR2X1_154 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_219_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_220_) );
OAI21X1 OAI21X1_126 ( .A(_219_), .B(_220_), .C(w_cout_4_), .Y(_221_) );
NAND2X1 NAND2X1_143 ( .A(_221_), .B(_225_), .Y(_0__16_) );
OAI21X1 OAI21X1_127 ( .A(_222_), .B(_219_), .C(_224_), .Y(_14__1_) );
INVX1 INVX1_127 ( .A(_14__3_), .Y(_229_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_230_) );
NAND2X1 NAND2X1_144 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_231_) );
NAND3X1 NAND3X1_57 ( .A(_229_), .B(_231_), .C(_230_), .Y(_232_) );
NOR2X1 NOR2X1_155 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_226_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_227_) );
OAI21X1 OAI21X1_128 ( .A(_226_), .B(_227_), .C(_14__3_), .Y(_228_) );
NAND2X1 NAND2X1_145 ( .A(_228_), .B(_232_), .Y(_0__19_) );
OAI21X1 OAI21X1_129 ( .A(_229_), .B(_226_), .C(_231_), .Y(_13_) );
INVX1 INVX1_128 ( .A(_14__1_), .Y(_236_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_237_) );
NAND2X1 NAND2X1_146 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_238_) );
NAND3X1 NAND3X1_58 ( .A(_236_), .B(_238_), .C(_237_), .Y(_239_) );
NOR2X1 NOR2X1_156 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_233_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_234_) );
OAI21X1 OAI21X1_130 ( .A(_233_), .B(_234_), .C(_14__1_), .Y(_235_) );
NAND2X1 NAND2X1_147 ( .A(_235_), .B(_239_), .Y(_0__17_) );
OAI21X1 OAI21X1_131 ( .A(_236_), .B(_233_), .C(_238_), .Y(_14__2_) );
INVX1 INVX1_129 ( .A(_14__2_), .Y(_243_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_244_) );
NAND2X1 NAND2X1_148 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_245_) );
NAND3X1 NAND3X1_59 ( .A(_243_), .B(_245_), .C(_244_), .Y(_246_) );
NOR2X1 NOR2X1_157 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_240_) );
AND2X2 AND2X2_73 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_241_) );
OAI21X1 OAI21X1_132 ( .A(_240_), .B(_241_), .C(_14__2_), .Y(_242_) );
NAND2X1 NAND2X1_149 ( .A(_242_), .B(_246_), .Y(_0__18_) );
OAI21X1 OAI21X1_133 ( .A(_243_), .B(_240_), .C(_245_), .Y(_14__3_) );
INVX1 INVX1_130 ( .A(i_add_term1[16]), .Y(_247_) );
BUFX2 BUFX2_61 ( .A(cskip3_inst_rca0_fa0_o_sum), .Y(_0__56_) );
BUFX2 BUFX2_62 ( .A(cskip3_inst_rca0_fa1_o_sum), .Y(_0__57_) );
BUFX2 BUFX2_63 ( .A(cskip3_inst_rca0_fa2_o_sum), .Y(_0__58_) );
BUFX2 BUFX2_64 ( .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_65 ( .A(cskip3_inst_cin), .Y(w_cout_14_) );
endmodule
