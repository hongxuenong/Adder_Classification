module cla_43bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [42:0] i_add1;
input [42:0] i_add2;
output [43:0] o_result;

NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_349_), .C(_348_), .Y(_350_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_344_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_345_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_345_), .C(w_C_17_), .Y(_346_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_350_), .Y(_252__17_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(w_C_18_), .Y(_354_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_355_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_356_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_356_), .C(_355_), .Y(_357_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_351_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_352_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_352_), .C(w_C_18_), .Y(_353_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_357_), .Y(_252__18_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(w_C_19_), .Y(_361_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_362_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_363_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_363_), .C(_362_), .Y(_364_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_358_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_359_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_358_), .B(_359_), .C(w_C_19_), .Y(_360_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_364_), .Y(_252__19_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(w_C_20_), .Y(_368_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_369_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_370_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_370_), .C(_369_), .Y(_371_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_365_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_366_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_365_), .B(_366_), .C(w_C_20_), .Y(_367_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_371_), .Y(_252__20_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(w_C_21_), .Y(_375_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_376_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_377_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_377_), .C(_376_), .Y(_378_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_372_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_373_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_373_), .C(w_C_21_), .Y(_374_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_378_), .Y(_252__21_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(w_C_22_), .Y(_382_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_383_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_384_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_382_), .B(_384_), .C(_383_), .Y(_385_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_379_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_380_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_380_), .C(w_C_22_), .Y(_381_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_385_), .Y(_252__22_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(w_C_23_), .Y(_389_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_390_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_391_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_391_), .C(_390_), .Y(_392_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_386_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_387_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_387_), .C(w_C_23_), .Y(_388_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(_392_), .Y(_252__23_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(w_C_24_), .Y(_396_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_397_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_398_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_398_), .C(_397_), .Y(_399_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_393_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_394_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_394_), .C(w_C_24_), .Y(_395_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_399_), .Y(_252__24_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(w_C_25_), .Y(_403_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_404_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_405_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_405_), .C(_404_), .Y(_406_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_400_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_401_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_400_), .B(_401_), .C(w_C_25_), .Y(_402_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_406_), .Y(_252__25_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(w_C_26_), .Y(_410_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_411_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_412_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(_412_), .C(_411_), .Y(_413_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_407_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_408_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_408_), .C(w_C_26_), .Y(_409_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_413_), .Y(_252__26_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(w_C_27_), .Y(_417_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_418_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_419_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_419_), .C(_418_), .Y(_420_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_414_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_415_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_414_), .B(_415_), .C(w_C_27_), .Y(_416_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_420_), .Y(_252__27_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(w_C_28_), .Y(_424_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_425_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_426_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_426_), .C(_425_), .Y(_427_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_421_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_422_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_422_), .C(w_C_28_), .Y(_423_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_427_), .Y(_252__28_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(w_C_29_), .Y(_431_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_432_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_433_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_433_), .C(_432_), .Y(_434_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_428_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_429_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_429_), .C(w_C_29_), .Y(_430_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_434_), .Y(_252__29_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(w_C_30_), .Y(_438_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_439_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_440_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_440_), .C(_439_), .Y(_441_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_435_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_436_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_436_), .C(w_C_30_), .Y(_437_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_441_), .Y(_252__30_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(w_C_31_), .Y(_445_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_446_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_447_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_445_), .B(_447_), .C(_446_), .Y(_448_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_442_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_443_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_443_), .C(w_C_31_), .Y(_444_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_448_), .Y(_252__31_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(w_C_32_), .Y(_452_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_453_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_454_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_454_), .C(_453_), .Y(_455_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_449_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_450_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_450_), .C(w_C_32_), .Y(_451_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_455_), .Y(_252__32_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(w_C_33_), .Y(_459_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_460_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_461_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_461_), .C(_460_), .Y(_462_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_456_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_457_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_456_), .B(_457_), .C(w_C_33_), .Y(_458_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_462_), .Y(_252__33_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(w_C_34_), .Y(_466_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_467_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_468_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_466_), .B(_468_), .C(_467_), .Y(_469_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_463_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_464_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_464_), .C(w_C_34_), .Y(_465_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_469_), .Y(_252__34_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(w_C_35_), .Y(_473_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_474_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_475_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_475_), .C(_474_), .Y(_476_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_470_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_471_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_470_), .B(_471_), .C(w_C_35_), .Y(_472_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_476_), .Y(_252__35_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(w_C_36_), .Y(_480_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_481_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_482_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_482_), .C(_481_), .Y(_483_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_477_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_478_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_477_), .B(_478_), .C(w_C_36_), .Y(_479_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_483_), .Y(_252__36_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(w_C_37_), .Y(_487_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_488_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_489_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_489_), .C(_488_), .Y(_490_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_484_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_485_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_484_), .B(_485_), .C(w_C_37_), .Y(_486_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_490_), .Y(_252__37_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(w_C_38_), .Y(_494_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_495_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_496_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_496_), .C(_495_), .Y(_497_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_491_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_492_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_492_), .C(w_C_38_), .Y(_493_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_497_), .Y(_252__38_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(w_C_39_), .Y(_501_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_502_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_503_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_501_), .B(_503_), .C(_502_), .Y(_504_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_498_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_499_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_499_), .C(w_C_39_), .Y(_500_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_504_), .Y(_252__39_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(w_C_40_), .Y(_508_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_509_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_510_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_510_), .C(_509_), .Y(_511_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_505_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_506_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(_506_), .C(w_C_40_), .Y(_507_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_511_), .Y(_252__40_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(w_C_41_), .Y(_515_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_516_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_517_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_517_), .C(_516_), .Y(_518_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_512_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_513_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_513_), .C(w_C_41_), .Y(_514_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_518_), .Y(_252__41_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(w_C_42_), .Y(_522_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_523_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_524_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_522_), .B(_524_), .C(_523_), .Y(_525_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_519_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_520_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_520_), .C(w_C_42_), .Y(_521_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_525_), .Y(_252__42_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_529_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_530_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_531_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_531_), .C(_530_), .Y(_532_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_526_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_527_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_527_), .C(gnd), .Y(_528_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_532_), .Y(_252__0_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_536_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_537_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_538_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_536_), .B(_538_), .C(_537_), .Y(_539_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_533_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_534_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_534_), .C(w_C_1_), .Y(_535_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_539_), .Y(_252__1_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_543_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_544_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_545_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_545_), .C(_544_), .Y(_546_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_540_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_541_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_541_), .C(w_C_2_), .Y(_542_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_542_), .B(_546_), .Y(_252__2_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_550_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_551_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_552_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_550_), .B(_552_), .C(_551_), .Y(_553_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_547_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_548_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_548_), .C(w_C_3_), .Y(_549_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(_553_), .Y(_252__3_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_7_), .Y(w_C_3_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .Y(_8_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add1[3]), .Y(_9_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_9_), .Y(_10_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_11_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_11_), .C(_7_), .Y(_12_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_10_), .Y(w_C_4_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_14_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_14_), .C(_12_), .Y(_15_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_15_), .Y(w_C_5_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_16_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_16_), .C(_15_), .Y(_17_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .C(_17_), .Y(_18_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_18_), .Y(w_C_6_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .Y(_19_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add1[6]), .Y(_20_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_21_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_21_), .Y(_22_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_23_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_23_), .Y(_24_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_24_), .C(_17_), .Y(_25_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_20_), .C(_25_), .Y(w_C_7_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_20_), .Y(_26_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_26_), .Y(_27_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_28_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_28_), .Y(_29_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_29_), .C(_25_), .Y(_30_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .C(_30_), .Y(_31_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_31_), .Y(w_C_8_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .Y(_32_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add1[8]), .Y(_33_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_34_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_34_), .Y(_35_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_36_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_36_), .Y(_37_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_37_), .C(_30_), .Y(_38_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_33_), .C(_38_), .Y(w_C_9_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_33_), .Y(_39_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_39_), .Y(_40_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_41_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_41_), .Y(_42_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_42_), .C(_38_), .Y(_43_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .C(_43_), .Y(_44_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_44_), .Y(w_C_10_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .Y(_45_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add1[10]), .Y(_46_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_47_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_47_), .Y(_48_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_49_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_49_), .Y(_50_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_50_), .C(_43_), .Y(_51_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_46_), .C(_51_), .Y(w_C_11_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_46_), .Y(_52_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_52_), .Y(_53_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_54_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_54_), .Y(_55_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_55_), .C(_51_), .Y(_56_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .C(_56_), .Y(_57_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_57_), .Y(w_C_12_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .Y(_58_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add1[12]), .Y(_59_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_60_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_60_), .Y(_61_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_62_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_62_), .Y(_63_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_63_), .C(_56_), .Y(_64_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_59_), .C(_64_), .Y(w_C_13_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_59_), .Y(_65_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_65_), .Y(_66_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_67_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_67_), .Y(_68_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_68_), .C(_64_), .Y(_69_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .C(_69_), .Y(_70_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_70_), .Y(w_C_14_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .Y(_71_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add1[14]), .Y(_72_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_72_), .Y(_73_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_73_), .Y(_74_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_75_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_75_), .Y(_76_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_77_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(_78_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_78_), .C(_69_), .Y(_79_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_74_), .Y(_80_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_80_), .Y(w_C_15_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_81_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_81_), .Y(_82_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_82_), .C(_79_), .Y(_83_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .C(_83_), .Y(_84_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_84_), .Y(w_C_16_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .Y(_85_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add1[16]), .Y(_86_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_86_), .Y(_87_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(_87_), .Y(_88_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_89_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_89_), .Y(_90_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_91_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_91_), .Y(_92_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_92_), .C(_83_), .Y(_93_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_88_), .Y(_94_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_94_), .Y(w_C_17_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_95_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_95_), .Y(_96_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_96_), .C(_93_), .Y(_97_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .C(_97_), .Y(_98_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_98_), .Y(w_C_18_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .Y(_99_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add1[18]), .Y(_100_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_100_), .Y(_101_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_101_), .Y(_102_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_103_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_103_), .Y(_104_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_105_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_105_), .Y(_106_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_106_), .C(_97_), .Y(_107_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_102_), .Y(_108_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(_108_), .Y(w_C_19_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_109_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_109_), .Y(_110_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_110_), .C(_107_), .Y(_111_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .C(_111_), .Y(_112_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_112_), .Y(w_C_20_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .Y(_113_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add1[20]), .Y(_114_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_114_), .Y(_115_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(_115_), .Y(_116_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_117_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_117_), .Y(_118_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_119_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(_119_), .Y(_120_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_120_), .C(_111_), .Y(_121_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_116_), .Y(_122_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(_122_), .Y(w_C_21_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_123_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(_123_), .Y(_124_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_124_), .C(_121_), .Y(_125_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .C(_125_), .Y(_126_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_126_), .Y(w_C_22_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .Y(_127_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add1[22]), .Y(_128_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_128_), .Y(_129_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(_129_), .Y(_130_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_131_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(_131_), .Y(_132_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_133_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(_133_), .Y(_134_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_134_), .C(_125_), .Y(_135_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_130_), .Y(_136_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(_136_), .Y(w_C_23_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_137_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(_137_), .Y(_138_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_138_), .C(_135_), .Y(_139_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .C(_139_), .Y(_140_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(_140_), .Y(w_C_24_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .Y(_141_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add1[24]), .Y(_142_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_142_), .Y(_143_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_143_), .Y(_144_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_145_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_145_), .Y(_146_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_147_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_147_), .Y(_148_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_148_), .C(_139_), .Y(_149_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_144_), .Y(_150_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_150_), .Y(w_C_25_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_151_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_151_), .Y(_152_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_152_), .C(_149_), .Y(_153_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .C(_153_), .Y(_154_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(_154_), .Y(w_C_26_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .Y(_155_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(i_add1[26]), .Y(_156_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_156_), .Y(_157_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(_157_), .Y(_158_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_159_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(_159_), .Y(_160_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_161_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(_161_), .Y(_162_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_162_), .C(_153_), .Y(_163_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_158_), .Y(_164_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(_164_), .Y(w_C_27_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_165_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(_165_), .Y(_166_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_166_), .C(_163_), .Y(_167_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .C(_167_), .Y(_168_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(_168_), .Y(w_C_28_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .Y(_169_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(i_add1[28]), .Y(_170_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_170_), .Y(_171_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(_171_), .Y(_172_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_173_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(_173_), .Y(_174_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_175_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(_175_), .Y(_176_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_176_), .C(_167_), .Y(_177_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_172_), .Y(_178_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(_178_), .Y(w_C_29_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_179_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(_179_), .Y(_180_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_180_), .C(_177_), .Y(_181_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .C(_181_), .Y(_182_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(_182_), .Y(w_C_30_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .Y(_183_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(i_add1[30]), .Y(_184_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_184_), .Y(_185_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(_185_), .Y(_186_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_187_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(_187_), .Y(_188_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_189_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(_189_), .Y(_190_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_190_), .C(_181_), .Y(_191_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_186_), .Y(_192_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(_192_), .Y(w_C_31_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_193_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(_193_), .Y(_194_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_194_), .C(_191_), .Y(_195_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .C(_195_), .Y(_196_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(_196_), .Y(w_C_32_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .Y(_197_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(i_add1[32]), .Y(_198_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_198_), .Y(_199_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(_199_), .Y(_200_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_201_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(_201_), .Y(_202_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_203_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(_203_), .Y(_204_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_204_), .C(_195_), .Y(_205_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_200_), .Y(_206_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(_206_), .Y(w_C_33_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_207_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(_207_), .Y(_208_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_208_), .C(_205_), .Y(_209_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .C(_209_), .Y(_210_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(_210_), .Y(w_C_34_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_211_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_212_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_210_), .C(_211_), .Y(w_C_35_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_213_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_214_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(_214_), .Y(_215_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(_212_), .Y(_216_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_216_), .C(_209_), .Y(_217_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_218_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_218_), .C(_217_), .Y(_219_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_213_), .Y(w_C_36_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .Y(_220_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(i_add1[36]), .Y(_221_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_221_), .Y(_222_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_222_), .C(_219_), .Y(_223_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_221_), .C(_223_), .Y(w_C_37_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .Y(_224_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(i_add1[37]), .Y(_225_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .C(w_C_37_), .Y(_226_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_225_), .C(_226_), .Y(w_C_38_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .Y(_227_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(i_add1[38]), .Y(_228_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_228_), .Y(_229_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(w_C_38_), .B(_229_), .Y(_230_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .C(_230_), .Y(_231_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(_231_), .Y(w_C_39_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_232_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_233_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_231_), .C(_232_), .Y(w_C_40_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_234_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(_233_), .Y(_235_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(_229_), .Y(_236_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_225_), .Y(_237_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_238_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_239_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_238_), .B(_239_), .C(_223_), .Y(_240_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_228_), .Y(_241_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_241_), .C(_240_), .Y(_242_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_232_), .C(_242_), .Y(_243_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_244_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_244_), .C(_243_), .Y(_245_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_245_), .Y(w_C_41_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_246_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_247_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_247_), .C(_245_), .Y(_248_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_246_), .Y(w_C_42_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_249_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_250_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_250_), .C(_248_), .Y(_251_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_251_), .Y(w_C_43_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_252__19_), .Y(o_result[19]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_252__20_), .Y(o_result[20]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_252__21_), .Y(o_result[21]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_252__22_), .Y(o_result[22]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_252__23_), .Y(o_result[23]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_252__24_), .Y(o_result[24]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_252__25_), .Y(o_result[25]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_252__26_), .Y(o_result[26]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_252__27_), .Y(o_result[27]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_252__28_), .Y(o_result[28]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_252__29_), .Y(o_result[29]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_252__30_), .Y(o_result[30]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_252__31_), .Y(o_result[31]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_252__32_), .Y(o_result[32]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_252__33_), .Y(o_result[33]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_252__34_), .Y(o_result[34]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_252__35_), .Y(o_result[35]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_252__36_), .Y(o_result[36]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_252__37_), .Y(o_result[37]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_252__38_), .Y(o_result[38]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_252__39_), .Y(o_result[39]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_252__40_), .Y(o_result[40]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_252__41_), .Y(o_result[41]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_252__42_), .Y(o_result[42]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(w_C_43_), .Y(o_result[43]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_252__0_), .Y(o_result[0]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_252__1_), .Y(o_result[1]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_252__2_), .Y(o_result[2]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_252__3_), .Y(o_result[3]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_252__4_), .Y(o_result[4]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_252__5_), .Y(o_result[5]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_252__6_), .Y(o_result[6]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_252__7_), .Y(o_result[7]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_252__8_), .Y(o_result[8]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_252__9_), .Y(o_result[9]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_252__10_), .Y(o_result[10]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_252__11_), .Y(o_result[11]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_252__12_), .Y(o_result[12]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_252__13_), .Y(o_result[13]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_252__14_), .Y(o_result[14]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_252__15_), .Y(o_result[15]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_252__16_), .Y(o_result[16]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_252__17_), .Y(o_result[17]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_252__18_), .Y(o_result[18]) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_256_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_257_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_258_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_258_), .C(_257_), .Y(_259_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_253_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_254_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_253_), .B(_254_), .C(w_C_4_), .Y(_255_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_259_), .Y(_252__4_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_263_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_264_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_265_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_265_), .C(_264_), .Y(_266_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_260_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_261_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_261_), .C(w_C_5_), .Y(_262_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_266_), .Y(_252__5_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_270_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_271_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_272_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_272_), .C(_271_), .Y(_273_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_267_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_268_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_268_), .C(w_C_6_), .Y(_269_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_273_), .Y(_252__6_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_277_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_278_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_279_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_279_), .C(_278_), .Y(_280_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_274_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_275_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_275_), .C(w_C_7_), .Y(_276_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_280_), .Y(_252__7_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_284_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_285_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_286_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_286_), .C(_285_), .Y(_287_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_281_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_282_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_282_), .C(w_C_8_), .Y(_283_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_283_), .B(_287_), .Y(_252__8_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_291_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_292_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_293_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_293_), .C(_292_), .Y(_294_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_288_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_289_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_289_), .C(w_C_9_), .Y(_290_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_294_), .Y(_252__9_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_298_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_299_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_300_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_300_), .C(_299_), .Y(_301_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_295_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_296_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_296_), .C(w_C_10_), .Y(_297_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_301_), .Y(_252__10_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_305_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_306_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_307_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_307_), .C(_306_), .Y(_308_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_302_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_303_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_303_), .C(w_C_11_), .Y(_304_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_308_), .Y(_252__11_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(w_C_12_), .Y(_312_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_313_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_314_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_314_), .C(_313_), .Y(_315_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_309_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_310_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_310_), .C(w_C_12_), .Y(_311_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_315_), .Y(_252__12_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(w_C_13_), .Y(_319_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_320_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_321_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_321_), .C(_320_), .Y(_322_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_316_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_317_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_316_), .B(_317_), .C(w_C_13_), .Y(_318_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_322_), .Y(_252__13_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(w_C_14_), .Y(_326_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_327_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_328_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_328_), .C(_327_), .Y(_329_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_323_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_324_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_324_), .C(w_C_14_), .Y(_325_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_329_), .Y(_252__14_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(_333_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_334_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_335_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_335_), .C(_334_), .Y(_336_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_330_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_331_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_331_), .C(w_C_15_), .Y(_332_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_336_), .Y(_252__15_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(w_C_16_), .Y(_340_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_341_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_342_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_342_), .C(_341_), .Y(_343_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_337_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_338_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_338_), .C(w_C_16_), .Y(_339_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_343_), .Y(_252__16_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(w_C_17_), .Y(_347_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_348_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_349_) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(w_C_43_), .Y(_252__43_) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
