module CSkipA_40bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_9_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_19_) );
OAI21X1 OAI21X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .C(1'b0), .Y(_20_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_21_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_22_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_23_) );
NAND3X1 NAND3X1_1 ( .A(_21_), .B(_22_), .C(_23_), .Y(_24_) );
OAI21X1 OAI21X1_2 ( .A(_20_), .B(_24_), .C(_19_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3_), .Y(_25_) );
OAI21X1 OAI21X1_3 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .C(1'b0), .Y(_26_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_27_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_28_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_29_) );
NAND3X1 NAND3X1_2 ( .A(_27_), .B(_28_), .C(_29_), .Y(_30_) );
OAI21X1 OAI21X1_4 ( .A(_26_), .B(_30_), .C(_25_), .Y(w_cout_2_) );
INVX1 INVX1_3 ( .A(_5_), .Y(_31_) );
OAI21X1 OAI21X1_5 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .C(1'b0), .Y(_32_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_33_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_34_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_35_) );
NAND3X1 NAND3X1_3 ( .A(_33_), .B(_34_), .C(_35_), .Y(_36_) );
OAI21X1 OAI21X1_6 ( .A(_32_), .B(_36_), .C(_31_), .Y(w_cout_3_) );
INVX1 INVX1_4 ( .A(_7_), .Y(_37_) );
OAI21X1 OAI21X1_7 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .C(1'b0), .Y(_38_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_39_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_40_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_41_) );
NAND3X1 NAND3X1_4 ( .A(_39_), .B(_40_), .C(_41_), .Y(_42_) );
OAI21X1 OAI21X1_8 ( .A(_38_), .B(_42_), .C(_37_), .Y(w_cout_4_) );
INVX1 INVX1_5 ( .A(_9_), .Y(_43_) );
OAI21X1 OAI21X1_9 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .C(1'b0), .Y(_44_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_45_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_46_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_47_) );
NAND3X1 NAND3X1_5 ( .A(_45_), .B(_46_), .C(_47_), .Y(_48_) );
OAI21X1 OAI21X1_10 ( .A(_44_), .B(_48_), .C(_43_), .Y(w_cout_5_) );
INVX1 INVX1_6 ( .A(_11_), .Y(_49_) );
OAI21X1 OAI21X1_11 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .C(1'b0), .Y(_50_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_51_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_52_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_53_) );
NAND3X1 NAND3X1_6 ( .A(_51_), .B(_52_), .C(_53_), .Y(_54_) );
OAI21X1 OAI21X1_12 ( .A(_50_), .B(_54_), .C(_49_), .Y(w_cout_6_) );
INVX1 INVX1_7 ( .A(_13_), .Y(_55_) );
OAI21X1 OAI21X1_13 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .C(1'b0), .Y(_56_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_57_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_58_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_59_) );
NAND3X1 NAND3X1_7 ( .A(_57_), .B(_58_), .C(_59_), .Y(_60_) );
OAI21X1 OAI21X1_14 ( .A(_56_), .B(_60_), .C(_55_), .Y(w_cout_7_) );
INVX1 INVX1_8 ( .A(_15_), .Y(_61_) );
OAI21X1 OAI21X1_15 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .C(1'b0), .Y(_62_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_63_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_64_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_65_) );
NAND3X1 NAND3X1_8 ( .A(_63_), .B(_64_), .C(_65_), .Y(_66_) );
OAI21X1 OAI21X1_16 ( .A(_62_), .B(_66_), .C(_61_), .Y(w_cout_8_) );
INVX1 INVX1_9 ( .A(_17_), .Y(_67_) );
OAI21X1 OAI21X1_17 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .C(1'b0), .Y(_68_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_69_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_70_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_71_) );
NAND3X1 NAND3X1_9 ( .A(_69_), .B(_70_), .C(_71_), .Y(_72_) );
OAI21X1 OAI21X1_18 ( .A(_68_), .B(_72_), .C(_67_), .Y(w_cout_9_) );
INVX1 INVX1_10 ( .A(skip0_cin_next), .Y(_76_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_77_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_78_) );
NAND3X1 NAND3X1_10 ( .A(_76_), .B(_78_), .C(_77_), .Y(_79_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_73_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_74_) );
OAI21X1 OAI21X1_19 ( .A(_73_), .B(_74_), .C(skip0_cin_next), .Y(_75_) );
NAND2X1 NAND2X1_2 ( .A(_75_), .B(_79_), .Y(_0__4_) );
OAI21X1 OAI21X1_20 ( .A(_76_), .B(_73_), .C(_78_), .Y(_2__1_) );
INVX1 INVX1_11 ( .A(_2__1_), .Y(_83_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_84_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_85_) );
NAND3X1 NAND3X1_11 ( .A(_83_), .B(_85_), .C(_84_), .Y(_86_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_80_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_81_) );
OAI21X1 OAI21X1_21 ( .A(_80_), .B(_81_), .C(_2__1_), .Y(_82_) );
NAND2X1 NAND2X1_4 ( .A(_82_), .B(_86_), .Y(_0__5_) );
OAI21X1 OAI21X1_22 ( .A(_83_), .B(_80_), .C(_85_), .Y(_2__2_) );
INVX1 INVX1_12 ( .A(_2__2_), .Y(_90_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_91_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_92_) );
NAND3X1 NAND3X1_12 ( .A(_90_), .B(_92_), .C(_91_), .Y(_93_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_87_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_88_) );
OAI21X1 OAI21X1_23 ( .A(_87_), .B(_88_), .C(_2__2_), .Y(_89_) );
NAND2X1 NAND2X1_6 ( .A(_89_), .B(_93_), .Y(_0__6_) );
OAI21X1 OAI21X1_24 ( .A(_90_), .B(_87_), .C(_92_), .Y(_2__3_) );
INVX1 INVX1_13 ( .A(_2__3_), .Y(_97_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_98_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_99_) );
NAND3X1 NAND3X1_13 ( .A(_97_), .B(_99_), .C(_98_), .Y(_100_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_94_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_95_) );
OAI21X1 OAI21X1_25 ( .A(_94_), .B(_95_), .C(_2__3_), .Y(_96_) );
NAND2X1 NAND2X1_8 ( .A(_96_), .B(_100_), .Y(_0__7_) );
OAI21X1 OAI21X1_26 ( .A(_97_), .B(_94_), .C(_99_), .Y(_1_) );
INVX1 INVX1_14 ( .A(w_cout_1_), .Y(_104_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_105_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_106_) );
NAND3X1 NAND3X1_14 ( .A(_104_), .B(_106_), .C(_105_), .Y(_107_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_101_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_102_) );
OAI21X1 OAI21X1_27 ( .A(_101_), .B(_102_), .C(w_cout_1_), .Y(_103_) );
NAND2X1 NAND2X1_10 ( .A(_103_), .B(_107_), .Y(_0__8_) );
OAI21X1 OAI21X1_28 ( .A(_104_), .B(_101_), .C(_106_), .Y(_4__1_) );
INVX1 INVX1_15 ( .A(_4__1_), .Y(_111_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_112_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_113_) );
NAND3X1 NAND3X1_15 ( .A(_111_), .B(_113_), .C(_112_), .Y(_114_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_108_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_109_) );
OAI21X1 OAI21X1_29 ( .A(_108_), .B(_109_), .C(_4__1_), .Y(_110_) );
NAND2X1 NAND2X1_12 ( .A(_110_), .B(_114_), .Y(_0__9_) );
OAI21X1 OAI21X1_30 ( .A(_111_), .B(_108_), .C(_113_), .Y(_4__2_) );
INVX1 INVX1_16 ( .A(_4__2_), .Y(_118_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_119_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_120_) );
NAND3X1 NAND3X1_16 ( .A(_118_), .B(_120_), .C(_119_), .Y(_121_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_115_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_116_) );
OAI21X1 OAI21X1_31 ( .A(_115_), .B(_116_), .C(_4__2_), .Y(_117_) );
NAND2X1 NAND2X1_14 ( .A(_117_), .B(_121_), .Y(_0__10_) );
OAI21X1 OAI21X1_32 ( .A(_118_), .B(_115_), .C(_120_), .Y(_4__3_) );
INVX1 INVX1_17 ( .A(_4__3_), .Y(_125_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_126_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_127_) );
NAND3X1 NAND3X1_17 ( .A(_125_), .B(_127_), .C(_126_), .Y(_128_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_122_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_123_) );
OAI21X1 OAI21X1_33 ( .A(_122_), .B(_123_), .C(_4__3_), .Y(_124_) );
NAND2X1 NAND2X1_16 ( .A(_124_), .B(_128_), .Y(_0__11_) );
OAI21X1 OAI21X1_34 ( .A(_125_), .B(_122_), .C(_127_), .Y(_3_) );
INVX1 INVX1_18 ( .A(w_cout_2_), .Y(_132_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_133_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_134_) );
NAND3X1 NAND3X1_18 ( .A(_132_), .B(_134_), .C(_133_), .Y(_135_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_129_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_130_) );
OAI21X1 OAI21X1_35 ( .A(_129_), .B(_130_), .C(w_cout_2_), .Y(_131_) );
NAND2X1 NAND2X1_18 ( .A(_131_), .B(_135_), .Y(_0__12_) );
OAI21X1 OAI21X1_36 ( .A(_132_), .B(_129_), .C(_134_), .Y(_6__1_) );
INVX1 INVX1_19 ( .A(_6__1_), .Y(_139_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_140_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_141_) );
NAND3X1 NAND3X1_19 ( .A(_139_), .B(_141_), .C(_140_), .Y(_142_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_136_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_137_) );
OAI21X1 OAI21X1_37 ( .A(_136_), .B(_137_), .C(_6__1_), .Y(_138_) );
NAND2X1 NAND2X1_20 ( .A(_138_), .B(_142_), .Y(_0__13_) );
OAI21X1 OAI21X1_38 ( .A(_139_), .B(_136_), .C(_141_), .Y(_6__2_) );
INVX1 INVX1_20 ( .A(_6__2_), .Y(_146_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_147_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_148_) );
NAND3X1 NAND3X1_20 ( .A(_146_), .B(_148_), .C(_147_), .Y(_149_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_143_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_144_) );
OAI21X1 OAI21X1_39 ( .A(_143_), .B(_144_), .C(_6__2_), .Y(_145_) );
NAND2X1 NAND2X1_22 ( .A(_145_), .B(_149_), .Y(_0__14_) );
OAI21X1 OAI21X1_40 ( .A(_146_), .B(_143_), .C(_148_), .Y(_6__3_) );
INVX1 INVX1_21 ( .A(_6__3_), .Y(_153_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_154_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_155_) );
NAND3X1 NAND3X1_21 ( .A(_153_), .B(_155_), .C(_154_), .Y(_156_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_150_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_151_) );
OAI21X1 OAI21X1_41 ( .A(_150_), .B(_151_), .C(_6__3_), .Y(_152_) );
NAND2X1 NAND2X1_24 ( .A(_152_), .B(_156_), .Y(_0__15_) );
OAI21X1 OAI21X1_42 ( .A(_153_), .B(_150_), .C(_155_), .Y(_5_) );
INVX1 INVX1_22 ( .A(w_cout_3_), .Y(_160_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_161_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_162_) );
NAND3X1 NAND3X1_22 ( .A(_160_), .B(_162_), .C(_161_), .Y(_163_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_157_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_158_) );
OAI21X1 OAI21X1_43 ( .A(_157_), .B(_158_), .C(w_cout_3_), .Y(_159_) );
NAND2X1 NAND2X1_26 ( .A(_159_), .B(_163_), .Y(_0__16_) );
OAI21X1 OAI21X1_44 ( .A(_160_), .B(_157_), .C(_162_), .Y(_8__1_) );
INVX1 INVX1_23 ( .A(_8__1_), .Y(_167_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_168_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_169_) );
NAND3X1 NAND3X1_23 ( .A(_167_), .B(_169_), .C(_168_), .Y(_170_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_164_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_165_) );
OAI21X1 OAI21X1_45 ( .A(_164_), .B(_165_), .C(_8__1_), .Y(_166_) );
NAND2X1 NAND2X1_28 ( .A(_166_), .B(_170_), .Y(_0__17_) );
OAI21X1 OAI21X1_46 ( .A(_167_), .B(_164_), .C(_169_), .Y(_8__2_) );
INVX1 INVX1_24 ( .A(_8__2_), .Y(_174_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_175_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_176_) );
NAND3X1 NAND3X1_24 ( .A(_174_), .B(_176_), .C(_175_), .Y(_177_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_171_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_172_) );
OAI21X1 OAI21X1_47 ( .A(_171_), .B(_172_), .C(_8__2_), .Y(_173_) );
NAND2X1 NAND2X1_30 ( .A(_173_), .B(_177_), .Y(_0__18_) );
OAI21X1 OAI21X1_48 ( .A(_174_), .B(_171_), .C(_176_), .Y(_8__3_) );
INVX1 INVX1_25 ( .A(_8__3_), .Y(_181_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_182_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_183_) );
NAND3X1 NAND3X1_25 ( .A(_181_), .B(_183_), .C(_182_), .Y(_184_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_178_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_179_) );
OAI21X1 OAI21X1_49 ( .A(_178_), .B(_179_), .C(_8__3_), .Y(_180_) );
NAND2X1 NAND2X1_32 ( .A(_180_), .B(_184_), .Y(_0__19_) );
OAI21X1 OAI21X1_50 ( .A(_181_), .B(_178_), .C(_183_), .Y(_7_) );
INVX1 INVX1_26 ( .A(w_cout_4_), .Y(_188_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_189_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_190_) );
NAND3X1 NAND3X1_26 ( .A(_188_), .B(_190_), .C(_189_), .Y(_191_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_185_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_186_) );
OAI21X1 OAI21X1_51 ( .A(_185_), .B(_186_), .C(w_cout_4_), .Y(_187_) );
NAND2X1 NAND2X1_34 ( .A(_187_), .B(_191_), .Y(_0__20_) );
OAI21X1 OAI21X1_52 ( .A(_188_), .B(_185_), .C(_190_), .Y(_10__1_) );
INVX1 INVX1_27 ( .A(_10__1_), .Y(_195_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_196_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_197_) );
NAND3X1 NAND3X1_27 ( .A(_195_), .B(_197_), .C(_196_), .Y(_198_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_192_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_193_) );
OAI21X1 OAI21X1_53 ( .A(_192_), .B(_193_), .C(_10__1_), .Y(_194_) );
NAND2X1 NAND2X1_36 ( .A(_194_), .B(_198_), .Y(_0__21_) );
OAI21X1 OAI21X1_54 ( .A(_195_), .B(_192_), .C(_197_), .Y(_10__2_) );
INVX1 INVX1_28 ( .A(_10__2_), .Y(_202_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_203_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_204_) );
NAND3X1 NAND3X1_28 ( .A(_202_), .B(_204_), .C(_203_), .Y(_205_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_199_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_200_) );
OAI21X1 OAI21X1_55 ( .A(_199_), .B(_200_), .C(_10__2_), .Y(_201_) );
NAND2X1 NAND2X1_38 ( .A(_201_), .B(_205_), .Y(_0__22_) );
OAI21X1 OAI21X1_56 ( .A(_202_), .B(_199_), .C(_204_), .Y(_10__3_) );
INVX1 INVX1_29 ( .A(_10__3_), .Y(_209_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_210_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_211_) );
NAND3X1 NAND3X1_29 ( .A(_209_), .B(_211_), .C(_210_), .Y(_212_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_206_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_207_) );
OAI21X1 OAI21X1_57 ( .A(_206_), .B(_207_), .C(_10__3_), .Y(_208_) );
NAND2X1 NAND2X1_40 ( .A(_208_), .B(_212_), .Y(_0__23_) );
OAI21X1 OAI21X1_58 ( .A(_209_), .B(_206_), .C(_211_), .Y(_9_) );
INVX1 INVX1_30 ( .A(w_cout_5_), .Y(_216_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_217_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_218_) );
NAND3X1 NAND3X1_30 ( .A(_216_), .B(_218_), .C(_217_), .Y(_219_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_213_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_214_) );
OAI21X1 OAI21X1_59 ( .A(_213_), .B(_214_), .C(w_cout_5_), .Y(_215_) );
NAND2X1 NAND2X1_42 ( .A(_215_), .B(_219_), .Y(_0__24_) );
OAI21X1 OAI21X1_60 ( .A(_216_), .B(_213_), .C(_218_), .Y(_12__1_) );
INVX1 INVX1_31 ( .A(_12__1_), .Y(_223_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_224_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_225_) );
NAND3X1 NAND3X1_31 ( .A(_223_), .B(_225_), .C(_224_), .Y(_226_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_220_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_221_) );
OAI21X1 OAI21X1_61 ( .A(_220_), .B(_221_), .C(_12__1_), .Y(_222_) );
NAND2X1 NAND2X1_44 ( .A(_222_), .B(_226_), .Y(_0__25_) );
OAI21X1 OAI21X1_62 ( .A(_223_), .B(_220_), .C(_225_), .Y(_12__2_) );
INVX1 INVX1_32 ( .A(_12__2_), .Y(_230_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_231_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_232_) );
NAND3X1 NAND3X1_32 ( .A(_230_), .B(_232_), .C(_231_), .Y(_233_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_227_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_228_) );
OAI21X1 OAI21X1_63 ( .A(_227_), .B(_228_), .C(_12__2_), .Y(_229_) );
NAND2X1 NAND2X1_46 ( .A(_229_), .B(_233_), .Y(_0__26_) );
OAI21X1 OAI21X1_64 ( .A(_230_), .B(_227_), .C(_232_), .Y(_12__3_) );
INVX1 INVX1_33 ( .A(_12__3_), .Y(_237_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_238_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_239_) );
NAND3X1 NAND3X1_33 ( .A(_237_), .B(_239_), .C(_238_), .Y(_240_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_234_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_235_) );
OAI21X1 OAI21X1_65 ( .A(_234_), .B(_235_), .C(_12__3_), .Y(_236_) );
NAND2X1 NAND2X1_48 ( .A(_236_), .B(_240_), .Y(_0__27_) );
OAI21X1 OAI21X1_66 ( .A(_237_), .B(_234_), .C(_239_), .Y(_11_) );
INVX1 INVX1_34 ( .A(w_cout_6_), .Y(_244_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_245_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_246_) );
NAND3X1 NAND3X1_34 ( .A(_244_), .B(_246_), .C(_245_), .Y(_247_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_241_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_242_) );
OAI21X1 OAI21X1_67 ( .A(_241_), .B(_242_), .C(w_cout_6_), .Y(_243_) );
NAND2X1 NAND2X1_50 ( .A(_243_), .B(_247_), .Y(_0__28_) );
OAI21X1 OAI21X1_68 ( .A(_244_), .B(_241_), .C(_246_), .Y(_14__1_) );
INVX1 INVX1_35 ( .A(_14__1_), .Y(_251_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_252_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_253_) );
NAND3X1 NAND3X1_35 ( .A(_251_), .B(_253_), .C(_252_), .Y(_254_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_248_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_249_) );
OAI21X1 OAI21X1_69 ( .A(_248_), .B(_249_), .C(_14__1_), .Y(_250_) );
NAND2X1 NAND2X1_52 ( .A(_250_), .B(_254_), .Y(_0__29_) );
OAI21X1 OAI21X1_70 ( .A(_251_), .B(_248_), .C(_253_), .Y(_14__2_) );
INVX1 INVX1_36 ( .A(_14__2_), .Y(_258_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_259_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_260_) );
NAND3X1 NAND3X1_36 ( .A(_258_), .B(_260_), .C(_259_), .Y(_261_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_255_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_256_) );
OAI21X1 OAI21X1_71 ( .A(_255_), .B(_256_), .C(_14__2_), .Y(_257_) );
NAND2X1 NAND2X1_54 ( .A(_257_), .B(_261_), .Y(_0__30_) );
OAI21X1 OAI21X1_72 ( .A(_258_), .B(_255_), .C(_260_), .Y(_14__3_) );
INVX1 INVX1_37 ( .A(_14__3_), .Y(_265_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_266_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_267_) );
NAND3X1 NAND3X1_37 ( .A(_265_), .B(_267_), .C(_266_), .Y(_268_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_262_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_263_) );
OAI21X1 OAI21X1_73 ( .A(_262_), .B(_263_), .C(_14__3_), .Y(_264_) );
NAND2X1 NAND2X1_56 ( .A(_264_), .B(_268_), .Y(_0__31_) );
OAI21X1 OAI21X1_74 ( .A(_265_), .B(_262_), .C(_267_), .Y(_13_) );
INVX1 INVX1_38 ( .A(w_cout_7_), .Y(_272_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_273_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_274_) );
NAND3X1 NAND3X1_38 ( .A(_272_), .B(_274_), .C(_273_), .Y(_275_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_269_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_270_) );
OAI21X1 OAI21X1_75 ( .A(_269_), .B(_270_), .C(w_cout_7_), .Y(_271_) );
NAND2X1 NAND2X1_58 ( .A(_271_), .B(_275_), .Y(_0__32_) );
OAI21X1 OAI21X1_76 ( .A(_272_), .B(_269_), .C(_274_), .Y(_16__1_) );
INVX1 INVX1_39 ( .A(_16__1_), .Y(_279_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_280_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_281_) );
NAND3X1 NAND3X1_39 ( .A(_279_), .B(_281_), .C(_280_), .Y(_282_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_276_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_277_) );
OAI21X1 OAI21X1_77 ( .A(_276_), .B(_277_), .C(_16__1_), .Y(_278_) );
NAND2X1 NAND2X1_60 ( .A(_278_), .B(_282_), .Y(_0__33_) );
OAI21X1 OAI21X1_78 ( .A(_279_), .B(_276_), .C(_281_), .Y(_16__2_) );
INVX1 INVX1_40 ( .A(_16__2_), .Y(_286_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_287_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_288_) );
NAND3X1 NAND3X1_40 ( .A(_286_), .B(_288_), .C(_287_), .Y(_289_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_283_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_284_) );
OAI21X1 OAI21X1_79 ( .A(_283_), .B(_284_), .C(_16__2_), .Y(_285_) );
NAND2X1 NAND2X1_62 ( .A(_285_), .B(_289_), .Y(_0__34_) );
OAI21X1 OAI21X1_80 ( .A(_286_), .B(_283_), .C(_288_), .Y(_16__3_) );
INVX1 INVX1_41 ( .A(_16__3_), .Y(_293_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_294_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_295_) );
NAND3X1 NAND3X1_41 ( .A(_293_), .B(_295_), .C(_294_), .Y(_296_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_290_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_291_) );
OAI21X1 OAI21X1_81 ( .A(_290_), .B(_291_), .C(_16__3_), .Y(_292_) );
NAND2X1 NAND2X1_64 ( .A(_292_), .B(_296_), .Y(_0__35_) );
OAI21X1 OAI21X1_82 ( .A(_293_), .B(_290_), .C(_295_), .Y(_15_) );
INVX1 INVX1_42 ( .A(w_cout_8_), .Y(_300_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_301_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_302_) );
NAND3X1 NAND3X1_42 ( .A(_300_), .B(_302_), .C(_301_), .Y(_303_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_297_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_298_) );
OAI21X1 OAI21X1_83 ( .A(_297_), .B(_298_), .C(w_cout_8_), .Y(_299_) );
NAND2X1 NAND2X1_66 ( .A(_299_), .B(_303_), .Y(_0__36_) );
OAI21X1 OAI21X1_84 ( .A(_300_), .B(_297_), .C(_302_), .Y(_18__1_) );
INVX1 INVX1_43 ( .A(_18__1_), .Y(_307_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_308_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_309_) );
NAND3X1 NAND3X1_43 ( .A(_307_), .B(_309_), .C(_308_), .Y(_310_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_304_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_305_) );
OAI21X1 OAI21X1_85 ( .A(_304_), .B(_305_), .C(_18__1_), .Y(_306_) );
NAND2X1 NAND2X1_68 ( .A(_306_), .B(_310_), .Y(_0__37_) );
OAI21X1 OAI21X1_86 ( .A(_307_), .B(_304_), .C(_309_), .Y(_18__2_) );
INVX1 INVX1_44 ( .A(_18__2_), .Y(_314_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_315_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_316_) );
NAND3X1 NAND3X1_44 ( .A(_314_), .B(_316_), .C(_315_), .Y(_317_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_311_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_312_) );
OAI21X1 OAI21X1_87 ( .A(_311_), .B(_312_), .C(_18__2_), .Y(_313_) );
NAND2X1 NAND2X1_70 ( .A(_313_), .B(_317_), .Y(_0__38_) );
OAI21X1 OAI21X1_88 ( .A(_314_), .B(_311_), .C(_316_), .Y(_18__3_) );
INVX1 INVX1_45 ( .A(_18__3_), .Y(_321_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_322_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_323_) );
NAND3X1 NAND3X1_45 ( .A(_321_), .B(_323_), .C(_322_), .Y(_324_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_318_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_319_) );
OAI21X1 OAI21X1_89 ( .A(_318_), .B(_319_), .C(_18__3_), .Y(_320_) );
NAND2X1 NAND2X1_72 ( .A(_320_), .B(_324_), .Y(_0__39_) );
OAI21X1 OAI21X1_90 ( .A(_321_), .B(_318_), .C(_323_), .Y(_17_) );
INVX1 INVX1_46 ( .A(1'b0), .Y(_328_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_329_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_330_) );
NAND3X1 NAND3X1_46 ( .A(_328_), .B(_330_), .C(_329_), .Y(_331_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_325_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_326_) );
OAI21X1 OAI21X1_91 ( .A(_325_), .B(_326_), .C(1'b0), .Y(_327_) );
NAND2X1 NAND2X1_74 ( .A(_327_), .B(_331_), .Y(_0__0_) );
OAI21X1 OAI21X1_92 ( .A(_328_), .B(_325_), .C(_330_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_47 ( .A(rca_inst_w_CARRY_1_), .Y(_335_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_336_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_337_) );
NAND3X1 NAND3X1_47 ( .A(_335_), .B(_337_), .C(_336_), .Y(_338_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_332_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_333_) );
OAI21X1 OAI21X1_93 ( .A(_332_), .B(_333_), .C(rca_inst_w_CARRY_1_), .Y(_334_) );
NAND2X1 NAND2X1_76 ( .A(_334_), .B(_338_), .Y(_0__1_) );
OAI21X1 OAI21X1_94 ( .A(_335_), .B(_332_), .C(_337_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_48 ( .A(rca_inst_w_CARRY_2_), .Y(_342_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_343_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_344_) );
NAND3X1 NAND3X1_48 ( .A(_342_), .B(_344_), .C(_343_), .Y(_345_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_339_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_340_) );
OAI21X1 OAI21X1_95 ( .A(_339_), .B(_340_), .C(rca_inst_w_CARRY_2_), .Y(_341_) );
NAND2X1 NAND2X1_78 ( .A(_341_), .B(_345_), .Y(_0__2_) );
OAI21X1 OAI21X1_96 ( .A(_342_), .B(_339_), .C(_344_), .Y(rca_inst_w_CARRY_3_) );
INVX1 INVX1_49 ( .A(rca_inst_w_CARRY_3_), .Y(_349_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_350_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_351_) );
NAND3X1 NAND3X1_49 ( .A(_349_), .B(_351_), .C(_350_), .Y(_352_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_346_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_347_) );
OAI21X1 OAI21X1_97 ( .A(_346_), .B(_347_), .C(rca_inst_w_CARRY_3_), .Y(_348_) );
NAND2X1 NAND2X1_80 ( .A(_348_), .B(_352_), .Y(_0__3_) );
OAI21X1 OAI21X1_98 ( .A(_349_), .B(_346_), .C(_351_), .Y(cout0) );
INVX1 INVX1_50 ( .A(cout0), .Y(_353_) );
OAI21X1 OAI21X1_99 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .C(1'b0), .Y(_354_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_355_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_356_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_357_) );
NAND3X1 NAND3X1_50 ( .A(_355_), .B(_356_), .C(_357_), .Y(_358_) );
OAI21X1 OAI21X1_100 ( .A(_354_), .B(_358_), .C(_353_), .Y(skip0_cin_next) );
BUFX2 BUFX2_42 ( .A(skip0_cin_next), .Y(_2__0_) );
BUFX2 BUFX2_43 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_44 ( .A(w_cout_1_), .Y(_4__0_) );
BUFX2 BUFX2_45 ( .A(_3_), .Y(_4__4_) );
BUFX2 BUFX2_46 ( .A(w_cout_2_), .Y(_6__0_) );
BUFX2 BUFX2_47 ( .A(_5_), .Y(_6__4_) );
BUFX2 BUFX2_48 ( .A(w_cout_3_), .Y(_8__0_) );
BUFX2 BUFX2_49 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_50 ( .A(w_cout_4_), .Y(_10__0_) );
BUFX2 BUFX2_51 ( .A(_9_), .Y(_10__4_) );
BUFX2 BUFX2_52 ( .A(w_cout_5_), .Y(_12__0_) );
BUFX2 BUFX2_53 ( .A(_11_), .Y(_12__4_) );
BUFX2 BUFX2_54 ( .A(w_cout_6_), .Y(_14__0_) );
BUFX2 BUFX2_55 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_56 ( .A(w_cout_7_), .Y(_16__0_) );
BUFX2 BUFX2_57 ( .A(_15_), .Y(_16__4_) );
BUFX2 BUFX2_58 ( .A(w_cout_8_), .Y(_18__0_) );
BUFX2 BUFX2_59 ( .A(_17_), .Y(_18__4_) );
BUFX2 BUFX2_60 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_61 ( .A(cout0), .Y(rca_inst_w_CARRY_4_) );
BUFX2 BUFX2_62 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
