module CSkipA_21bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_6_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(cskip1_inst_rca0_fa0_o_sum), .Y(sum[20]) );
INVX1 INVX1_1 ( .A(1'b0), .Y(_19_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_20_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_21_) );
NAND3X1 NAND3X1_1 ( .A(_19_), .B(_21_), .C(_20_), .Y(_22_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_16_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_17_) );
OAI21X1 OAI21X1_1 ( .A(_16_), .B(_17_), .C(1'b0), .Y(_18_) );
NAND2X1 NAND2X1_2 ( .A(_18_), .B(_22_), .Y(_0__0_) );
OAI21X1 OAI21X1_2 ( .A(_19_), .B(_16_), .C(_21_), .Y(_2__1_) );
INVX1 INVX1_2 ( .A(_2__3_), .Y(_26_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_27_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_28_) );
NAND3X1 NAND3X1_2 ( .A(_26_), .B(_28_), .C(_27_), .Y(_29_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_23_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_24_) );
OAI21X1 OAI21X1_3 ( .A(_23_), .B(_24_), .C(_2__3_), .Y(_25_) );
NAND2X1 NAND2X1_4 ( .A(_25_), .B(_29_), .Y(_0__3_) );
OAI21X1 OAI21X1_4 ( .A(_26_), .B(_23_), .C(_28_), .Y(_1_) );
INVX1 INVX1_3 ( .A(_2__1_), .Y(_33_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_34_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_35_) );
NAND3X1 NAND3X1_3 ( .A(_33_), .B(_35_), .C(_34_), .Y(_36_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_30_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_31_) );
OAI21X1 OAI21X1_5 ( .A(_30_), .B(_31_), .C(_2__1_), .Y(_32_) );
NAND2X1 NAND2X1_6 ( .A(_32_), .B(_36_), .Y(_0__1_) );
OAI21X1 OAI21X1_6 ( .A(_33_), .B(_30_), .C(_35_), .Y(_2__2_) );
INVX1 INVX1_4 ( .A(_2__2_), .Y(_40_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_41_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_42_) );
NAND3X1 NAND3X1_4 ( .A(_40_), .B(_42_), .C(_41_), .Y(_43_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_37_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_38_) );
OAI21X1 OAI21X1_7 ( .A(_37_), .B(_38_), .C(_2__2_), .Y(_39_) );
NAND2X1 NAND2X1_8 ( .A(_39_), .B(_43_), .Y(_0__2_) );
OAI21X1 OAI21X1_8 ( .A(_40_), .B(_37_), .C(_42_), .Y(_2__3_) );
INVX1 INVX1_5 ( .A(i_add_term1[0]), .Y(_44_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[0]), .B(_44_), .Y(_45_) );
INVX1 INVX1_6 ( .A(i_add_term2[0]), .Y(_46_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term1[0]), .B(_46_), .Y(_47_) );
INVX1 INVX1_7 ( .A(i_add_term1[1]), .Y(_48_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[1]), .B(_48_), .Y(_49_) );
INVX1 INVX1_8 ( .A(i_add_term2[1]), .Y(_50_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term1[1]), .B(_50_), .Y(_51_) );
OAI22X1 OAI22X1_1 ( .A(_45_), .B(_47_), .C(_49_), .D(_51_), .Y(_52_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_53_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_54_) );
NOR2X1 NOR2X1_10 ( .A(_53_), .B(_54_), .Y(_55_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_56_) );
NAND2X1 NAND2X1_9 ( .A(_55_), .B(_56_), .Y(_57_) );
NOR2X1 NOR2X1_11 ( .A(_52_), .B(_57_), .Y(_3_) );
INVX1 INVX1_9 ( .A(_1_), .Y(_58_) );
NAND2X1 NAND2X1_10 ( .A(1'b0), .B(_3_), .Y(_59_) );
OAI21X1 OAI21X1_9 ( .A(_3_), .B(_58_), .C(_59_), .Y(w_cout_1_) );
INVX1 INVX1_10 ( .A(w_cout_1_), .Y(_63_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_64_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_65_) );
NAND3X1 NAND3X1_5 ( .A(_63_), .B(_65_), .C(_64_), .Y(_66_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_60_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_61_) );
OAI21X1 OAI21X1_10 ( .A(_60_), .B(_61_), .C(w_cout_1_), .Y(_62_) );
NAND2X1 NAND2X1_12 ( .A(_62_), .B(_66_), .Y(_0__4_) );
OAI21X1 OAI21X1_11 ( .A(_63_), .B(_60_), .C(_65_), .Y(_5__1_) );
INVX1 INVX1_11 ( .A(_5__3_), .Y(_70_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_71_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_72_) );
NAND3X1 NAND3X1_6 ( .A(_70_), .B(_72_), .C(_71_), .Y(_73_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_67_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_68_) );
OAI21X1 OAI21X1_12 ( .A(_67_), .B(_68_), .C(_5__3_), .Y(_69_) );
NAND2X1 NAND2X1_14 ( .A(_69_), .B(_73_), .Y(_0__7_) );
OAI21X1 OAI21X1_13 ( .A(_70_), .B(_67_), .C(_72_), .Y(_4_) );
INVX1 INVX1_12 ( .A(_5__1_), .Y(_77_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_78_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_79_) );
NAND3X1 NAND3X1_7 ( .A(_77_), .B(_79_), .C(_78_), .Y(_80_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_74_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_75_) );
OAI21X1 OAI21X1_14 ( .A(_74_), .B(_75_), .C(_5__1_), .Y(_76_) );
NAND2X1 NAND2X1_16 ( .A(_76_), .B(_80_), .Y(_0__5_) );
OAI21X1 OAI21X1_15 ( .A(_77_), .B(_74_), .C(_79_), .Y(_5__2_) );
INVX1 INVX1_13 ( .A(_5__2_), .Y(_84_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_85_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_86_) );
NAND3X1 NAND3X1_8 ( .A(_84_), .B(_86_), .C(_85_), .Y(_87_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_81_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_82_) );
OAI21X1 OAI21X1_16 ( .A(_81_), .B(_82_), .C(_5__2_), .Y(_83_) );
NAND2X1 NAND2X1_18 ( .A(_83_), .B(_87_), .Y(_0__6_) );
OAI21X1 OAI21X1_17 ( .A(_84_), .B(_81_), .C(_86_), .Y(_5__3_) );
INVX1 INVX1_14 ( .A(i_add_term1[4]), .Y(_88_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[4]), .B(_88_), .Y(_89_) );
INVX1 INVX1_15 ( .A(i_add_term2[4]), .Y(_90_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term1[4]), .B(_90_), .Y(_91_) );
INVX1 INVX1_16 ( .A(i_add_term1[5]), .Y(_92_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[5]), .B(_92_), .Y(_93_) );
INVX1 INVX1_17 ( .A(i_add_term2[5]), .Y(_94_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term1[5]), .B(_94_), .Y(_95_) );
OAI22X1 OAI22X1_2 ( .A(_89_), .B(_91_), .C(_93_), .D(_95_), .Y(_96_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_97_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_98_) );
NOR2X1 NOR2X1_21 ( .A(_97_), .B(_98_), .Y(_99_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_100_) );
NAND2X1 NAND2X1_19 ( .A(_99_), .B(_100_), .Y(_101_) );
NOR2X1 NOR2X1_22 ( .A(_96_), .B(_101_), .Y(_6_) );
INVX1 INVX1_18 ( .A(_4_), .Y(_102_) );
NAND2X1 NAND2X1_20 ( .A(1'b0), .B(_6_), .Y(_103_) );
OAI21X1 OAI21X1_18 ( .A(_6_), .B(_102_), .C(_103_), .Y(w_cout_2_) );
INVX1 INVX1_19 ( .A(w_cout_2_), .Y(_107_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_108_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_109_) );
NAND3X1 NAND3X1_9 ( .A(_107_), .B(_109_), .C(_108_), .Y(_110_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_104_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_105_) );
OAI21X1 OAI21X1_19 ( .A(_104_), .B(_105_), .C(w_cout_2_), .Y(_106_) );
NAND2X1 NAND2X1_22 ( .A(_106_), .B(_110_), .Y(_0__8_) );
OAI21X1 OAI21X1_20 ( .A(_107_), .B(_104_), .C(_109_), .Y(_8__1_) );
INVX1 INVX1_20 ( .A(_8__3_), .Y(_114_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_115_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_116_) );
NAND3X1 NAND3X1_10 ( .A(_114_), .B(_116_), .C(_115_), .Y(_117_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_111_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_112_) );
OAI21X1 OAI21X1_21 ( .A(_111_), .B(_112_), .C(_8__3_), .Y(_113_) );
NAND2X1 NAND2X1_24 ( .A(_113_), .B(_117_), .Y(_0__11_) );
OAI21X1 OAI21X1_22 ( .A(_114_), .B(_111_), .C(_116_), .Y(_7_) );
INVX1 INVX1_21 ( .A(_8__1_), .Y(_121_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_122_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_123_) );
NAND3X1 NAND3X1_11 ( .A(_121_), .B(_123_), .C(_122_), .Y(_124_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_118_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_119_) );
OAI21X1 OAI21X1_23 ( .A(_118_), .B(_119_), .C(_8__1_), .Y(_120_) );
NAND2X1 NAND2X1_26 ( .A(_120_), .B(_124_), .Y(_0__9_) );
OAI21X1 OAI21X1_24 ( .A(_121_), .B(_118_), .C(_123_), .Y(_8__2_) );
INVX1 INVX1_22 ( .A(_8__2_), .Y(_128_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_129_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_130_) );
NAND3X1 NAND3X1_12 ( .A(_128_), .B(_130_), .C(_129_), .Y(_131_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_125_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_126_) );
OAI21X1 OAI21X1_25 ( .A(_125_), .B(_126_), .C(_8__2_), .Y(_127_) );
NAND2X1 NAND2X1_28 ( .A(_127_), .B(_131_), .Y(_0__10_) );
OAI21X1 OAI21X1_26 ( .A(_128_), .B(_125_), .C(_130_), .Y(_8__3_) );
INVX1 INVX1_23 ( .A(i_add_term1[8]), .Y(_132_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[8]), .B(_132_), .Y(_133_) );
INVX1 INVX1_24 ( .A(i_add_term2[8]), .Y(_134_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term1[8]), .B(_134_), .Y(_135_) );
INVX1 INVX1_25 ( .A(i_add_term1[9]), .Y(_136_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[9]), .B(_136_), .Y(_137_) );
INVX1 INVX1_26 ( .A(i_add_term2[9]), .Y(_138_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term1[9]), .B(_138_), .Y(_139_) );
OAI22X1 OAI22X1_3 ( .A(_133_), .B(_135_), .C(_137_), .D(_139_), .Y(_140_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_141_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_142_) );
NOR2X1 NOR2X1_32 ( .A(_141_), .B(_142_), .Y(_143_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_144_) );
NAND2X1 NAND2X1_29 ( .A(_143_), .B(_144_), .Y(_145_) );
NOR2X1 NOR2X1_33 ( .A(_140_), .B(_145_), .Y(_9_) );
INVX1 INVX1_27 ( .A(_7_), .Y(_146_) );
NAND2X1 NAND2X1_30 ( .A(1'b0), .B(_9_), .Y(_147_) );
OAI21X1 OAI21X1_27 ( .A(_9_), .B(_146_), .C(_147_), .Y(w_cout_3_) );
INVX1 INVX1_28 ( .A(w_cout_3_), .Y(_151_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_152_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_153_) );
NAND3X1 NAND3X1_13 ( .A(_151_), .B(_153_), .C(_152_), .Y(_154_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_148_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_149_) );
OAI21X1 OAI21X1_28 ( .A(_148_), .B(_149_), .C(w_cout_3_), .Y(_150_) );
NAND2X1 NAND2X1_32 ( .A(_150_), .B(_154_), .Y(_0__12_) );
OAI21X1 OAI21X1_29 ( .A(_151_), .B(_148_), .C(_153_), .Y(_11__1_) );
INVX1 INVX1_29 ( .A(_11__3_), .Y(_158_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_159_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_160_) );
NAND3X1 NAND3X1_14 ( .A(_158_), .B(_160_), .C(_159_), .Y(_161_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_155_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_156_) );
OAI21X1 OAI21X1_30 ( .A(_155_), .B(_156_), .C(_11__3_), .Y(_157_) );
NAND2X1 NAND2X1_34 ( .A(_157_), .B(_161_), .Y(_0__15_) );
OAI21X1 OAI21X1_31 ( .A(_158_), .B(_155_), .C(_160_), .Y(_10_) );
INVX1 INVX1_30 ( .A(_11__1_), .Y(_165_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_166_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_167_) );
NAND3X1 NAND3X1_15 ( .A(_165_), .B(_167_), .C(_166_), .Y(_168_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_162_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_163_) );
OAI21X1 OAI21X1_32 ( .A(_162_), .B(_163_), .C(_11__1_), .Y(_164_) );
NAND2X1 NAND2X1_36 ( .A(_164_), .B(_168_), .Y(_0__13_) );
OAI21X1 OAI21X1_33 ( .A(_165_), .B(_162_), .C(_167_), .Y(_11__2_) );
INVX1 INVX1_31 ( .A(_11__2_), .Y(_172_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_173_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_174_) );
NAND3X1 NAND3X1_16 ( .A(_172_), .B(_174_), .C(_173_), .Y(_175_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_169_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_170_) );
OAI21X1 OAI21X1_34 ( .A(_169_), .B(_170_), .C(_11__2_), .Y(_171_) );
NAND2X1 NAND2X1_38 ( .A(_171_), .B(_175_), .Y(_0__14_) );
OAI21X1 OAI21X1_35 ( .A(_172_), .B(_169_), .C(_174_), .Y(_11__3_) );
INVX1 INVX1_32 ( .A(i_add_term1[12]), .Y(_176_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[12]), .B(_176_), .Y(_177_) );
INVX1 INVX1_33 ( .A(i_add_term2[12]), .Y(_178_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term1[12]), .B(_178_), .Y(_179_) );
INVX1 INVX1_34 ( .A(i_add_term1[13]), .Y(_180_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[13]), .B(_180_), .Y(_181_) );
INVX1 INVX1_35 ( .A(i_add_term2[13]), .Y(_182_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term1[13]), .B(_182_), .Y(_183_) );
OAI22X1 OAI22X1_4 ( .A(_177_), .B(_179_), .C(_181_), .D(_183_), .Y(_184_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_185_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_186_) );
NOR2X1 NOR2X1_43 ( .A(_185_), .B(_186_), .Y(_187_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_188_) );
NAND2X1 NAND2X1_39 ( .A(_187_), .B(_188_), .Y(_189_) );
NOR2X1 NOR2X1_44 ( .A(_184_), .B(_189_), .Y(_12_) );
INVX1 INVX1_36 ( .A(_10_), .Y(_190_) );
NAND2X1 NAND2X1_40 ( .A(1'b0), .B(_12_), .Y(_191_) );
OAI21X1 OAI21X1_36 ( .A(_12_), .B(_190_), .C(_191_), .Y(w_cout_4_) );
INVX1 INVX1_37 ( .A(w_cout_4_), .Y(_195_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_196_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_197_) );
NAND3X1 NAND3X1_17 ( .A(_195_), .B(_197_), .C(_196_), .Y(_198_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_192_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_193_) );
OAI21X1 OAI21X1_37 ( .A(_192_), .B(_193_), .C(w_cout_4_), .Y(_194_) );
NAND2X1 NAND2X1_42 ( .A(_194_), .B(_198_), .Y(_0__16_) );
OAI21X1 OAI21X1_38 ( .A(_195_), .B(_192_), .C(_197_), .Y(_14__1_) );
INVX1 INVX1_38 ( .A(_14__3_), .Y(_202_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_203_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_204_) );
NAND3X1 NAND3X1_18 ( .A(_202_), .B(_204_), .C(_203_), .Y(_205_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_199_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_200_) );
OAI21X1 OAI21X1_39 ( .A(_199_), .B(_200_), .C(_14__3_), .Y(_201_) );
NAND2X1 NAND2X1_44 ( .A(_201_), .B(_205_), .Y(_0__19_) );
OAI21X1 OAI21X1_40 ( .A(_202_), .B(_199_), .C(_204_), .Y(_13_) );
INVX1 INVX1_39 ( .A(_14__1_), .Y(_209_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_210_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_211_) );
NAND3X1 NAND3X1_19 ( .A(_209_), .B(_211_), .C(_210_), .Y(_212_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_206_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_207_) );
OAI21X1 OAI21X1_41 ( .A(_206_), .B(_207_), .C(_14__1_), .Y(_208_) );
NAND2X1 NAND2X1_46 ( .A(_208_), .B(_212_), .Y(_0__17_) );
OAI21X1 OAI21X1_42 ( .A(_209_), .B(_206_), .C(_211_), .Y(_14__2_) );
INVX1 INVX1_40 ( .A(_14__2_), .Y(_216_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_217_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_218_) );
NAND3X1 NAND3X1_20 ( .A(_216_), .B(_218_), .C(_217_), .Y(_219_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_213_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_214_) );
OAI21X1 OAI21X1_43 ( .A(_213_), .B(_214_), .C(_14__2_), .Y(_215_) );
NAND2X1 NAND2X1_48 ( .A(_215_), .B(_219_), .Y(_0__18_) );
OAI21X1 OAI21X1_44 ( .A(_216_), .B(_213_), .C(_218_), .Y(_14__3_) );
INVX1 INVX1_41 ( .A(i_add_term1[16]), .Y(_220_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[16]), .B(_220_), .Y(_221_) );
INVX1 INVX1_42 ( .A(i_add_term2[16]), .Y(_222_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term1[16]), .B(_222_), .Y(_223_) );
INVX1 INVX1_43 ( .A(i_add_term1[17]), .Y(_224_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[17]), .B(_224_), .Y(_225_) );
INVX1 INVX1_44 ( .A(i_add_term2[17]), .Y(_226_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term1[17]), .B(_226_), .Y(_227_) );
OAI22X1 OAI22X1_5 ( .A(_221_), .B(_223_), .C(_225_), .D(_227_), .Y(_228_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_229_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_230_) );
NOR2X1 NOR2X1_54 ( .A(_229_), .B(_230_), .Y(_231_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_232_) );
NAND2X1 NAND2X1_49 ( .A(_231_), .B(_232_), .Y(_233_) );
NOR2X1 NOR2X1_55 ( .A(_228_), .B(_233_), .Y(_15_) );
INVX1 INVX1_45 ( .A(_13_), .Y(_234_) );
NAND2X1 NAND2X1_50 ( .A(1'b0), .B(_15_), .Y(_235_) );
OAI21X1 OAI21X1_45 ( .A(_15_), .B(_234_), .C(_235_), .Y(cskip1_inst_cin) );
INVX1 INVX1_46 ( .A(cskip1_inst_cin), .Y(_239_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_240_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_241_) );
NAND3X1 NAND3X1_21 ( .A(_239_), .B(_241_), .C(_240_), .Y(_242_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_236_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_237_) );
OAI21X1 OAI21X1_46 ( .A(_236_), .B(_237_), .C(cskip1_inst_cin), .Y(_238_) );
NAND2X1 NAND2X1_52 ( .A(_238_), .B(_242_), .Y(cskip1_inst_rca0_fa0_o_sum) );
OAI21X1 OAI21X1_47 ( .A(_239_), .B(_236_), .C(_241_), .Y(cskip1_inst_cout0) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_243_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_244_) );
NOR2X1 NOR2X1_58 ( .A(_243_), .B(_244_), .Y(cskip1_inst_skip0_P) );
INVX1 INVX1_47 ( .A(cskip1_inst_cout0), .Y(_245_) );
NAND2X1 NAND2X1_53 ( .A(1'b0), .B(cskip1_inst_skip0_P), .Y(_246_) );
OAI21X1 OAI21X1_48 ( .A(cskip1_inst_skip0_P), .B(_245_), .C(_246_), .Y(w_cout_6_) );
BUFX2 BUFX2_23 ( .A(cskip1_inst_rca0_fa0_o_sum), .Y(_0__20_) );
BUFX2 BUFX2_24 ( .A(1'b0), .Y(w_cout_0_) );
BUFX2 BUFX2_25 ( .A(cskip1_inst_cin), .Y(w_cout_5_) );
endmodule
