module CSkipA_57bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term1[45], i_add_term1[46], i_add_term1[47], i_add_term1[48], i_add_term1[49], i_add_term1[50], i_add_term1[51], i_add_term1[52], i_add_term1[53], i_add_term1[54], i_add_term1[55], i_add_term1[56], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], i_add_term2[45], i_add_term2[46], i_add_term2[47], i_add_term2[48], i_add_term2[49], i_add_term2[50], i_add_term2[51], i_add_term2[52], i_add_term2[53], i_add_term2[54], i_add_term2[55], i_add_term2[56], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], sum[45], sum[46], sum[47], sum[48], sum[49], sum[50], sum[51], sum[52], sum[53], sum[54], sum[55], sum[56], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term1[45];
input i_add_term1[46];
input i_add_term1[47];
input i_add_term1[48];
input i_add_term1[49];
input i_add_term1[50];
input i_add_term1[51];
input i_add_term1[52];
input i_add_term1[53];
input i_add_term1[54];
input i_add_term1[55];
input i_add_term1[56];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
input i_add_term2[45];
input i_add_term2[46];
input i_add_term2[47];
input i_add_term2[48];
input i_add_term2[49];
input i_add_term2[50];
input i_add_term2[51];
input i_add_term2[52];
input i_add_term2[53];
input i_add_term2[54];
input i_add_term2[55];
input i_add_term2[56];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output sum[45];
output sum[46];
output sum[47];
output sum[48];
output sum[49];
output sum[50];
output sum[51];
output sum[52];
output sum[53];
output sum[54];
output sum[55];
output sum[56];
output cout;

NOR2X1 NOR2X1_1 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_269_) );
OAI21X1 OAI21X1_1 ( .A(_267_), .B(_269_), .C(_268_), .Y(_17__1_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_263_) );
NAND3X1 NAND3X1_1 ( .A(_267_), .B(_268_), .C(_263_), .Y(_264_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_265_) );
OAI21X1 OAI21X1_2 ( .A(_269_), .B(_265_), .C(w_cout_5_), .Y(_266_) );
NAND2X1 NAND2X1_1 ( .A(_266_), .B(_264_), .Y(_0__20_) );
INVX1 INVX1_1 ( .A(_17__3_), .Y(_274_) );
NAND2X1 NAND2X1_2 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_275_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_276_) );
OAI21X1 OAI21X1_3 ( .A(_274_), .B(_276_), .C(_275_), .Y(_16_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_270_) );
NAND3X1 NAND3X1_2 ( .A(_274_), .B(_275_), .C(_270_), .Y(_271_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_272_) );
OAI21X1 OAI21X1_4 ( .A(_276_), .B(_272_), .C(_17__3_), .Y(_273_) );
NAND2X1 NAND2X1_3 ( .A(_273_), .B(_271_), .Y(_0__23_) );
INVX1 INVX1_2 ( .A(_17__1_), .Y(_281_) );
NAND2X1 NAND2X1_4 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_282_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_283_) );
OAI21X1 OAI21X1_5 ( .A(_281_), .B(_283_), .C(_282_), .Y(_17__2_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_277_) );
NAND3X1 NAND3X1_3 ( .A(_281_), .B(_282_), .C(_277_), .Y(_278_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_279_) );
OAI21X1 OAI21X1_6 ( .A(_283_), .B(_279_), .C(_17__1_), .Y(_280_) );
NAND2X1 NAND2X1_5 ( .A(_280_), .B(_278_), .Y(_0__21_) );
INVX1 INVX1_3 ( .A(_17__2_), .Y(_288_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_289_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_290_) );
OAI21X1 OAI21X1_7 ( .A(_288_), .B(_290_), .C(_289_), .Y(_17__3_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_284_) );
NAND3X1 NAND3X1_4 ( .A(_288_), .B(_289_), .C(_284_), .Y(_285_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_286_) );
OAI21X1 OAI21X1_8 ( .A(_290_), .B(_286_), .C(_17__2_), .Y(_287_) );
NAND2X1 NAND2X1_7 ( .A(_287_), .B(_285_), .Y(_0__22_) );
INVX1 INVX1_4 ( .A(i_add_term1[20]), .Y(_291_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[20]), .B(_291_), .Y(_292_) );
INVX1 INVX1_5 ( .A(i_add_term2[20]), .Y(_293_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term1[20]), .B(_293_), .Y(_294_) );
INVX1 INVX1_6 ( .A(i_add_term1[21]), .Y(_295_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[21]), .B(_295_), .Y(_296_) );
INVX1 INVX1_7 ( .A(i_add_term2[21]), .Y(_297_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term1[21]), .B(_297_), .Y(_298_) );
OAI22X1 OAI22X1_1 ( .A(_292_), .B(_294_), .C(_296_), .D(_298_), .Y(_299_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_300_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_301_) );
NOR2X1 NOR2X1_10 ( .A(_300_), .B(_301_), .Y(_302_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_303_) );
NAND2X1 NAND2X1_8 ( .A(_302_), .B(_303_), .Y(_304_) );
NOR2X1 NOR2X1_11 ( .A(_299_), .B(_304_), .Y(_18_) );
INVX1 INVX1_8 ( .A(_16_), .Y(_305_) );
NAND2X1 NAND2X1_9 ( .A(1'b0), .B(_18_), .Y(_306_) );
OAI21X1 OAI21X1_9 ( .A(_18_), .B(_305_), .C(_306_), .Y(w_cout_6_) );
INVX1 INVX1_9 ( .A(w_cout_6_), .Y(_311_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_312_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_313_) );
OAI21X1 OAI21X1_10 ( .A(_311_), .B(_313_), .C(_312_), .Y(_20__1_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_307_) );
NAND3X1 NAND3X1_5 ( .A(_311_), .B(_312_), .C(_307_), .Y(_308_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_309_) );
OAI21X1 OAI21X1_11 ( .A(_313_), .B(_309_), .C(w_cout_6_), .Y(_310_) );
NAND2X1 NAND2X1_11 ( .A(_310_), .B(_308_), .Y(_0__24_) );
INVX1 INVX1_10 ( .A(_20__3_), .Y(_318_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_319_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_320_) );
OAI21X1 OAI21X1_12 ( .A(_318_), .B(_320_), .C(_319_), .Y(_19_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_314_) );
NAND3X1 NAND3X1_6 ( .A(_318_), .B(_319_), .C(_314_), .Y(_315_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_316_) );
OAI21X1 OAI21X1_13 ( .A(_320_), .B(_316_), .C(_20__3_), .Y(_317_) );
NAND2X1 NAND2X1_13 ( .A(_317_), .B(_315_), .Y(_0__27_) );
INVX1 INVX1_11 ( .A(_20__1_), .Y(_325_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_326_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_327_) );
OAI21X1 OAI21X1_14 ( .A(_325_), .B(_327_), .C(_326_), .Y(_20__2_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_321_) );
NAND3X1 NAND3X1_7 ( .A(_325_), .B(_326_), .C(_321_), .Y(_322_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_323_) );
OAI21X1 OAI21X1_15 ( .A(_327_), .B(_323_), .C(_20__1_), .Y(_324_) );
NAND2X1 NAND2X1_15 ( .A(_324_), .B(_322_), .Y(_0__25_) );
INVX1 INVX1_12 ( .A(_20__2_), .Y(_332_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_333_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_334_) );
OAI21X1 OAI21X1_16 ( .A(_332_), .B(_334_), .C(_333_), .Y(_20__3_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_328_) );
NAND3X1 NAND3X1_8 ( .A(_332_), .B(_333_), .C(_328_), .Y(_329_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_330_) );
OAI21X1 OAI21X1_17 ( .A(_334_), .B(_330_), .C(_20__2_), .Y(_331_) );
NAND2X1 NAND2X1_17 ( .A(_331_), .B(_329_), .Y(_0__26_) );
INVX1 INVX1_13 ( .A(i_add_term1[24]), .Y(_335_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[24]), .B(_335_), .Y(_336_) );
INVX1 INVX1_14 ( .A(i_add_term2[24]), .Y(_337_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term1[24]), .B(_337_), .Y(_338_) );
INVX1 INVX1_15 ( .A(i_add_term1[25]), .Y(_339_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[25]), .B(_339_), .Y(_340_) );
INVX1 INVX1_16 ( .A(i_add_term2[25]), .Y(_341_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term1[25]), .B(_341_), .Y(_342_) );
OAI22X1 OAI22X1_2 ( .A(_336_), .B(_338_), .C(_340_), .D(_342_), .Y(_343_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_344_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_345_) );
NOR2X1 NOR2X1_21 ( .A(_344_), .B(_345_), .Y(_346_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_347_) );
NAND2X1 NAND2X1_18 ( .A(_346_), .B(_347_), .Y(_348_) );
NOR2X1 NOR2X1_22 ( .A(_343_), .B(_348_), .Y(_21_) );
INVX1 INVX1_17 ( .A(_19_), .Y(_349_) );
NAND2X1 NAND2X1_19 ( .A(1'b0), .B(_21_), .Y(_350_) );
OAI21X1 OAI21X1_18 ( .A(_21_), .B(_349_), .C(_350_), .Y(w_cout_7_) );
INVX1 INVX1_18 ( .A(w_cout_7_), .Y(_355_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_356_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_357_) );
OAI21X1 OAI21X1_19 ( .A(_355_), .B(_357_), .C(_356_), .Y(_23__1_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_351_) );
NAND3X1 NAND3X1_9 ( .A(_355_), .B(_356_), .C(_351_), .Y(_352_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_353_) );
OAI21X1 OAI21X1_20 ( .A(_357_), .B(_353_), .C(w_cout_7_), .Y(_354_) );
NAND2X1 NAND2X1_21 ( .A(_354_), .B(_352_), .Y(_0__28_) );
INVX1 INVX1_19 ( .A(_23__3_), .Y(_362_) );
NAND2X1 NAND2X1_22 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_363_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_364_) );
OAI21X1 OAI21X1_21 ( .A(_362_), .B(_364_), .C(_363_), .Y(_22_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_358_) );
NAND3X1 NAND3X1_10 ( .A(_362_), .B(_363_), .C(_358_), .Y(_359_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_360_) );
OAI21X1 OAI21X1_22 ( .A(_364_), .B(_360_), .C(_23__3_), .Y(_361_) );
NAND2X1 NAND2X1_23 ( .A(_361_), .B(_359_), .Y(_0__31_) );
INVX1 INVX1_20 ( .A(_23__1_), .Y(_369_) );
NAND2X1 NAND2X1_24 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_370_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_371_) );
OAI21X1 OAI21X1_23 ( .A(_369_), .B(_371_), .C(_370_), .Y(_23__2_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_365_) );
NAND3X1 NAND3X1_11 ( .A(_369_), .B(_370_), .C(_365_), .Y(_366_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_367_) );
OAI21X1 OAI21X1_24 ( .A(_371_), .B(_367_), .C(_23__1_), .Y(_368_) );
NAND2X1 NAND2X1_25 ( .A(_368_), .B(_366_), .Y(_0__29_) );
INVX1 INVX1_21 ( .A(_23__2_), .Y(_376_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_377_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_378_) );
OAI21X1 OAI21X1_25 ( .A(_376_), .B(_378_), .C(_377_), .Y(_23__3_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_372_) );
NAND3X1 NAND3X1_12 ( .A(_376_), .B(_377_), .C(_372_), .Y(_373_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_374_) );
OAI21X1 OAI21X1_26 ( .A(_378_), .B(_374_), .C(_23__2_), .Y(_375_) );
NAND2X1 NAND2X1_27 ( .A(_375_), .B(_373_), .Y(_0__30_) );
INVX1 INVX1_22 ( .A(i_add_term1[28]), .Y(_379_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[28]), .B(_379_), .Y(_380_) );
INVX1 INVX1_23 ( .A(i_add_term2[28]), .Y(_381_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term1[28]), .B(_381_), .Y(_382_) );
INVX1 INVX1_24 ( .A(i_add_term1[29]), .Y(_383_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[29]), .B(_383_), .Y(_384_) );
INVX1 INVX1_25 ( .A(i_add_term2[29]), .Y(_385_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term1[29]), .B(_385_), .Y(_386_) );
OAI22X1 OAI22X1_3 ( .A(_380_), .B(_382_), .C(_384_), .D(_386_), .Y(_387_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_388_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_389_) );
NOR2X1 NOR2X1_32 ( .A(_388_), .B(_389_), .Y(_390_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_391_) );
NAND2X1 NAND2X1_28 ( .A(_390_), .B(_391_), .Y(_392_) );
NOR2X1 NOR2X1_33 ( .A(_387_), .B(_392_), .Y(_24_) );
INVX1 INVX1_26 ( .A(_22_), .Y(_393_) );
NAND2X1 NAND2X1_29 ( .A(1'b0), .B(_24_), .Y(_394_) );
OAI21X1 OAI21X1_27 ( .A(_24_), .B(_393_), .C(_394_), .Y(w_cout_8_) );
INVX1 INVX1_27 ( .A(w_cout_8_), .Y(_399_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_400_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_401_) );
OAI21X1 OAI21X1_28 ( .A(_399_), .B(_401_), .C(_400_), .Y(_26__1_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_395_) );
NAND3X1 NAND3X1_13 ( .A(_399_), .B(_400_), .C(_395_), .Y(_396_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_397_) );
OAI21X1 OAI21X1_29 ( .A(_401_), .B(_397_), .C(w_cout_8_), .Y(_398_) );
NAND2X1 NAND2X1_31 ( .A(_398_), .B(_396_), .Y(_0__32_) );
INVX1 INVX1_28 ( .A(_26__3_), .Y(_406_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_407_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_408_) );
OAI21X1 OAI21X1_30 ( .A(_406_), .B(_408_), .C(_407_), .Y(_25_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_402_) );
NAND3X1 NAND3X1_14 ( .A(_406_), .B(_407_), .C(_402_), .Y(_403_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_404_) );
OAI21X1 OAI21X1_31 ( .A(_408_), .B(_404_), .C(_26__3_), .Y(_405_) );
NAND2X1 NAND2X1_33 ( .A(_405_), .B(_403_), .Y(_0__35_) );
INVX1 INVX1_29 ( .A(_26__1_), .Y(_413_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_414_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_415_) );
OAI21X1 OAI21X1_32 ( .A(_413_), .B(_415_), .C(_414_), .Y(_26__2_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_409_) );
NAND3X1 NAND3X1_15 ( .A(_413_), .B(_414_), .C(_409_), .Y(_410_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_411_) );
OAI21X1 OAI21X1_33 ( .A(_415_), .B(_411_), .C(_26__1_), .Y(_412_) );
NAND2X1 NAND2X1_35 ( .A(_412_), .B(_410_), .Y(_0__33_) );
INVX1 INVX1_30 ( .A(_26__2_), .Y(_420_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_421_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_422_) );
OAI21X1 OAI21X1_34 ( .A(_420_), .B(_422_), .C(_421_), .Y(_26__3_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_416_) );
NAND3X1 NAND3X1_16 ( .A(_420_), .B(_421_), .C(_416_), .Y(_417_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_418_) );
OAI21X1 OAI21X1_35 ( .A(_422_), .B(_418_), .C(_26__2_), .Y(_419_) );
NAND2X1 NAND2X1_37 ( .A(_419_), .B(_417_), .Y(_0__34_) );
INVX1 INVX1_31 ( .A(i_add_term1[32]), .Y(_423_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[32]), .B(_423_), .Y(_424_) );
INVX1 INVX1_32 ( .A(i_add_term2[32]), .Y(_425_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term1[32]), .B(_425_), .Y(_426_) );
INVX1 INVX1_33 ( .A(i_add_term1[33]), .Y(_427_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[33]), .B(_427_), .Y(_428_) );
INVX1 INVX1_34 ( .A(i_add_term2[33]), .Y(_429_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term1[33]), .B(_429_), .Y(_430_) );
OAI22X1 OAI22X1_4 ( .A(_424_), .B(_426_), .C(_428_), .D(_430_), .Y(_431_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_432_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_433_) );
NOR2X1 NOR2X1_43 ( .A(_432_), .B(_433_), .Y(_434_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_435_) );
NAND2X1 NAND2X1_38 ( .A(_434_), .B(_435_), .Y(_436_) );
NOR2X1 NOR2X1_44 ( .A(_431_), .B(_436_), .Y(_27_) );
INVX1 INVX1_35 ( .A(_25_), .Y(_437_) );
NAND2X1 NAND2X1_39 ( .A(1'b0), .B(_27_), .Y(_438_) );
OAI21X1 OAI21X1_36 ( .A(_27_), .B(_437_), .C(_438_), .Y(w_cout_9_) );
INVX1 INVX1_36 ( .A(w_cout_9_), .Y(_443_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_444_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_445_) );
OAI21X1 OAI21X1_37 ( .A(_443_), .B(_445_), .C(_444_), .Y(_29__1_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_439_) );
NAND3X1 NAND3X1_17 ( .A(_443_), .B(_444_), .C(_439_), .Y(_440_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_441_) );
OAI21X1 OAI21X1_38 ( .A(_445_), .B(_441_), .C(w_cout_9_), .Y(_442_) );
NAND2X1 NAND2X1_41 ( .A(_442_), .B(_440_), .Y(_0__36_) );
INVX1 INVX1_37 ( .A(_29__3_), .Y(_450_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_451_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_452_) );
OAI21X1 OAI21X1_39 ( .A(_450_), .B(_452_), .C(_451_), .Y(_28_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_446_) );
NAND3X1 NAND3X1_18 ( .A(_450_), .B(_451_), .C(_446_), .Y(_447_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_448_) );
OAI21X1 OAI21X1_40 ( .A(_452_), .B(_448_), .C(_29__3_), .Y(_449_) );
NAND2X1 NAND2X1_43 ( .A(_449_), .B(_447_), .Y(_0__39_) );
INVX1 INVX1_38 ( .A(_29__1_), .Y(_457_) );
NAND2X1 NAND2X1_44 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_458_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_459_) );
OAI21X1 OAI21X1_41 ( .A(_457_), .B(_459_), .C(_458_), .Y(_29__2_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_453_) );
NAND3X1 NAND3X1_19 ( .A(_457_), .B(_458_), .C(_453_), .Y(_454_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_455_) );
OAI21X1 OAI21X1_42 ( .A(_459_), .B(_455_), .C(_29__1_), .Y(_456_) );
NAND2X1 NAND2X1_45 ( .A(_456_), .B(_454_), .Y(_0__37_) );
INVX1 INVX1_39 ( .A(_29__2_), .Y(_464_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_465_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_466_) );
OAI21X1 OAI21X1_43 ( .A(_464_), .B(_466_), .C(_465_), .Y(_29__3_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_460_) );
NAND3X1 NAND3X1_20 ( .A(_464_), .B(_465_), .C(_460_), .Y(_461_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_462_) );
OAI21X1 OAI21X1_44 ( .A(_466_), .B(_462_), .C(_29__2_), .Y(_463_) );
NAND2X1 NAND2X1_47 ( .A(_463_), .B(_461_), .Y(_0__38_) );
INVX1 INVX1_40 ( .A(i_add_term1[36]), .Y(_467_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[36]), .B(_467_), .Y(_468_) );
INVX1 INVX1_41 ( .A(i_add_term2[36]), .Y(_469_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term1[36]), .B(_469_), .Y(_470_) );
INVX1 INVX1_42 ( .A(i_add_term1[37]), .Y(_471_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[37]), .B(_471_), .Y(_472_) );
INVX1 INVX1_43 ( .A(i_add_term2[37]), .Y(_473_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term1[37]), .B(_473_), .Y(_474_) );
OAI22X1 OAI22X1_5 ( .A(_468_), .B(_470_), .C(_472_), .D(_474_), .Y(_475_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_476_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_477_) );
NOR2X1 NOR2X1_54 ( .A(_476_), .B(_477_), .Y(_478_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_479_) );
NAND2X1 NAND2X1_48 ( .A(_478_), .B(_479_), .Y(_480_) );
NOR2X1 NOR2X1_55 ( .A(_475_), .B(_480_), .Y(_30_) );
INVX1 INVX1_44 ( .A(_28_), .Y(_481_) );
NAND2X1 NAND2X1_49 ( .A(1'b0), .B(_30_), .Y(_482_) );
OAI21X1 OAI21X1_45 ( .A(_30_), .B(_481_), .C(_482_), .Y(w_cout_10_) );
INVX1 INVX1_45 ( .A(w_cout_10_), .Y(_487_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_488_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_489_) );
OAI21X1 OAI21X1_46 ( .A(_487_), .B(_489_), .C(_488_), .Y(_32__1_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_483_) );
NAND3X1 NAND3X1_21 ( .A(_487_), .B(_488_), .C(_483_), .Y(_484_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_485_) );
OAI21X1 OAI21X1_47 ( .A(_489_), .B(_485_), .C(w_cout_10_), .Y(_486_) );
NAND2X1 NAND2X1_51 ( .A(_486_), .B(_484_), .Y(_0__40_) );
INVX1 INVX1_46 ( .A(_32__3_), .Y(_494_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_495_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_496_) );
OAI21X1 OAI21X1_48 ( .A(_494_), .B(_496_), .C(_495_), .Y(_31_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_490_) );
NAND3X1 NAND3X1_22 ( .A(_494_), .B(_495_), .C(_490_), .Y(_491_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_492_) );
OAI21X1 OAI21X1_49 ( .A(_496_), .B(_492_), .C(_32__3_), .Y(_493_) );
NAND2X1 NAND2X1_53 ( .A(_493_), .B(_491_), .Y(_0__43_) );
INVX1 INVX1_47 ( .A(_32__1_), .Y(_501_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_502_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_503_) );
OAI21X1 OAI21X1_50 ( .A(_501_), .B(_503_), .C(_502_), .Y(_32__2_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_497_) );
NAND3X1 NAND3X1_23 ( .A(_501_), .B(_502_), .C(_497_), .Y(_498_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_499_) );
OAI21X1 OAI21X1_51 ( .A(_503_), .B(_499_), .C(_32__1_), .Y(_500_) );
NAND2X1 NAND2X1_55 ( .A(_500_), .B(_498_), .Y(_0__41_) );
INVX1 INVX1_48 ( .A(_32__2_), .Y(_508_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_509_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_510_) );
OAI21X1 OAI21X1_52 ( .A(_508_), .B(_510_), .C(_509_), .Y(_32__3_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_504_) );
NAND3X1 NAND3X1_24 ( .A(_508_), .B(_509_), .C(_504_), .Y(_505_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_506_) );
OAI21X1 OAI21X1_53 ( .A(_510_), .B(_506_), .C(_32__2_), .Y(_507_) );
NAND2X1 NAND2X1_57 ( .A(_507_), .B(_505_), .Y(_0__42_) );
INVX1 INVX1_49 ( .A(i_add_term1[40]), .Y(_511_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[40]), .B(_511_), .Y(_512_) );
INVX1 INVX1_50 ( .A(i_add_term2[40]), .Y(_513_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term1[40]), .B(_513_), .Y(_514_) );
INVX1 INVX1_51 ( .A(i_add_term1[41]), .Y(_515_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[41]), .B(_515_), .Y(_516_) );
INVX1 INVX1_52 ( .A(i_add_term2[41]), .Y(_517_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term1[41]), .B(_517_), .Y(_518_) );
OAI22X1 OAI22X1_6 ( .A(_512_), .B(_514_), .C(_516_), .D(_518_), .Y(_519_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_520_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_521_) );
NOR2X1 NOR2X1_65 ( .A(_520_), .B(_521_), .Y(_522_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_523_) );
NAND2X1 NAND2X1_58 ( .A(_522_), .B(_523_), .Y(_524_) );
NOR2X1 NOR2X1_66 ( .A(_519_), .B(_524_), .Y(_33_) );
INVX1 INVX1_53 ( .A(_31_), .Y(_525_) );
NAND2X1 NAND2X1_59 ( .A(1'b0), .B(_33_), .Y(_526_) );
OAI21X1 OAI21X1_54 ( .A(_33_), .B(_525_), .C(_526_), .Y(w_cout_11_) );
INVX1 INVX1_54 ( .A(w_cout_11_), .Y(_531_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_532_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_533_) );
OAI21X1 OAI21X1_55 ( .A(_531_), .B(_533_), .C(_532_), .Y(_35__1_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_527_) );
NAND3X1 NAND3X1_25 ( .A(_531_), .B(_532_), .C(_527_), .Y(_528_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_529_) );
OAI21X1 OAI21X1_56 ( .A(_533_), .B(_529_), .C(w_cout_11_), .Y(_530_) );
NAND2X1 NAND2X1_61 ( .A(_530_), .B(_528_), .Y(_0__44_) );
INVX1 INVX1_55 ( .A(_35__3_), .Y(_538_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_539_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_540_) );
OAI21X1 OAI21X1_57 ( .A(_538_), .B(_540_), .C(_539_), .Y(_34_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_534_) );
NAND3X1 NAND3X1_26 ( .A(_538_), .B(_539_), .C(_534_), .Y(_535_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_536_) );
OAI21X1 OAI21X1_58 ( .A(_540_), .B(_536_), .C(_35__3_), .Y(_537_) );
NAND2X1 NAND2X1_63 ( .A(_537_), .B(_535_), .Y(_0__47_) );
INVX1 INVX1_56 ( .A(_35__1_), .Y(_545_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_546_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_547_) );
OAI21X1 OAI21X1_59 ( .A(_545_), .B(_547_), .C(_546_), .Y(_35__2_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_541_) );
NAND3X1 NAND3X1_27 ( .A(_545_), .B(_546_), .C(_541_), .Y(_542_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_543_) );
OAI21X1 OAI21X1_60 ( .A(_547_), .B(_543_), .C(_35__1_), .Y(_544_) );
NAND2X1 NAND2X1_65 ( .A(_544_), .B(_542_), .Y(_0__45_) );
INVX1 INVX1_57 ( .A(_35__2_), .Y(_552_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_553_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_554_) );
OAI21X1 OAI21X1_61 ( .A(_552_), .B(_554_), .C(_553_), .Y(_35__3_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_548_) );
NAND3X1 NAND3X1_28 ( .A(_552_), .B(_553_), .C(_548_), .Y(_549_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_550_) );
OAI21X1 OAI21X1_62 ( .A(_554_), .B(_550_), .C(_35__2_), .Y(_551_) );
NAND2X1 NAND2X1_67 ( .A(_551_), .B(_549_), .Y(_0__46_) );
INVX1 INVX1_58 ( .A(i_add_term1[44]), .Y(_555_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[44]), .B(_555_), .Y(_556_) );
INVX1 INVX1_59 ( .A(i_add_term2[44]), .Y(_557_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term1[44]), .B(_557_), .Y(_558_) );
INVX1 INVX1_60 ( .A(i_add_term1[45]), .Y(_559_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[45]), .B(_559_), .Y(_560_) );
INVX1 INVX1_61 ( .A(i_add_term2[45]), .Y(_561_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term1[45]), .B(_561_), .Y(_562_) );
OAI22X1 OAI22X1_7 ( .A(_556_), .B(_558_), .C(_560_), .D(_562_), .Y(_563_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_564_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_565_) );
NOR2X1 NOR2X1_76 ( .A(_564_), .B(_565_), .Y(_566_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_567_) );
NAND2X1 NAND2X1_68 ( .A(_566_), .B(_567_), .Y(_568_) );
NOR2X1 NOR2X1_77 ( .A(_563_), .B(_568_), .Y(_36_) );
INVX1 INVX1_62 ( .A(_34_), .Y(_569_) );
NAND2X1 NAND2X1_69 ( .A(1'b0), .B(_36_), .Y(_570_) );
OAI21X1 OAI21X1_63 ( .A(_36_), .B(_569_), .C(_570_), .Y(w_cout_12_) );
INVX1 INVX1_63 ( .A(w_cout_12_), .Y(_575_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_576_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_577_) );
OAI21X1 OAI21X1_64 ( .A(_575_), .B(_577_), .C(_576_), .Y(_38__1_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_571_) );
NAND3X1 NAND3X1_29 ( .A(_575_), .B(_576_), .C(_571_), .Y(_572_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_573_) );
OAI21X1 OAI21X1_65 ( .A(_577_), .B(_573_), .C(w_cout_12_), .Y(_574_) );
NAND2X1 NAND2X1_71 ( .A(_574_), .B(_572_), .Y(_0__48_) );
INVX1 INVX1_64 ( .A(_38__3_), .Y(_582_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_583_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_584_) );
OAI21X1 OAI21X1_66 ( .A(_582_), .B(_584_), .C(_583_), .Y(_37_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_578_) );
NAND3X1 NAND3X1_30 ( .A(_582_), .B(_583_), .C(_578_), .Y(_579_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_580_) );
OAI21X1 OAI21X1_67 ( .A(_584_), .B(_580_), .C(_38__3_), .Y(_581_) );
NAND2X1 NAND2X1_73 ( .A(_581_), .B(_579_), .Y(_0__51_) );
INVX1 INVX1_65 ( .A(_38__1_), .Y(_589_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_590_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_591_) );
OAI21X1 OAI21X1_68 ( .A(_589_), .B(_591_), .C(_590_), .Y(_38__2_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_585_) );
NAND3X1 NAND3X1_31 ( .A(_589_), .B(_590_), .C(_585_), .Y(_586_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_587_) );
OAI21X1 OAI21X1_69 ( .A(_591_), .B(_587_), .C(_38__1_), .Y(_588_) );
NAND2X1 NAND2X1_75 ( .A(_588_), .B(_586_), .Y(_0__49_) );
INVX1 INVX1_66 ( .A(_38__2_), .Y(_596_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_597_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_598_) );
OAI21X1 OAI21X1_70 ( .A(_596_), .B(_598_), .C(_597_), .Y(_38__3_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_592_) );
NAND3X1 NAND3X1_32 ( .A(_596_), .B(_597_), .C(_592_), .Y(_593_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_594_) );
OAI21X1 OAI21X1_71 ( .A(_598_), .B(_594_), .C(_38__2_), .Y(_595_) );
NAND2X1 NAND2X1_77 ( .A(_595_), .B(_593_), .Y(_0__50_) );
INVX1 INVX1_67 ( .A(i_add_term1[48]), .Y(_599_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[48]), .B(_599_), .Y(_600_) );
INVX1 INVX1_68 ( .A(i_add_term2[48]), .Y(_601_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term1[48]), .B(_601_), .Y(_602_) );
INVX1 INVX1_69 ( .A(i_add_term1[49]), .Y(_603_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[49]), .B(_603_), .Y(_604_) );
INVX1 INVX1_70 ( .A(i_add_term2[49]), .Y(_605_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term1[49]), .B(_605_), .Y(_606_) );
OAI22X1 OAI22X1_8 ( .A(_600_), .B(_602_), .C(_604_), .D(_606_), .Y(_607_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_608_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_609_) );
NOR2X1 NOR2X1_87 ( .A(_608_), .B(_609_), .Y(_610_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_611_) );
NAND2X1 NAND2X1_78 ( .A(_610_), .B(_611_), .Y(_612_) );
NOR2X1 NOR2X1_88 ( .A(_607_), .B(_612_), .Y(_39_) );
INVX1 INVX1_71 ( .A(_37_), .Y(_613_) );
NAND2X1 NAND2X1_79 ( .A(1'b0), .B(_39_), .Y(_614_) );
OAI21X1 OAI21X1_72 ( .A(_39_), .B(_613_), .C(_614_), .Y(w_cout_13_) );
INVX1 INVX1_72 ( .A(w_cout_13_), .Y(_619_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_620_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_621_) );
OAI21X1 OAI21X1_73 ( .A(_619_), .B(_621_), .C(_620_), .Y(_41__1_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_615_) );
NAND3X1 NAND3X1_33 ( .A(_619_), .B(_620_), .C(_615_), .Y(_616_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_617_) );
OAI21X1 OAI21X1_74 ( .A(_621_), .B(_617_), .C(w_cout_13_), .Y(_618_) );
NAND2X1 NAND2X1_81 ( .A(_618_), .B(_616_), .Y(_0__52_) );
INVX1 INVX1_73 ( .A(_41__3_), .Y(_626_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_627_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_628_) );
OAI21X1 OAI21X1_75 ( .A(_626_), .B(_628_), .C(_627_), .Y(_40_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_622_) );
NAND3X1 NAND3X1_34 ( .A(_626_), .B(_627_), .C(_622_), .Y(_623_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_624_) );
OAI21X1 OAI21X1_76 ( .A(_628_), .B(_624_), .C(_41__3_), .Y(_625_) );
NAND2X1 NAND2X1_83 ( .A(_625_), .B(_623_), .Y(_0__55_) );
INVX1 INVX1_74 ( .A(_41__1_), .Y(_633_) );
NAND2X1 NAND2X1_84 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_634_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_635_) );
OAI21X1 OAI21X1_77 ( .A(_633_), .B(_635_), .C(_634_), .Y(_41__2_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_629_) );
NAND3X1 NAND3X1_35 ( .A(_633_), .B(_634_), .C(_629_), .Y(_630_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_631_) );
OAI21X1 OAI21X1_78 ( .A(_635_), .B(_631_), .C(_41__1_), .Y(_632_) );
NAND2X1 NAND2X1_85 ( .A(_632_), .B(_630_), .Y(_0__53_) );
INVX1 INVX1_75 ( .A(_41__2_), .Y(_640_) );
NAND2X1 NAND2X1_86 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_641_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_642_) );
OAI21X1 OAI21X1_79 ( .A(_640_), .B(_642_), .C(_641_), .Y(_41__3_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_636_) );
NAND3X1 NAND3X1_36 ( .A(_640_), .B(_641_), .C(_636_), .Y(_637_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_638_) );
OAI21X1 OAI21X1_80 ( .A(_642_), .B(_638_), .C(_41__2_), .Y(_639_) );
NAND2X1 NAND2X1_87 ( .A(_639_), .B(_637_), .Y(_0__54_) );
INVX1 INVX1_76 ( .A(i_add_term1[52]), .Y(_643_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[52]), .B(_643_), .Y(_644_) );
INVX1 INVX1_77 ( .A(i_add_term2[52]), .Y(_645_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term1[52]), .B(_645_), .Y(_646_) );
INVX1 INVX1_78 ( .A(i_add_term1[53]), .Y(_647_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[53]), .B(_647_), .Y(_648_) );
INVX1 INVX1_79 ( .A(i_add_term2[53]), .Y(_649_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term1[53]), .B(_649_), .Y(_650_) );
OAI22X1 OAI22X1_9 ( .A(_644_), .B(_646_), .C(_648_), .D(_650_), .Y(_651_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_652_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_653_) );
NOR2X1 NOR2X1_98 ( .A(_652_), .B(_653_), .Y(_654_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_655_) );
NAND2X1 NAND2X1_88 ( .A(_654_), .B(_655_), .Y(_656_) );
NOR2X1 NOR2X1_99 ( .A(_651_), .B(_656_), .Y(_42_) );
INVX1 INVX1_80 ( .A(_40_), .Y(_657_) );
NAND2X1 NAND2X1_89 ( .A(1'b0), .B(_42_), .Y(_658_) );
OAI21X1 OAI21X1_81 ( .A(_42_), .B(_657_), .C(_658_), .Y(cskip1_inst_cin) );
INVX1 INVX1_81 ( .A(cskip1_inst_cin), .Y(_663_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_664_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_665_) );
OAI21X1 OAI21X1_82 ( .A(_663_), .B(_665_), .C(_664_), .Y(cskip1_inst_cout0) );
OR2X2 OR2X2_37 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_659_) );
NAND3X1 NAND3X1_37 ( .A(_663_), .B(_664_), .C(_659_), .Y(_660_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_661_) );
OAI21X1 OAI21X1_83 ( .A(_665_), .B(_661_), .C(cskip1_inst_cin), .Y(_662_) );
NAND2X1 NAND2X1_91 ( .A(_662_), .B(_660_), .Y(cskip1_inst_rca0_fa0_o_sum) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_666_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_667_) );
NOR2X1 NOR2X1_102 ( .A(_666_), .B(_667_), .Y(cskip1_inst_skip0_P) );
INVX1 INVX1_82 ( .A(cskip1_inst_cout0), .Y(_668_) );
NAND2X1 NAND2X1_92 ( .A(1'b0), .B(cskip1_inst_skip0_P), .Y(_669_) );
OAI21X1 OAI21X1_84 ( .A(cskip1_inst_skip0_P), .B(_668_), .C(_669_), .Y(w_cout_15_) );
BUFX2 BUFX2_1 ( .A(w_cout_15_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .A(_0__54_), .Y(sum[54]) );
BUFX2 BUFX2_57 ( .A(_0__55_), .Y(sum[55]) );
BUFX2 BUFX2_58 ( .A(cskip1_inst_rca0_fa0_o_sum), .Y(sum[56]) );
INVX1 INVX1_83 ( .A(1'b0), .Y(_47_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_48_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_49_) );
OAI21X1 OAI21X1_85 ( .A(_47_), .B(_49_), .C(_48_), .Y(_2__1_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_43_) );
NAND3X1 NAND3X1_38 ( .A(_47_), .B(_48_), .C(_43_), .Y(_44_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_45_) );
OAI21X1 OAI21X1_86 ( .A(_49_), .B(_45_), .C(1'b0), .Y(_46_) );
NAND2X1 NAND2X1_94 ( .A(_46_), .B(_44_), .Y(_0__0_) );
INVX1 INVX1_84 ( .A(_2__3_), .Y(_54_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_55_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_56_) );
OAI21X1 OAI21X1_87 ( .A(_54_), .B(_56_), .C(_55_), .Y(_1_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_50_) );
NAND3X1 NAND3X1_39 ( .A(_54_), .B(_55_), .C(_50_), .Y(_51_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_52_) );
OAI21X1 OAI21X1_88 ( .A(_56_), .B(_52_), .C(_2__3_), .Y(_53_) );
NAND2X1 NAND2X1_96 ( .A(_53_), .B(_51_), .Y(_0__3_) );
INVX1 INVX1_85 ( .A(_2__1_), .Y(_61_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_62_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_63_) );
OAI21X1 OAI21X1_89 ( .A(_61_), .B(_63_), .C(_62_), .Y(_2__2_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_57_) );
NAND3X1 NAND3X1_40 ( .A(_61_), .B(_62_), .C(_57_), .Y(_58_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_59_) );
OAI21X1 OAI21X1_90 ( .A(_63_), .B(_59_), .C(_2__1_), .Y(_60_) );
NAND2X1 NAND2X1_98 ( .A(_60_), .B(_58_), .Y(_0__1_) );
INVX1 INVX1_86 ( .A(_2__2_), .Y(_68_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_69_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_70_) );
OAI21X1 OAI21X1_91 ( .A(_68_), .B(_70_), .C(_69_), .Y(_2__3_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_64_) );
NAND3X1 NAND3X1_41 ( .A(_68_), .B(_69_), .C(_64_), .Y(_65_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_66_) );
OAI21X1 OAI21X1_92 ( .A(_70_), .B(_66_), .C(_2__2_), .Y(_67_) );
NAND2X1 NAND2X1_100 ( .A(_67_), .B(_65_), .Y(_0__2_) );
INVX1 INVX1_87 ( .A(i_add_term1[0]), .Y(_71_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term2[0]), .B(_71_), .Y(_72_) );
INVX1 INVX1_88 ( .A(i_add_term2[0]), .Y(_73_) );
NOR2X1 NOR2X1_108 ( .A(i_add_term1[0]), .B(_73_), .Y(_74_) );
INVX1 INVX1_89 ( .A(i_add_term1[1]), .Y(_75_) );
NOR2X1 NOR2X1_109 ( .A(i_add_term2[1]), .B(_75_), .Y(_76_) );
INVX1 INVX1_90 ( .A(i_add_term2[1]), .Y(_77_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term1[1]), .B(_77_), .Y(_78_) );
OAI22X1 OAI22X1_10 ( .A(_72_), .B(_74_), .C(_76_), .D(_78_), .Y(_79_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_80_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_81_) );
NOR2X1 NOR2X1_112 ( .A(_80_), .B(_81_), .Y(_82_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_83_) );
NAND2X1 NAND2X1_101 ( .A(_82_), .B(_83_), .Y(_84_) );
NOR2X1 NOR2X1_113 ( .A(_79_), .B(_84_), .Y(_3_) );
INVX1 INVX1_91 ( .A(_1_), .Y(_85_) );
NAND2X1 NAND2X1_102 ( .A(1'b0), .B(_3_), .Y(_86_) );
OAI21X1 OAI21X1_93 ( .A(_3_), .B(_85_), .C(_86_), .Y(w_cout_1_) );
INVX1 INVX1_92 ( .A(w_cout_1_), .Y(_91_) );
NAND2X1 NAND2X1_103 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_92_) );
NOR2X1 NOR2X1_114 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_93_) );
OAI21X1 OAI21X1_94 ( .A(_91_), .B(_93_), .C(_92_), .Y(_5__1_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_87_) );
NAND3X1 NAND3X1_42 ( .A(_91_), .B(_92_), .C(_87_), .Y(_88_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_89_) );
OAI21X1 OAI21X1_95 ( .A(_93_), .B(_89_), .C(w_cout_1_), .Y(_90_) );
NAND2X1 NAND2X1_104 ( .A(_90_), .B(_88_), .Y(_0__4_) );
INVX1 INVX1_93 ( .A(_5__3_), .Y(_98_) );
NAND2X1 NAND2X1_105 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_99_) );
NOR2X1 NOR2X1_115 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_100_) );
OAI21X1 OAI21X1_96 ( .A(_98_), .B(_100_), .C(_99_), .Y(_4_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_94_) );
NAND3X1 NAND3X1_43 ( .A(_98_), .B(_99_), .C(_94_), .Y(_95_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_96_) );
OAI21X1 OAI21X1_97 ( .A(_100_), .B(_96_), .C(_5__3_), .Y(_97_) );
NAND2X1 NAND2X1_106 ( .A(_97_), .B(_95_), .Y(_0__7_) );
INVX1 INVX1_94 ( .A(_5__1_), .Y(_105_) );
NAND2X1 NAND2X1_107 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_106_) );
NOR2X1 NOR2X1_116 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_107_) );
OAI21X1 OAI21X1_98 ( .A(_105_), .B(_107_), .C(_106_), .Y(_5__2_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_101_) );
NAND3X1 NAND3X1_44 ( .A(_105_), .B(_106_), .C(_101_), .Y(_102_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_103_) );
OAI21X1 OAI21X1_99 ( .A(_107_), .B(_103_), .C(_5__1_), .Y(_104_) );
NAND2X1 NAND2X1_108 ( .A(_104_), .B(_102_), .Y(_0__5_) );
INVX1 INVX1_95 ( .A(_5__2_), .Y(_112_) );
NAND2X1 NAND2X1_109 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_113_) );
NOR2X1 NOR2X1_117 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_114_) );
OAI21X1 OAI21X1_100 ( .A(_112_), .B(_114_), .C(_113_), .Y(_5__3_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_108_) );
NAND3X1 NAND3X1_45 ( .A(_112_), .B(_113_), .C(_108_), .Y(_109_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_110_) );
OAI21X1 OAI21X1_101 ( .A(_114_), .B(_110_), .C(_5__2_), .Y(_111_) );
NAND2X1 NAND2X1_110 ( .A(_111_), .B(_109_), .Y(_0__6_) );
INVX1 INVX1_96 ( .A(i_add_term1[4]), .Y(_115_) );
NOR2X1 NOR2X1_118 ( .A(i_add_term2[4]), .B(_115_), .Y(_116_) );
INVX1 INVX1_97 ( .A(i_add_term2[4]), .Y(_117_) );
NOR2X1 NOR2X1_119 ( .A(i_add_term1[4]), .B(_117_), .Y(_118_) );
INVX1 INVX1_98 ( .A(i_add_term1[5]), .Y(_119_) );
NOR2X1 NOR2X1_120 ( .A(i_add_term2[5]), .B(_119_), .Y(_120_) );
INVX1 INVX1_99 ( .A(i_add_term2[5]), .Y(_121_) );
NOR2X1 NOR2X1_121 ( .A(i_add_term1[5]), .B(_121_), .Y(_122_) );
OAI22X1 OAI22X1_11 ( .A(_116_), .B(_118_), .C(_120_), .D(_122_), .Y(_123_) );
NOR2X1 NOR2X1_122 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_124_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_125_) );
NOR2X1 NOR2X1_123 ( .A(_124_), .B(_125_), .Y(_126_) );
XOR2X1 XOR2X1_11 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_127_) );
NAND2X1 NAND2X1_111 ( .A(_126_), .B(_127_), .Y(_128_) );
NOR2X1 NOR2X1_124 ( .A(_123_), .B(_128_), .Y(_6_) );
INVX1 INVX1_100 ( .A(_4_), .Y(_129_) );
NAND2X1 NAND2X1_112 ( .A(1'b0), .B(_6_), .Y(_130_) );
OAI21X1 OAI21X1_102 ( .A(_6_), .B(_129_), .C(_130_), .Y(w_cout_2_) );
INVX1 INVX1_101 ( .A(w_cout_2_), .Y(_135_) );
NAND2X1 NAND2X1_113 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_136_) );
NOR2X1 NOR2X1_125 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_137_) );
OAI21X1 OAI21X1_103 ( .A(_135_), .B(_137_), .C(_136_), .Y(_8__1_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_131_) );
NAND3X1 NAND3X1_46 ( .A(_135_), .B(_136_), .C(_131_), .Y(_132_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_133_) );
OAI21X1 OAI21X1_104 ( .A(_137_), .B(_133_), .C(w_cout_2_), .Y(_134_) );
NAND2X1 NAND2X1_114 ( .A(_134_), .B(_132_), .Y(_0__8_) );
INVX1 INVX1_102 ( .A(_8__3_), .Y(_142_) );
NAND2X1 NAND2X1_115 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_143_) );
NOR2X1 NOR2X1_126 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_144_) );
OAI21X1 OAI21X1_105 ( .A(_142_), .B(_144_), .C(_143_), .Y(_7_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_138_) );
NAND3X1 NAND3X1_47 ( .A(_142_), .B(_143_), .C(_138_), .Y(_139_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_140_) );
OAI21X1 OAI21X1_106 ( .A(_144_), .B(_140_), .C(_8__3_), .Y(_141_) );
NAND2X1 NAND2X1_116 ( .A(_141_), .B(_139_), .Y(_0__11_) );
INVX1 INVX1_103 ( .A(_8__1_), .Y(_149_) );
NAND2X1 NAND2X1_117 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_150_) );
NOR2X1 NOR2X1_127 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_151_) );
OAI21X1 OAI21X1_107 ( .A(_149_), .B(_151_), .C(_150_), .Y(_8__2_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_145_) );
NAND3X1 NAND3X1_48 ( .A(_149_), .B(_150_), .C(_145_), .Y(_146_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_147_) );
OAI21X1 OAI21X1_108 ( .A(_151_), .B(_147_), .C(_8__1_), .Y(_148_) );
NAND2X1 NAND2X1_118 ( .A(_148_), .B(_146_), .Y(_0__9_) );
INVX1 INVX1_104 ( .A(_8__2_), .Y(_156_) );
NAND2X1 NAND2X1_119 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_157_) );
NOR2X1 NOR2X1_128 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_158_) );
OAI21X1 OAI21X1_109 ( .A(_156_), .B(_158_), .C(_157_), .Y(_8__3_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_152_) );
NAND3X1 NAND3X1_49 ( .A(_156_), .B(_157_), .C(_152_), .Y(_153_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_154_) );
OAI21X1 OAI21X1_110 ( .A(_158_), .B(_154_), .C(_8__2_), .Y(_155_) );
NAND2X1 NAND2X1_120 ( .A(_155_), .B(_153_), .Y(_0__10_) );
INVX1 INVX1_105 ( .A(i_add_term1[8]), .Y(_159_) );
NOR2X1 NOR2X1_129 ( .A(i_add_term2[8]), .B(_159_), .Y(_160_) );
INVX1 INVX1_106 ( .A(i_add_term2[8]), .Y(_161_) );
NOR2X1 NOR2X1_130 ( .A(i_add_term1[8]), .B(_161_), .Y(_162_) );
INVX1 INVX1_107 ( .A(i_add_term1[9]), .Y(_163_) );
NOR2X1 NOR2X1_131 ( .A(i_add_term2[9]), .B(_163_), .Y(_164_) );
INVX1 INVX1_108 ( .A(i_add_term2[9]), .Y(_165_) );
NOR2X1 NOR2X1_132 ( .A(i_add_term1[9]), .B(_165_), .Y(_166_) );
OAI22X1 OAI22X1_12 ( .A(_160_), .B(_162_), .C(_164_), .D(_166_), .Y(_167_) );
NOR2X1 NOR2X1_133 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_168_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_169_) );
NOR2X1 NOR2X1_134 ( .A(_168_), .B(_169_), .Y(_170_) );
XOR2X1 XOR2X1_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_171_) );
NAND2X1 NAND2X1_121 ( .A(_170_), .B(_171_), .Y(_172_) );
NOR2X1 NOR2X1_135 ( .A(_167_), .B(_172_), .Y(_9_) );
INVX1 INVX1_109 ( .A(_7_), .Y(_173_) );
NAND2X1 NAND2X1_122 ( .A(1'b0), .B(_9_), .Y(_174_) );
OAI21X1 OAI21X1_111 ( .A(_9_), .B(_173_), .C(_174_), .Y(w_cout_3_) );
INVX1 INVX1_110 ( .A(w_cout_3_), .Y(_179_) );
NAND2X1 NAND2X1_123 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_180_) );
NOR2X1 NOR2X1_136 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_181_) );
OAI21X1 OAI21X1_112 ( .A(_179_), .B(_181_), .C(_180_), .Y(_11__1_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_175_) );
NAND3X1 NAND3X1_50 ( .A(_179_), .B(_180_), .C(_175_), .Y(_176_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_177_) );
OAI21X1 OAI21X1_113 ( .A(_181_), .B(_177_), .C(w_cout_3_), .Y(_178_) );
NAND2X1 NAND2X1_124 ( .A(_178_), .B(_176_), .Y(_0__12_) );
INVX1 INVX1_111 ( .A(_11__3_), .Y(_186_) );
NAND2X1 NAND2X1_125 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_187_) );
NOR2X1 NOR2X1_137 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_188_) );
OAI21X1 OAI21X1_114 ( .A(_186_), .B(_188_), .C(_187_), .Y(_10_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_182_) );
NAND3X1 NAND3X1_51 ( .A(_186_), .B(_187_), .C(_182_), .Y(_183_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_184_) );
OAI21X1 OAI21X1_115 ( .A(_188_), .B(_184_), .C(_11__3_), .Y(_185_) );
NAND2X1 NAND2X1_126 ( .A(_185_), .B(_183_), .Y(_0__15_) );
INVX1 INVX1_112 ( .A(_11__1_), .Y(_193_) );
NAND2X1 NAND2X1_127 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_194_) );
NOR2X1 NOR2X1_138 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_195_) );
OAI21X1 OAI21X1_116 ( .A(_193_), .B(_195_), .C(_194_), .Y(_11__2_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_189_) );
NAND3X1 NAND3X1_52 ( .A(_193_), .B(_194_), .C(_189_), .Y(_190_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_191_) );
OAI21X1 OAI21X1_117 ( .A(_195_), .B(_191_), .C(_11__1_), .Y(_192_) );
NAND2X1 NAND2X1_128 ( .A(_192_), .B(_190_), .Y(_0__13_) );
INVX1 INVX1_113 ( .A(_11__2_), .Y(_200_) );
NAND2X1 NAND2X1_129 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_201_) );
NOR2X1 NOR2X1_139 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_202_) );
OAI21X1 OAI21X1_118 ( .A(_200_), .B(_202_), .C(_201_), .Y(_11__3_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_196_) );
NAND3X1 NAND3X1_53 ( .A(_200_), .B(_201_), .C(_196_), .Y(_197_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_198_) );
OAI21X1 OAI21X1_119 ( .A(_202_), .B(_198_), .C(_11__2_), .Y(_199_) );
NAND2X1 NAND2X1_130 ( .A(_199_), .B(_197_), .Y(_0__14_) );
INVX1 INVX1_114 ( .A(i_add_term1[12]), .Y(_203_) );
NOR2X1 NOR2X1_140 ( .A(i_add_term2[12]), .B(_203_), .Y(_204_) );
INVX1 INVX1_115 ( .A(i_add_term2[12]), .Y(_205_) );
NOR2X1 NOR2X1_141 ( .A(i_add_term1[12]), .B(_205_), .Y(_206_) );
INVX1 INVX1_116 ( .A(i_add_term1[13]), .Y(_207_) );
NOR2X1 NOR2X1_142 ( .A(i_add_term2[13]), .B(_207_), .Y(_208_) );
INVX1 INVX1_117 ( .A(i_add_term2[13]), .Y(_209_) );
NOR2X1 NOR2X1_143 ( .A(i_add_term1[13]), .B(_209_), .Y(_210_) );
OAI22X1 OAI22X1_13 ( .A(_204_), .B(_206_), .C(_208_), .D(_210_), .Y(_211_) );
NOR2X1 NOR2X1_144 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_212_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_213_) );
NOR2X1 NOR2X1_145 ( .A(_212_), .B(_213_), .Y(_214_) );
XOR2X1 XOR2X1_13 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_215_) );
NAND2X1 NAND2X1_131 ( .A(_214_), .B(_215_), .Y(_216_) );
NOR2X1 NOR2X1_146 ( .A(_211_), .B(_216_), .Y(_12_) );
INVX1 INVX1_118 ( .A(_10_), .Y(_217_) );
NAND2X1 NAND2X1_132 ( .A(1'b0), .B(_12_), .Y(_218_) );
OAI21X1 OAI21X1_120 ( .A(_12_), .B(_217_), .C(_218_), .Y(w_cout_4_) );
INVX1 INVX1_119 ( .A(w_cout_4_), .Y(_223_) );
NAND2X1 NAND2X1_133 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_224_) );
NOR2X1 NOR2X1_147 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_225_) );
OAI21X1 OAI21X1_121 ( .A(_223_), .B(_225_), .C(_224_), .Y(_14__1_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_219_) );
NAND3X1 NAND3X1_54 ( .A(_223_), .B(_224_), .C(_219_), .Y(_220_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_221_) );
OAI21X1 OAI21X1_122 ( .A(_225_), .B(_221_), .C(w_cout_4_), .Y(_222_) );
NAND2X1 NAND2X1_134 ( .A(_222_), .B(_220_), .Y(_0__16_) );
INVX1 INVX1_120 ( .A(_14__3_), .Y(_230_) );
NAND2X1 NAND2X1_135 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_231_) );
NOR2X1 NOR2X1_148 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_232_) );
OAI21X1 OAI21X1_123 ( .A(_230_), .B(_232_), .C(_231_), .Y(_13_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_226_) );
NAND3X1 NAND3X1_55 ( .A(_230_), .B(_231_), .C(_226_), .Y(_227_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_228_) );
OAI21X1 OAI21X1_124 ( .A(_232_), .B(_228_), .C(_14__3_), .Y(_229_) );
NAND2X1 NAND2X1_136 ( .A(_229_), .B(_227_), .Y(_0__19_) );
INVX1 INVX1_121 ( .A(_14__1_), .Y(_237_) );
NAND2X1 NAND2X1_137 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_238_) );
NOR2X1 NOR2X1_149 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_239_) );
OAI21X1 OAI21X1_125 ( .A(_237_), .B(_239_), .C(_238_), .Y(_14__2_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_233_) );
NAND3X1 NAND3X1_56 ( .A(_237_), .B(_238_), .C(_233_), .Y(_234_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_235_) );
OAI21X1 OAI21X1_126 ( .A(_239_), .B(_235_), .C(_14__1_), .Y(_236_) );
NAND2X1 NAND2X1_138 ( .A(_236_), .B(_234_), .Y(_0__17_) );
INVX1 INVX1_122 ( .A(_14__2_), .Y(_244_) );
NAND2X1 NAND2X1_139 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_245_) );
NOR2X1 NOR2X1_150 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_246_) );
OAI21X1 OAI21X1_127 ( .A(_244_), .B(_246_), .C(_245_), .Y(_14__3_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_240_) );
NAND3X1 NAND3X1_57 ( .A(_244_), .B(_245_), .C(_240_), .Y(_241_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_242_) );
OAI21X1 OAI21X1_128 ( .A(_246_), .B(_242_), .C(_14__2_), .Y(_243_) );
NAND2X1 NAND2X1_140 ( .A(_243_), .B(_241_), .Y(_0__18_) );
INVX1 INVX1_123 ( .A(i_add_term1[16]), .Y(_247_) );
NOR2X1 NOR2X1_151 ( .A(i_add_term2[16]), .B(_247_), .Y(_248_) );
INVX1 INVX1_124 ( .A(i_add_term2[16]), .Y(_249_) );
NOR2X1 NOR2X1_152 ( .A(i_add_term1[16]), .B(_249_), .Y(_250_) );
INVX1 INVX1_125 ( .A(i_add_term1[17]), .Y(_251_) );
NOR2X1 NOR2X1_153 ( .A(i_add_term2[17]), .B(_251_), .Y(_252_) );
INVX1 INVX1_126 ( .A(i_add_term2[17]), .Y(_253_) );
NOR2X1 NOR2X1_154 ( .A(i_add_term1[17]), .B(_253_), .Y(_254_) );
OAI22X1 OAI22X1_14 ( .A(_248_), .B(_250_), .C(_252_), .D(_254_), .Y(_255_) );
NOR2X1 NOR2X1_155 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_256_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_257_) );
NOR2X1 NOR2X1_156 ( .A(_256_), .B(_257_), .Y(_258_) );
XOR2X1 XOR2X1_14 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_259_) );
NAND2X1 NAND2X1_141 ( .A(_258_), .B(_259_), .Y(_260_) );
NOR2X1 NOR2X1_157 ( .A(_255_), .B(_260_), .Y(_15_) );
INVX1 INVX1_127 ( .A(_13_), .Y(_261_) );
NAND2X1 NAND2X1_142 ( .A(1'b0), .B(_15_), .Y(_262_) );
OAI21X1 OAI21X1_129 ( .A(_15_), .B(_261_), .C(_262_), .Y(w_cout_5_) );
INVX1 INVX1_128 ( .A(w_cout_5_), .Y(_267_) );
NAND2X1 NAND2X1_143 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_268_) );
BUFX2 BUFX2_59 ( .A(cskip1_inst_rca0_fa0_o_sum), .Y(_0__56_) );
BUFX2 BUFX2_60 ( .A(1'b0), .Y(w_cout_0_) );
BUFX2 BUFX2_61 ( .A(cskip1_inst_cin), .Y(w_cout_14_) );
endmodule
