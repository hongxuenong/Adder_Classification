module cla_51bit (i_add1, i_add2, o_result);

input [50:0] i_add1;
input [50:0] i_add2;
output [51:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

INVX1 INVX1_1 ( .A(_161_), .Y(_162_) );
NAND3X1 NAND3X1_1 ( .A(_160_), .B(_162_), .C(_153_), .Y(_163_) );
AND2X2 AND2X2_1 ( .A(_163_), .B(_158_), .Y(_164_) );
INVX1 INVX1_2 ( .A(_164_), .Y(w_C_27_) );
AND2X2 AND2X2_2 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_165_) );
INVX1 INVX1_3 ( .A(_165_), .Y(_166_) );
NAND3X1 NAND3X1_2 ( .A(_158_), .B(_166_), .C(_163_), .Y(_167_) );
OAI21X1 OAI21X1_1 ( .A(i_add2[27]), .B(i_add1[27]), .C(_167_), .Y(_168_) );
INVX1 INVX1_4 ( .A(_168_), .Y(w_C_28_) );
INVX1 INVX1_5 ( .A(i_add2[28]), .Y(_169_) );
INVX1 INVX1_6 ( .A(i_add1[28]), .Y(_170_) );
NOR2X1 NOR2X1_1 ( .A(_169_), .B(_170_), .Y(_171_) );
INVX1 INVX1_7 ( .A(_171_), .Y(_172_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_173_) );
INVX1 INVX1_8 ( .A(_173_), .Y(_174_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_175_) );
INVX1 INVX1_9 ( .A(_175_), .Y(_176_) );
NAND3X1 NAND3X1_3 ( .A(_174_), .B(_176_), .C(_167_), .Y(_177_) );
AND2X2 AND2X2_3 ( .A(_177_), .B(_172_), .Y(_178_) );
INVX1 INVX1_10 ( .A(_178_), .Y(w_C_29_) );
AND2X2 AND2X2_4 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_179_) );
BUFX2 BUFX2_1 ( .A(_306__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_306__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_306__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_306__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_306__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_306__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_306__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_306__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_306__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_306__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_306__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_306__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_306__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_306__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_306__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_306__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_306__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_306__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_306__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_306__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_306__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_306__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_306__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_306__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_306__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_306__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_306__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_306__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_306__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_306__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_306__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_306__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_306__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_306__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_306__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_306__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_306__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(_306__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .A(_306__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .A(_306__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .A(_306__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .A(_306__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .A(_306__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .A(_306__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .A(_306__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .A(_306__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .A(_306__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .A(_306__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .A(_306__48_), .Y(o_result[48]) );
BUFX2 BUFX2_50 ( .A(_306__49_), .Y(o_result[49]) );
BUFX2 BUFX2_51 ( .A(_306__50_), .Y(o_result[50]) );
BUFX2 BUFX2_52 ( .A(w_C_51_), .Y(o_result[51]) );
INVX1 INVX1_11 ( .A(w_C_4_), .Y(_310_) );
OR2X2 OR2X2_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_311_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_312_) );
NAND3X1 NAND3X1_4 ( .A(_310_), .B(_312_), .C(_311_), .Y(_313_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_307_) );
AND2X2 AND2X2_5 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_308_) );
OAI21X1 OAI21X1_2 ( .A(_307_), .B(_308_), .C(w_C_4_), .Y(_309_) );
NAND2X1 NAND2X1_2 ( .A(_309_), .B(_313_), .Y(_306__4_) );
INVX1 INVX1_12 ( .A(w_C_5_), .Y(_317_) );
OR2X2 OR2X2_2 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_318_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_319_) );
NAND3X1 NAND3X1_5 ( .A(_317_), .B(_319_), .C(_318_), .Y(_320_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_314_) );
AND2X2 AND2X2_6 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_315_) );
OAI21X1 OAI21X1_3 ( .A(_314_), .B(_315_), .C(w_C_5_), .Y(_316_) );
NAND2X1 NAND2X1_4 ( .A(_316_), .B(_320_), .Y(_306__5_) );
INVX1 INVX1_13 ( .A(w_C_6_), .Y(_324_) );
OR2X2 OR2X2_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_325_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_326_) );
NAND3X1 NAND3X1_6 ( .A(_324_), .B(_326_), .C(_325_), .Y(_327_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_321_) );
AND2X2 AND2X2_7 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_322_) );
OAI21X1 OAI21X1_4 ( .A(_321_), .B(_322_), .C(w_C_6_), .Y(_323_) );
NAND2X1 NAND2X1_6 ( .A(_323_), .B(_327_), .Y(_306__6_) );
INVX1 INVX1_14 ( .A(w_C_7_), .Y(_331_) );
OR2X2 OR2X2_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_332_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_333_) );
NAND3X1 NAND3X1_7 ( .A(_331_), .B(_333_), .C(_332_), .Y(_334_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_328_) );
AND2X2 AND2X2_8 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_329_) );
OAI21X1 OAI21X1_5 ( .A(_328_), .B(_329_), .C(w_C_7_), .Y(_330_) );
NAND2X1 NAND2X1_8 ( .A(_330_), .B(_334_), .Y(_306__7_) );
INVX1 INVX1_15 ( .A(w_C_8_), .Y(_338_) );
OR2X2 OR2X2_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_339_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_340_) );
NAND3X1 NAND3X1_8 ( .A(_338_), .B(_340_), .C(_339_), .Y(_341_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_335_) );
AND2X2 AND2X2_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_336_) );
OAI21X1 OAI21X1_6 ( .A(_335_), .B(_336_), .C(w_C_8_), .Y(_337_) );
NAND2X1 NAND2X1_10 ( .A(_337_), .B(_341_), .Y(_306__8_) );
INVX1 INVX1_16 ( .A(w_C_9_), .Y(_345_) );
OR2X2 OR2X2_6 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_346_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_347_) );
NAND3X1 NAND3X1_9 ( .A(_345_), .B(_347_), .C(_346_), .Y(_348_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_342_) );
AND2X2 AND2X2_10 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_343_) );
OAI21X1 OAI21X1_7 ( .A(_342_), .B(_343_), .C(w_C_9_), .Y(_344_) );
NAND2X1 NAND2X1_12 ( .A(_344_), .B(_348_), .Y(_306__9_) );
INVX1 INVX1_17 ( .A(w_C_10_), .Y(_352_) );
OR2X2 OR2X2_7 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_353_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_354_) );
NAND3X1 NAND3X1_10 ( .A(_352_), .B(_354_), .C(_353_), .Y(_355_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_349_) );
AND2X2 AND2X2_11 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_350_) );
OAI21X1 OAI21X1_8 ( .A(_349_), .B(_350_), .C(w_C_10_), .Y(_351_) );
NAND2X1 NAND2X1_14 ( .A(_351_), .B(_355_), .Y(_306__10_) );
INVX1 INVX1_18 ( .A(w_C_11_), .Y(_359_) );
OR2X2 OR2X2_8 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_360_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_361_) );
NAND3X1 NAND3X1_11 ( .A(_359_), .B(_361_), .C(_360_), .Y(_362_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_356_) );
AND2X2 AND2X2_12 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_357_) );
OAI21X1 OAI21X1_9 ( .A(_356_), .B(_357_), .C(w_C_11_), .Y(_358_) );
NAND2X1 NAND2X1_16 ( .A(_358_), .B(_362_), .Y(_306__11_) );
INVX1 INVX1_19 ( .A(w_C_12_), .Y(_366_) );
OR2X2 OR2X2_9 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_367_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_368_) );
NAND3X1 NAND3X1_12 ( .A(_366_), .B(_368_), .C(_367_), .Y(_369_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_363_) );
AND2X2 AND2X2_13 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_364_) );
OAI21X1 OAI21X1_10 ( .A(_363_), .B(_364_), .C(w_C_12_), .Y(_365_) );
NAND2X1 NAND2X1_18 ( .A(_365_), .B(_369_), .Y(_306__12_) );
INVX1 INVX1_20 ( .A(w_C_13_), .Y(_373_) );
OR2X2 OR2X2_10 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_374_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_375_) );
NAND3X1 NAND3X1_13 ( .A(_373_), .B(_375_), .C(_374_), .Y(_376_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_370_) );
AND2X2 AND2X2_14 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_371_) );
OAI21X1 OAI21X1_11 ( .A(_370_), .B(_371_), .C(w_C_13_), .Y(_372_) );
NAND2X1 NAND2X1_20 ( .A(_372_), .B(_376_), .Y(_306__13_) );
INVX1 INVX1_21 ( .A(w_C_14_), .Y(_380_) );
OR2X2 OR2X2_11 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_381_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_382_) );
NAND3X1 NAND3X1_14 ( .A(_380_), .B(_382_), .C(_381_), .Y(_383_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_377_) );
AND2X2 AND2X2_15 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_378_) );
OAI21X1 OAI21X1_12 ( .A(_377_), .B(_378_), .C(w_C_14_), .Y(_379_) );
NAND2X1 NAND2X1_22 ( .A(_379_), .B(_383_), .Y(_306__14_) );
INVX1 INVX1_22 ( .A(w_C_15_), .Y(_387_) );
OR2X2 OR2X2_12 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_388_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_389_) );
NAND3X1 NAND3X1_15 ( .A(_387_), .B(_389_), .C(_388_), .Y(_390_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_384_) );
AND2X2 AND2X2_16 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_385_) );
OAI21X1 OAI21X1_13 ( .A(_384_), .B(_385_), .C(w_C_15_), .Y(_386_) );
NAND2X1 NAND2X1_24 ( .A(_386_), .B(_390_), .Y(_306__15_) );
INVX1 INVX1_23 ( .A(w_C_16_), .Y(_394_) );
OR2X2 OR2X2_13 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_395_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_396_) );
NAND3X1 NAND3X1_16 ( .A(_394_), .B(_396_), .C(_395_), .Y(_397_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_391_) );
AND2X2 AND2X2_17 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_392_) );
OAI21X1 OAI21X1_14 ( .A(_391_), .B(_392_), .C(w_C_16_), .Y(_393_) );
NAND2X1 NAND2X1_26 ( .A(_393_), .B(_397_), .Y(_306__16_) );
INVX1 INVX1_24 ( .A(w_C_17_), .Y(_401_) );
OR2X2 OR2X2_14 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_402_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_403_) );
NAND3X1 NAND3X1_17 ( .A(_401_), .B(_403_), .C(_402_), .Y(_404_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_398_) );
AND2X2 AND2X2_18 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_399_) );
OAI21X1 OAI21X1_15 ( .A(_398_), .B(_399_), .C(w_C_17_), .Y(_400_) );
NAND2X1 NAND2X1_28 ( .A(_400_), .B(_404_), .Y(_306__17_) );
INVX1 INVX1_25 ( .A(w_C_18_), .Y(_408_) );
OR2X2 OR2X2_15 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_409_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_410_) );
NAND3X1 NAND3X1_18 ( .A(_408_), .B(_410_), .C(_409_), .Y(_411_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_405_) );
AND2X2 AND2X2_19 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_406_) );
OAI21X1 OAI21X1_16 ( .A(_405_), .B(_406_), .C(w_C_18_), .Y(_407_) );
NAND2X1 NAND2X1_30 ( .A(_407_), .B(_411_), .Y(_306__18_) );
INVX1 INVX1_26 ( .A(w_C_19_), .Y(_415_) );
OR2X2 OR2X2_16 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_416_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_417_) );
NAND3X1 NAND3X1_19 ( .A(_415_), .B(_417_), .C(_416_), .Y(_418_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_412_) );
AND2X2 AND2X2_20 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_413_) );
OAI21X1 OAI21X1_17 ( .A(_412_), .B(_413_), .C(w_C_19_), .Y(_414_) );
NAND2X1 NAND2X1_32 ( .A(_414_), .B(_418_), .Y(_306__19_) );
INVX1 INVX1_27 ( .A(w_C_20_), .Y(_422_) );
OR2X2 OR2X2_17 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_423_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_424_) );
NAND3X1 NAND3X1_20 ( .A(_422_), .B(_424_), .C(_423_), .Y(_425_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_419_) );
AND2X2 AND2X2_21 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_420_) );
OAI21X1 OAI21X1_18 ( .A(_419_), .B(_420_), .C(w_C_20_), .Y(_421_) );
NAND2X1 NAND2X1_34 ( .A(_421_), .B(_425_), .Y(_306__20_) );
INVX1 INVX1_28 ( .A(w_C_21_), .Y(_429_) );
OR2X2 OR2X2_18 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_430_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_431_) );
NAND3X1 NAND3X1_21 ( .A(_429_), .B(_431_), .C(_430_), .Y(_432_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_426_) );
AND2X2 AND2X2_22 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_427_) );
OAI21X1 OAI21X1_19 ( .A(_426_), .B(_427_), .C(w_C_21_), .Y(_428_) );
NAND2X1 NAND2X1_36 ( .A(_428_), .B(_432_), .Y(_306__21_) );
INVX1 INVX1_29 ( .A(w_C_22_), .Y(_436_) );
OR2X2 OR2X2_19 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_437_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_438_) );
NAND3X1 NAND3X1_22 ( .A(_436_), .B(_438_), .C(_437_), .Y(_439_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_433_) );
AND2X2 AND2X2_23 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_434_) );
OAI21X1 OAI21X1_20 ( .A(_433_), .B(_434_), .C(w_C_22_), .Y(_435_) );
NAND2X1 NAND2X1_38 ( .A(_435_), .B(_439_), .Y(_306__22_) );
INVX1 INVX1_30 ( .A(w_C_23_), .Y(_443_) );
OR2X2 OR2X2_20 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_444_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_445_) );
NAND3X1 NAND3X1_23 ( .A(_443_), .B(_445_), .C(_444_), .Y(_446_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_440_) );
AND2X2 AND2X2_24 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_441_) );
OAI21X1 OAI21X1_21 ( .A(_440_), .B(_441_), .C(w_C_23_), .Y(_442_) );
NAND2X1 NAND2X1_40 ( .A(_442_), .B(_446_), .Y(_306__23_) );
INVX1 INVX1_31 ( .A(w_C_24_), .Y(_450_) );
OR2X2 OR2X2_21 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_451_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_452_) );
NAND3X1 NAND3X1_24 ( .A(_450_), .B(_452_), .C(_451_), .Y(_453_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_447_) );
AND2X2 AND2X2_25 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_448_) );
OAI21X1 OAI21X1_22 ( .A(_447_), .B(_448_), .C(w_C_24_), .Y(_449_) );
NAND2X1 NAND2X1_42 ( .A(_449_), .B(_453_), .Y(_306__24_) );
INVX1 INVX1_32 ( .A(w_C_25_), .Y(_457_) );
OR2X2 OR2X2_22 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_458_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_459_) );
NAND3X1 NAND3X1_25 ( .A(_457_), .B(_459_), .C(_458_), .Y(_460_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_454_) );
AND2X2 AND2X2_26 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_455_) );
OAI21X1 OAI21X1_23 ( .A(_454_), .B(_455_), .C(w_C_25_), .Y(_456_) );
NAND2X1 NAND2X1_44 ( .A(_456_), .B(_460_), .Y(_306__25_) );
INVX1 INVX1_33 ( .A(w_C_26_), .Y(_464_) );
OR2X2 OR2X2_23 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_465_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_466_) );
NAND3X1 NAND3X1_26 ( .A(_464_), .B(_466_), .C(_465_), .Y(_467_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_461_) );
AND2X2 AND2X2_27 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_462_) );
OAI21X1 OAI21X1_24 ( .A(_461_), .B(_462_), .C(w_C_26_), .Y(_463_) );
NAND2X1 NAND2X1_46 ( .A(_463_), .B(_467_), .Y(_306__26_) );
INVX1 INVX1_34 ( .A(w_C_27_), .Y(_471_) );
OR2X2 OR2X2_24 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_472_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_473_) );
NAND3X1 NAND3X1_27 ( .A(_471_), .B(_473_), .C(_472_), .Y(_474_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_468_) );
AND2X2 AND2X2_28 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_469_) );
OAI21X1 OAI21X1_25 ( .A(_468_), .B(_469_), .C(w_C_27_), .Y(_470_) );
NAND2X1 NAND2X1_48 ( .A(_470_), .B(_474_), .Y(_306__27_) );
INVX1 INVX1_35 ( .A(w_C_28_), .Y(_478_) );
OR2X2 OR2X2_25 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_479_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_480_) );
NAND3X1 NAND3X1_28 ( .A(_478_), .B(_480_), .C(_479_), .Y(_481_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_475_) );
AND2X2 AND2X2_29 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_476_) );
OAI21X1 OAI21X1_26 ( .A(_475_), .B(_476_), .C(w_C_28_), .Y(_477_) );
NAND2X1 NAND2X1_50 ( .A(_477_), .B(_481_), .Y(_306__28_) );
INVX1 INVX1_36 ( .A(w_C_29_), .Y(_485_) );
OR2X2 OR2X2_26 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_486_) );
NAND2X1 NAND2X1_51 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_487_) );
NAND3X1 NAND3X1_29 ( .A(_485_), .B(_487_), .C(_486_), .Y(_488_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_482_) );
AND2X2 AND2X2_30 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_483_) );
OAI21X1 OAI21X1_27 ( .A(_482_), .B(_483_), .C(w_C_29_), .Y(_484_) );
NAND2X1 NAND2X1_52 ( .A(_484_), .B(_488_), .Y(_306__29_) );
INVX1 INVX1_37 ( .A(w_C_30_), .Y(_492_) );
OR2X2 OR2X2_27 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_493_) );
NAND2X1 NAND2X1_53 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_494_) );
NAND3X1 NAND3X1_30 ( .A(_492_), .B(_494_), .C(_493_), .Y(_495_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_489_) );
AND2X2 AND2X2_31 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_490_) );
OAI21X1 OAI21X1_28 ( .A(_489_), .B(_490_), .C(w_C_30_), .Y(_491_) );
NAND2X1 NAND2X1_54 ( .A(_491_), .B(_495_), .Y(_306__30_) );
INVX1 INVX1_38 ( .A(w_C_31_), .Y(_499_) );
OR2X2 OR2X2_28 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_500_) );
NAND2X1 NAND2X1_55 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_501_) );
NAND3X1 NAND3X1_31 ( .A(_499_), .B(_501_), .C(_500_), .Y(_502_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_496_) );
AND2X2 AND2X2_32 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_497_) );
OAI21X1 OAI21X1_29 ( .A(_496_), .B(_497_), .C(w_C_31_), .Y(_498_) );
NAND2X1 NAND2X1_56 ( .A(_498_), .B(_502_), .Y(_306__31_) );
INVX1 INVX1_39 ( .A(w_C_32_), .Y(_506_) );
OR2X2 OR2X2_29 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_507_) );
NAND2X1 NAND2X1_57 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_508_) );
NAND3X1 NAND3X1_32 ( .A(_506_), .B(_508_), .C(_507_), .Y(_509_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_503_) );
AND2X2 AND2X2_33 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_504_) );
OAI21X1 OAI21X1_30 ( .A(_503_), .B(_504_), .C(w_C_32_), .Y(_505_) );
NAND2X1 NAND2X1_58 ( .A(_505_), .B(_509_), .Y(_306__32_) );
INVX1 INVX1_40 ( .A(w_C_33_), .Y(_513_) );
OR2X2 OR2X2_30 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_514_) );
NAND2X1 NAND2X1_59 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_515_) );
NAND3X1 NAND3X1_33 ( .A(_513_), .B(_515_), .C(_514_), .Y(_516_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_510_) );
AND2X2 AND2X2_34 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_511_) );
OAI21X1 OAI21X1_31 ( .A(_510_), .B(_511_), .C(w_C_33_), .Y(_512_) );
NAND2X1 NAND2X1_60 ( .A(_512_), .B(_516_), .Y(_306__33_) );
INVX1 INVX1_41 ( .A(w_C_34_), .Y(_520_) );
OR2X2 OR2X2_31 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_521_) );
NAND2X1 NAND2X1_61 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_522_) );
NAND3X1 NAND3X1_34 ( .A(_520_), .B(_522_), .C(_521_), .Y(_523_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_517_) );
AND2X2 AND2X2_35 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_518_) );
OAI21X1 OAI21X1_32 ( .A(_517_), .B(_518_), .C(w_C_34_), .Y(_519_) );
NAND2X1 NAND2X1_62 ( .A(_519_), .B(_523_), .Y(_306__34_) );
INVX1 INVX1_42 ( .A(w_C_35_), .Y(_527_) );
OR2X2 OR2X2_32 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_528_) );
NAND2X1 NAND2X1_63 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_529_) );
NAND3X1 NAND3X1_35 ( .A(_527_), .B(_529_), .C(_528_), .Y(_530_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_524_) );
AND2X2 AND2X2_36 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_525_) );
OAI21X1 OAI21X1_33 ( .A(_524_), .B(_525_), .C(w_C_35_), .Y(_526_) );
NAND2X1 NAND2X1_64 ( .A(_526_), .B(_530_), .Y(_306__35_) );
INVX1 INVX1_43 ( .A(w_C_36_), .Y(_534_) );
OR2X2 OR2X2_33 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_535_) );
NAND2X1 NAND2X1_65 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_536_) );
NAND3X1 NAND3X1_36 ( .A(_534_), .B(_536_), .C(_535_), .Y(_537_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_531_) );
AND2X2 AND2X2_37 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_532_) );
OAI21X1 OAI21X1_34 ( .A(_531_), .B(_532_), .C(w_C_36_), .Y(_533_) );
NAND2X1 NAND2X1_66 ( .A(_533_), .B(_537_), .Y(_306__36_) );
INVX1 INVX1_44 ( .A(w_C_37_), .Y(_541_) );
OR2X2 OR2X2_34 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_542_) );
NAND2X1 NAND2X1_67 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_543_) );
NAND3X1 NAND3X1_37 ( .A(_541_), .B(_543_), .C(_542_), .Y(_544_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_538_) );
AND2X2 AND2X2_38 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_539_) );
OAI21X1 OAI21X1_35 ( .A(_538_), .B(_539_), .C(w_C_37_), .Y(_540_) );
NAND2X1 NAND2X1_68 ( .A(_540_), .B(_544_), .Y(_306__37_) );
INVX1 INVX1_45 ( .A(w_C_38_), .Y(_548_) );
OR2X2 OR2X2_35 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_549_) );
NAND2X1 NAND2X1_69 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_550_) );
NAND3X1 NAND3X1_38 ( .A(_548_), .B(_550_), .C(_549_), .Y(_551_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_545_) );
AND2X2 AND2X2_39 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_546_) );
OAI21X1 OAI21X1_36 ( .A(_545_), .B(_546_), .C(w_C_38_), .Y(_547_) );
NAND2X1 NAND2X1_70 ( .A(_547_), .B(_551_), .Y(_306__38_) );
INVX1 INVX1_46 ( .A(w_C_39_), .Y(_555_) );
OR2X2 OR2X2_36 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_556_) );
NAND2X1 NAND2X1_71 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_557_) );
NAND3X1 NAND3X1_39 ( .A(_555_), .B(_557_), .C(_556_), .Y(_558_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_552_) );
AND2X2 AND2X2_40 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_553_) );
OAI21X1 OAI21X1_37 ( .A(_552_), .B(_553_), .C(w_C_39_), .Y(_554_) );
NAND2X1 NAND2X1_72 ( .A(_554_), .B(_558_), .Y(_306__39_) );
INVX1 INVX1_47 ( .A(w_C_40_), .Y(_562_) );
OR2X2 OR2X2_37 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_563_) );
NAND2X1 NAND2X1_73 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_564_) );
NAND3X1 NAND3X1_40 ( .A(_562_), .B(_564_), .C(_563_), .Y(_565_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_559_) );
AND2X2 AND2X2_41 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_560_) );
OAI21X1 OAI21X1_38 ( .A(_559_), .B(_560_), .C(w_C_40_), .Y(_561_) );
NAND2X1 NAND2X1_74 ( .A(_561_), .B(_565_), .Y(_306__40_) );
INVX1 INVX1_48 ( .A(w_C_41_), .Y(_569_) );
OR2X2 OR2X2_38 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_570_) );
NAND2X1 NAND2X1_75 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_571_) );
NAND3X1 NAND3X1_41 ( .A(_569_), .B(_571_), .C(_570_), .Y(_572_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_566_) );
AND2X2 AND2X2_42 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_567_) );
OAI21X1 OAI21X1_39 ( .A(_566_), .B(_567_), .C(w_C_41_), .Y(_568_) );
NAND2X1 NAND2X1_76 ( .A(_568_), .B(_572_), .Y(_306__41_) );
INVX1 INVX1_49 ( .A(w_C_42_), .Y(_576_) );
OR2X2 OR2X2_39 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_577_) );
NAND2X1 NAND2X1_77 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_578_) );
NAND3X1 NAND3X1_42 ( .A(_576_), .B(_578_), .C(_577_), .Y(_579_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_573_) );
AND2X2 AND2X2_43 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_574_) );
OAI21X1 OAI21X1_40 ( .A(_573_), .B(_574_), .C(w_C_42_), .Y(_575_) );
NAND2X1 NAND2X1_78 ( .A(_575_), .B(_579_), .Y(_306__42_) );
INVX1 INVX1_50 ( .A(w_C_43_), .Y(_583_) );
OR2X2 OR2X2_40 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_584_) );
NAND2X1 NAND2X1_79 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_585_) );
NAND3X1 NAND3X1_43 ( .A(_583_), .B(_585_), .C(_584_), .Y(_586_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_580_) );
AND2X2 AND2X2_44 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_581_) );
OAI21X1 OAI21X1_41 ( .A(_580_), .B(_581_), .C(w_C_43_), .Y(_582_) );
NAND2X1 NAND2X1_80 ( .A(_582_), .B(_586_), .Y(_306__43_) );
INVX1 INVX1_51 ( .A(w_C_44_), .Y(_590_) );
OR2X2 OR2X2_41 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_591_) );
NAND2X1 NAND2X1_81 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_592_) );
NAND3X1 NAND3X1_44 ( .A(_590_), .B(_592_), .C(_591_), .Y(_593_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_587_) );
AND2X2 AND2X2_45 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_588_) );
OAI21X1 OAI21X1_42 ( .A(_587_), .B(_588_), .C(w_C_44_), .Y(_589_) );
NAND2X1 NAND2X1_82 ( .A(_589_), .B(_593_), .Y(_306__44_) );
INVX1 INVX1_52 ( .A(w_C_45_), .Y(_597_) );
OR2X2 OR2X2_42 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_598_) );
NAND2X1 NAND2X1_83 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_599_) );
NAND3X1 NAND3X1_45 ( .A(_597_), .B(_599_), .C(_598_), .Y(_600_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_594_) );
AND2X2 AND2X2_46 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_595_) );
OAI21X1 OAI21X1_43 ( .A(_594_), .B(_595_), .C(w_C_45_), .Y(_596_) );
NAND2X1 NAND2X1_84 ( .A(_596_), .B(_600_), .Y(_306__45_) );
INVX1 INVX1_53 ( .A(w_C_46_), .Y(_604_) );
OR2X2 OR2X2_43 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_605_) );
NAND2X1 NAND2X1_85 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_606_) );
NAND3X1 NAND3X1_46 ( .A(_604_), .B(_606_), .C(_605_), .Y(_607_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_601_) );
AND2X2 AND2X2_47 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_602_) );
OAI21X1 OAI21X1_44 ( .A(_601_), .B(_602_), .C(w_C_46_), .Y(_603_) );
NAND2X1 NAND2X1_86 ( .A(_603_), .B(_607_), .Y(_306__46_) );
INVX1 INVX1_54 ( .A(w_C_47_), .Y(_611_) );
OR2X2 OR2X2_44 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_612_) );
NAND2X1 NAND2X1_87 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_613_) );
NAND3X1 NAND3X1_47 ( .A(_611_), .B(_613_), .C(_612_), .Y(_614_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_608_) );
AND2X2 AND2X2_48 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_609_) );
OAI21X1 OAI21X1_45 ( .A(_608_), .B(_609_), .C(w_C_47_), .Y(_610_) );
NAND2X1 NAND2X1_88 ( .A(_610_), .B(_614_), .Y(_306__47_) );
INVX1 INVX1_55 ( .A(w_C_48_), .Y(_618_) );
OR2X2 OR2X2_45 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_619_) );
NAND2X1 NAND2X1_89 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_620_) );
NAND3X1 NAND3X1_48 ( .A(_618_), .B(_620_), .C(_619_), .Y(_621_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_615_) );
AND2X2 AND2X2_49 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_616_) );
OAI21X1 OAI21X1_46 ( .A(_615_), .B(_616_), .C(w_C_48_), .Y(_617_) );
NAND2X1 NAND2X1_90 ( .A(_617_), .B(_621_), .Y(_306__48_) );
INVX1 INVX1_56 ( .A(w_C_49_), .Y(_625_) );
OR2X2 OR2X2_46 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_626_) );
NAND2X1 NAND2X1_91 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_627_) );
NAND3X1 NAND3X1_49 ( .A(_625_), .B(_627_), .C(_626_), .Y(_628_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_622_) );
AND2X2 AND2X2_50 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_623_) );
OAI21X1 OAI21X1_47 ( .A(_622_), .B(_623_), .C(w_C_49_), .Y(_624_) );
NAND2X1 NAND2X1_92 ( .A(_624_), .B(_628_), .Y(_306__49_) );
INVX1 INVX1_57 ( .A(w_C_50_), .Y(_632_) );
OR2X2 OR2X2_47 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_633_) );
NAND2X1 NAND2X1_93 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_634_) );
NAND3X1 NAND3X1_50 ( .A(_632_), .B(_634_), .C(_633_), .Y(_635_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_629_) );
AND2X2 AND2X2_51 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_630_) );
OAI21X1 OAI21X1_48 ( .A(_629_), .B(_630_), .C(w_C_50_), .Y(_631_) );
NAND2X1 NAND2X1_94 ( .A(_631_), .B(_635_), .Y(_306__50_) );
INVX1 INVX1_58 ( .A(gnd), .Y(_639_) );
OR2X2 OR2X2_48 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_640_) );
NAND2X1 NAND2X1_95 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_641_) );
NAND3X1 NAND3X1_51 ( .A(_639_), .B(_641_), .C(_640_), .Y(_642_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_636_) );
AND2X2 AND2X2_52 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_637_) );
OAI21X1 OAI21X1_49 ( .A(_636_), .B(_637_), .C(gnd), .Y(_638_) );
NAND2X1 NAND2X1_96 ( .A(_638_), .B(_642_), .Y(_306__0_) );
INVX1 INVX1_59 ( .A(w_C_1_), .Y(_646_) );
OR2X2 OR2X2_49 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_647_) );
NAND2X1 NAND2X1_97 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_648_) );
NAND3X1 NAND3X1_52 ( .A(_646_), .B(_648_), .C(_647_), .Y(_649_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_643_) );
AND2X2 AND2X2_53 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_644_) );
OAI21X1 OAI21X1_50 ( .A(_643_), .B(_644_), .C(w_C_1_), .Y(_645_) );
NAND2X1 NAND2X1_98 ( .A(_645_), .B(_649_), .Y(_306__1_) );
INVX1 INVX1_60 ( .A(w_C_2_), .Y(_653_) );
OR2X2 OR2X2_50 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_654_) );
NAND2X1 NAND2X1_99 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_655_) );
NAND3X1 NAND3X1_53 ( .A(_653_), .B(_655_), .C(_654_), .Y(_656_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_650_) );
AND2X2 AND2X2_54 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_651_) );
OAI21X1 OAI21X1_51 ( .A(_650_), .B(_651_), .C(w_C_2_), .Y(_652_) );
NAND2X1 NAND2X1_100 ( .A(_652_), .B(_656_), .Y(_306__2_) );
INVX1 INVX1_61 ( .A(w_C_3_), .Y(_660_) );
OR2X2 OR2X2_51 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_661_) );
NAND2X1 NAND2X1_101 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_662_) );
NAND3X1 NAND3X1_54 ( .A(_660_), .B(_662_), .C(_661_), .Y(_663_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_657_) );
AND2X2 AND2X2_55 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_658_) );
OAI21X1 OAI21X1_52 ( .A(_657_), .B(_658_), .C(w_C_3_), .Y(_659_) );
NAND2X1 NAND2X1_102 ( .A(_659_), .B(_663_), .Y(_306__3_) );
INVX1 INVX1_62 ( .A(_179_), .Y(_180_) );
NAND3X1 NAND3X1_55 ( .A(_172_), .B(_180_), .C(_177_), .Y(_181_) );
OAI21X1 OAI21X1_53 ( .A(i_add2[29]), .B(i_add1[29]), .C(_181_), .Y(_182_) );
INVX1 INVX1_63 ( .A(_182_), .Y(w_C_30_) );
INVX1 INVX1_64 ( .A(i_add2[30]), .Y(_183_) );
INVX1 INVX1_65 ( .A(i_add1[30]), .Y(_184_) );
NOR2X1 NOR2X1_55 ( .A(_183_), .B(_184_), .Y(_185_) );
INVX1 INVX1_66 ( .A(_185_), .Y(_186_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_187_) );
INVX1 INVX1_67 ( .A(_187_), .Y(_188_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_189_) );
INVX1 INVX1_68 ( .A(_189_), .Y(_190_) );
NAND3X1 NAND3X1_56 ( .A(_188_), .B(_190_), .C(_181_), .Y(_191_) );
AND2X2 AND2X2_56 ( .A(_191_), .B(_186_), .Y(_192_) );
INVX1 INVX1_69 ( .A(_192_), .Y(w_C_31_) );
AND2X2 AND2X2_57 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_193_) );
INVX1 INVX1_70 ( .A(_193_), .Y(_194_) );
NAND3X1 NAND3X1_57 ( .A(_186_), .B(_194_), .C(_191_), .Y(_195_) );
OAI21X1 OAI21X1_54 ( .A(i_add2[31]), .B(i_add1[31]), .C(_195_), .Y(_196_) );
INVX1 INVX1_71 ( .A(_196_), .Y(w_C_32_) );
INVX1 INVX1_72 ( .A(i_add2[32]), .Y(_197_) );
INVX1 INVX1_73 ( .A(i_add1[32]), .Y(_198_) );
NOR2X1 NOR2X1_58 ( .A(_197_), .B(_198_), .Y(_199_) );
INVX1 INVX1_74 ( .A(_199_), .Y(_200_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_201_) );
INVX1 INVX1_75 ( .A(_201_), .Y(_202_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_203_) );
INVX1 INVX1_76 ( .A(_203_), .Y(_204_) );
NAND3X1 NAND3X1_58 ( .A(_202_), .B(_204_), .C(_195_), .Y(_205_) );
AND2X2 AND2X2_58 ( .A(_205_), .B(_200_), .Y(_206_) );
INVX1 INVX1_77 ( .A(_206_), .Y(w_C_33_) );
AND2X2 AND2X2_59 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_207_) );
INVX1 INVX1_78 ( .A(_207_), .Y(_208_) );
NAND3X1 NAND3X1_59 ( .A(_200_), .B(_208_), .C(_205_), .Y(_209_) );
OAI21X1 OAI21X1_55 ( .A(i_add2[33]), .B(i_add1[33]), .C(_209_), .Y(_210_) );
INVX1 INVX1_79 ( .A(_210_), .Y(w_C_34_) );
INVX1 INVX1_80 ( .A(i_add2[34]), .Y(_211_) );
INVX1 INVX1_81 ( .A(i_add1[34]), .Y(_212_) );
NOR2X1 NOR2X1_61 ( .A(_211_), .B(_212_), .Y(_213_) );
INVX1 INVX1_82 ( .A(_213_), .Y(_214_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_215_) );
INVX1 INVX1_83 ( .A(_215_), .Y(_216_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_217_) );
INVX1 INVX1_84 ( .A(_217_), .Y(_218_) );
NAND3X1 NAND3X1_60 ( .A(_216_), .B(_218_), .C(_209_), .Y(_219_) );
AND2X2 AND2X2_60 ( .A(_219_), .B(_214_), .Y(_220_) );
INVX1 INVX1_85 ( .A(_220_), .Y(w_C_35_) );
AND2X2 AND2X2_61 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_221_) );
INVX1 INVX1_86 ( .A(_221_), .Y(_222_) );
NAND3X1 NAND3X1_61 ( .A(_214_), .B(_222_), .C(_219_), .Y(_223_) );
OAI21X1 OAI21X1_56 ( .A(i_add2[35]), .B(i_add1[35]), .C(_223_), .Y(_224_) );
INVX1 INVX1_87 ( .A(_224_), .Y(w_C_36_) );
INVX1 INVX1_88 ( .A(i_add2[36]), .Y(_225_) );
INVX1 INVX1_89 ( .A(i_add1[36]), .Y(_226_) );
NOR2X1 NOR2X1_64 ( .A(_225_), .B(_226_), .Y(_227_) );
INVX1 INVX1_90 ( .A(_227_), .Y(_228_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_229_) );
INVX1 INVX1_91 ( .A(_229_), .Y(_230_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_231_) );
INVX1 INVX1_92 ( .A(_231_), .Y(_232_) );
NAND3X1 NAND3X1_62 ( .A(_230_), .B(_232_), .C(_223_), .Y(_233_) );
AND2X2 AND2X2_62 ( .A(_233_), .B(_228_), .Y(_234_) );
INVX1 INVX1_93 ( .A(_234_), .Y(w_C_37_) );
AND2X2 AND2X2_63 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_235_) );
INVX1 INVX1_94 ( .A(_235_), .Y(_236_) );
NAND3X1 NAND3X1_63 ( .A(_228_), .B(_236_), .C(_233_), .Y(_237_) );
OAI21X1 OAI21X1_57 ( .A(i_add2[37]), .B(i_add1[37]), .C(_237_), .Y(_238_) );
INVX1 INVX1_95 ( .A(_238_), .Y(w_C_38_) );
INVX1 INVX1_96 ( .A(i_add2[38]), .Y(_239_) );
INVX1 INVX1_97 ( .A(i_add1[38]), .Y(_240_) );
NOR2X1 NOR2X1_67 ( .A(_239_), .B(_240_), .Y(_241_) );
INVX1 INVX1_98 ( .A(_241_), .Y(_242_) );
NOR2X1 NOR2X1_68 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_243_) );
INVX1 INVX1_99 ( .A(_243_), .Y(_244_) );
NOR2X1 NOR2X1_69 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_245_) );
INVX1 INVX1_100 ( .A(_245_), .Y(_246_) );
NAND3X1 NAND3X1_64 ( .A(_244_), .B(_246_), .C(_237_), .Y(_247_) );
AND2X2 AND2X2_64 ( .A(_247_), .B(_242_), .Y(_248_) );
INVX1 INVX1_101 ( .A(_248_), .Y(w_C_39_) );
AND2X2 AND2X2_65 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_249_) );
INVX1 INVX1_102 ( .A(_249_), .Y(_250_) );
NAND3X1 NAND3X1_65 ( .A(_242_), .B(_250_), .C(_247_), .Y(_251_) );
OAI21X1 OAI21X1_58 ( .A(i_add2[39]), .B(i_add1[39]), .C(_251_), .Y(_252_) );
INVX1 INVX1_103 ( .A(_252_), .Y(w_C_40_) );
NAND2X1 NAND2X1_103 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_253_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_254_) );
OAI21X1 OAI21X1_59 ( .A(_254_), .B(_252_), .C(_253_), .Y(w_C_41_) );
OR2X2 OR2X2_52 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_255_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_256_) );
INVX1 INVX1_104 ( .A(_256_), .Y(_257_) );
INVX1 INVX1_105 ( .A(_254_), .Y(_258_) );
NAND3X1 NAND3X1_66 ( .A(_257_), .B(_258_), .C(_251_), .Y(_259_) );
NAND2X1 NAND2X1_104 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_260_) );
NAND3X1 NAND3X1_67 ( .A(_253_), .B(_260_), .C(_259_), .Y(_261_) );
AND2X2 AND2X2_66 ( .A(_261_), .B(_255_), .Y(w_C_42_) );
INVX1 INVX1_106 ( .A(i_add2[42]), .Y(_262_) );
INVX1 INVX1_107 ( .A(i_add1[42]), .Y(_263_) );
NAND2X1 NAND2X1_105 ( .A(_262_), .B(_263_), .Y(_264_) );
NAND3X1 NAND3X1_68 ( .A(_255_), .B(_264_), .C(_261_), .Y(_265_) );
OAI21X1 OAI21X1_60 ( .A(_262_), .B(_263_), .C(_265_), .Y(w_C_43_) );
INVX1 INVX1_108 ( .A(i_add2[43]), .Y(_266_) );
INVX1 INVX1_109 ( .A(i_add1[43]), .Y(_267_) );
NAND2X1 NAND2X1_106 ( .A(_266_), .B(_267_), .Y(_268_) );
NAND2X1 NAND2X1_107 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_269_) );
NAND2X1 NAND2X1_108 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_270_) );
NAND3X1 NAND3X1_69 ( .A(_269_), .B(_270_), .C(_265_), .Y(_271_) );
AND2X2 AND2X2_67 ( .A(_271_), .B(_268_), .Y(w_C_44_) );
INVX1 INVX1_110 ( .A(i_add2[44]), .Y(_272_) );
INVX1 INVX1_111 ( .A(i_add1[44]), .Y(_273_) );
NAND2X1 NAND2X1_109 ( .A(_272_), .B(_273_), .Y(_274_) );
NAND3X1 NAND3X1_70 ( .A(_268_), .B(_274_), .C(_271_), .Y(_275_) );
OAI21X1 OAI21X1_61 ( .A(_272_), .B(_273_), .C(_275_), .Y(w_C_45_) );
INVX1 INVX1_112 ( .A(i_add2[45]), .Y(_276_) );
INVX1 INVX1_113 ( .A(i_add1[45]), .Y(_277_) );
OAI21X1 OAI21X1_62 ( .A(i_add2[45]), .B(i_add1[45]), .C(w_C_45_), .Y(_278_) );
OAI21X1 OAI21X1_63 ( .A(_276_), .B(_277_), .C(_278_), .Y(w_C_46_) );
NOR2X1 NOR2X1_72 ( .A(_276_), .B(_277_), .Y(_279_) );
INVX1 INVX1_114 ( .A(_279_), .Y(_280_) );
AND2X2 AND2X2_68 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_281_) );
INVX1 INVX1_115 ( .A(_281_), .Y(_282_) );
NAND3X1 NAND3X1_71 ( .A(_280_), .B(_282_), .C(_278_), .Y(_283_) );
OAI21X1 OAI21X1_64 ( .A(i_add2[46]), .B(i_add1[46]), .C(_283_), .Y(_284_) );
INVX1 INVX1_116 ( .A(_284_), .Y(w_C_47_) );
NAND2X1 NAND2X1_110 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_285_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_286_) );
OAI21X1 OAI21X1_65 ( .A(_286_), .B(_284_), .C(_285_), .Y(w_C_48_) );
NAND2X1 NAND2X1_111 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_287_) );
INVX1 INVX1_117 ( .A(_286_), .Y(_288_) );
NOR2X1 NOR2X1_74 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_289_) );
INVX1 INVX1_118 ( .A(_289_), .Y(_290_) );
NOR2X1 NOR2X1_75 ( .A(_272_), .B(_273_), .Y(_291_) );
INVX1 INVX1_119 ( .A(_291_), .Y(_292_) );
NAND3X1 NAND3X1_72 ( .A(_292_), .B(_280_), .C(_275_), .Y(_293_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_294_) );
INVX1 INVX1_120 ( .A(_294_), .Y(_295_) );
NAND3X1 NAND3X1_73 ( .A(_290_), .B(_295_), .C(_293_), .Y(_296_) );
NAND3X1 NAND3X1_74 ( .A(_282_), .B(_285_), .C(_296_), .Y(_297_) );
OR2X2 OR2X2_53 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_298_) );
NAND3X1 NAND3X1_75 ( .A(_288_), .B(_298_), .C(_297_), .Y(_299_) );
NAND2X1 NAND2X1_112 ( .A(_287_), .B(_299_), .Y(w_C_49_) );
OR2X2 OR2X2_54 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_300_) );
NAND2X1 NAND2X1_113 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_301_) );
NAND3X1 NAND3X1_76 ( .A(_287_), .B(_301_), .C(_299_), .Y(_302_) );
AND2X2 AND2X2_69 ( .A(_302_), .B(_300_), .Y(w_C_50_) );
NAND2X1 NAND2X1_114 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_303_) );
OR2X2 OR2X2_55 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_304_) );
NAND3X1 NAND3X1_77 ( .A(_300_), .B(_304_), .C(_302_), .Y(_305_) );
NAND2X1 NAND2X1_115 ( .A(_303_), .B(_305_), .Y(w_C_51_) );
NAND2X1 NAND2X1_116 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_121 ( .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_117 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_118 ( .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_66 ( .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_122 ( .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_119 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_56 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_57 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_78 ( .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_120 ( .A(_4_), .B(_7_), .Y(w_C_3_) );
NAND2X1 NAND2X1_121 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
NAND3X1 NAND3X1_79 ( .A(_4_), .B(_8_), .C(_7_), .Y(_9_) );
OAI21X1 OAI21X1_67 ( .A(i_add2[3]), .B(i_add1[3]), .C(_9_), .Y(_10_) );
INVX1 INVX1_123 ( .A(_10_), .Y(w_C_4_) );
NAND2X1 NAND2X1_122 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
OR2X2 OR2X2_58 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_12_) );
OR2X2 OR2X2_59 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
NAND3X1 NAND3X1_80 ( .A(_12_), .B(_13_), .C(_9_), .Y(_14_) );
NAND2X1 NAND2X1_123 ( .A(_11_), .B(_14_), .Y(w_C_5_) );
NAND2X1 NAND2X1_124 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_15_) );
NAND3X1 NAND3X1_81 ( .A(_11_), .B(_15_), .C(_14_), .Y(_16_) );
OAI21X1 OAI21X1_68 ( .A(i_add2[5]), .B(i_add1[5]), .C(_16_), .Y(_17_) );
INVX1 INVX1_124 ( .A(_17_), .Y(w_C_6_) );
INVX1 INVX1_125 ( .A(i_add2[6]), .Y(_18_) );
INVX1 INVX1_126 ( .A(i_add1[6]), .Y(_19_) );
NOR2X1 NOR2X1_77 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_20_) );
INVX1 INVX1_127 ( .A(_20_), .Y(_21_) );
NOR2X1 NOR2X1_78 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_128 ( .A(_22_), .Y(_23_) );
NAND3X1 NAND3X1_82 ( .A(_21_), .B(_23_), .C(_16_), .Y(_24_) );
OAI21X1 OAI21X1_69 ( .A(_18_), .B(_19_), .C(_24_), .Y(w_C_7_) );
NOR2X1 NOR2X1_79 ( .A(_18_), .B(_19_), .Y(_25_) );
INVX1 INVX1_129 ( .A(_25_), .Y(_26_) );
AND2X2 AND2X2_70 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_27_) );
INVX1 INVX1_130 ( .A(_27_), .Y(_28_) );
NAND3X1 NAND3X1_83 ( .A(_26_), .B(_28_), .C(_24_), .Y(_29_) );
OAI21X1 OAI21X1_70 ( .A(i_add2[7]), .B(i_add1[7]), .C(_29_), .Y(_30_) );
INVX1 INVX1_131 ( .A(_30_), .Y(w_C_8_) );
INVX1 INVX1_132 ( .A(i_add2[8]), .Y(_31_) );
INVX1 INVX1_133 ( .A(i_add1[8]), .Y(_32_) );
NOR2X1 NOR2X1_80 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_33_) );
INVX1 INVX1_134 ( .A(_33_), .Y(_34_) );
NOR2X1 NOR2X1_81 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_35_) );
INVX1 INVX1_135 ( .A(_35_), .Y(_36_) );
NAND3X1 NAND3X1_84 ( .A(_34_), .B(_36_), .C(_29_), .Y(_37_) );
OAI21X1 OAI21X1_71 ( .A(_31_), .B(_32_), .C(_37_), .Y(w_C_9_) );
NOR2X1 NOR2X1_82 ( .A(_31_), .B(_32_), .Y(_38_) );
INVX1 INVX1_136 ( .A(_38_), .Y(_39_) );
AND2X2 AND2X2_71 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_40_) );
INVX1 INVX1_137 ( .A(_40_), .Y(_41_) );
NAND3X1 NAND3X1_85 ( .A(_39_), .B(_41_), .C(_37_), .Y(_42_) );
OAI21X1 OAI21X1_72 ( .A(i_add2[9]), .B(i_add1[9]), .C(_42_), .Y(_43_) );
INVX1 INVX1_138 ( .A(_43_), .Y(w_C_10_) );
INVX1 INVX1_139 ( .A(i_add2[10]), .Y(_44_) );
INVX1 INVX1_140 ( .A(i_add1[10]), .Y(_45_) );
NOR2X1 NOR2X1_83 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_46_) );
INVX1 INVX1_141 ( .A(_46_), .Y(_47_) );
NOR2X1 NOR2X1_84 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_48_) );
INVX1 INVX1_142 ( .A(_48_), .Y(_49_) );
NAND3X1 NAND3X1_86 ( .A(_47_), .B(_49_), .C(_42_), .Y(_50_) );
OAI21X1 OAI21X1_73 ( .A(_44_), .B(_45_), .C(_50_), .Y(w_C_11_) );
NOR2X1 NOR2X1_85 ( .A(_44_), .B(_45_), .Y(_51_) );
INVX1 INVX1_143 ( .A(_51_), .Y(_52_) );
AND2X2 AND2X2_72 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_53_) );
INVX1 INVX1_144 ( .A(_53_), .Y(_54_) );
NAND3X1 NAND3X1_87 ( .A(_52_), .B(_54_), .C(_50_), .Y(_55_) );
OAI21X1 OAI21X1_74 ( .A(i_add2[11]), .B(i_add1[11]), .C(_55_), .Y(_56_) );
INVX1 INVX1_145 ( .A(_56_), .Y(w_C_12_) );
INVX1 INVX1_146 ( .A(i_add2[12]), .Y(_57_) );
INVX1 INVX1_147 ( .A(i_add1[12]), .Y(_58_) );
NOR2X1 NOR2X1_86 ( .A(_57_), .B(_58_), .Y(_59_) );
INVX1 INVX1_148 ( .A(_59_), .Y(_60_) );
NOR2X1 NOR2X1_87 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_61_) );
INVX1 INVX1_149 ( .A(_61_), .Y(_62_) );
NOR2X1 NOR2X1_88 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_63_) );
INVX1 INVX1_150 ( .A(_63_), .Y(_64_) );
NAND3X1 NAND3X1_88 ( .A(_62_), .B(_64_), .C(_55_), .Y(_65_) );
AND2X2 AND2X2_73 ( .A(_65_), .B(_60_), .Y(_66_) );
INVX1 INVX1_151 ( .A(_66_), .Y(w_C_13_) );
AND2X2 AND2X2_74 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_67_) );
INVX1 INVX1_152 ( .A(_67_), .Y(_68_) );
NAND3X1 NAND3X1_89 ( .A(_60_), .B(_68_), .C(_65_), .Y(_69_) );
OAI21X1 OAI21X1_75 ( .A(i_add2[13]), .B(i_add1[13]), .C(_69_), .Y(_70_) );
INVX1 INVX1_153 ( .A(_70_), .Y(w_C_14_) );
INVX1 INVX1_154 ( .A(i_add2[14]), .Y(_71_) );
INVX1 INVX1_155 ( .A(i_add1[14]), .Y(_72_) );
NOR2X1 NOR2X1_89 ( .A(_71_), .B(_72_), .Y(_73_) );
INVX1 INVX1_156 ( .A(_73_), .Y(_74_) );
NOR2X1 NOR2X1_90 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_75_) );
INVX1 INVX1_157 ( .A(_75_), .Y(_76_) );
NOR2X1 NOR2X1_91 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_77_) );
INVX1 INVX1_158 ( .A(_77_), .Y(_78_) );
NAND3X1 NAND3X1_90 ( .A(_76_), .B(_78_), .C(_69_), .Y(_79_) );
AND2X2 AND2X2_75 ( .A(_79_), .B(_74_), .Y(_80_) );
INVX1 INVX1_159 ( .A(_80_), .Y(w_C_15_) );
AND2X2 AND2X2_76 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_81_) );
INVX1 INVX1_160 ( .A(_81_), .Y(_82_) );
NAND3X1 NAND3X1_91 ( .A(_74_), .B(_82_), .C(_79_), .Y(_83_) );
OAI21X1 OAI21X1_76 ( .A(i_add2[15]), .B(i_add1[15]), .C(_83_), .Y(_84_) );
INVX1 INVX1_161 ( .A(_84_), .Y(w_C_16_) );
INVX1 INVX1_162 ( .A(i_add2[16]), .Y(_85_) );
INVX1 INVX1_163 ( .A(i_add1[16]), .Y(_86_) );
NOR2X1 NOR2X1_92 ( .A(_85_), .B(_86_), .Y(_87_) );
INVX1 INVX1_164 ( .A(_87_), .Y(_88_) );
NOR2X1 NOR2X1_93 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_89_) );
INVX1 INVX1_165 ( .A(_89_), .Y(_90_) );
NOR2X1 NOR2X1_94 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_91_) );
INVX1 INVX1_166 ( .A(_91_), .Y(_92_) );
NAND3X1 NAND3X1_92 ( .A(_90_), .B(_92_), .C(_83_), .Y(_93_) );
AND2X2 AND2X2_77 ( .A(_93_), .B(_88_), .Y(_94_) );
INVX1 INVX1_167 ( .A(_94_), .Y(w_C_17_) );
AND2X2 AND2X2_78 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_95_) );
INVX1 INVX1_168 ( .A(_95_), .Y(_96_) );
NAND3X1 NAND3X1_93 ( .A(_88_), .B(_96_), .C(_93_), .Y(_97_) );
OAI21X1 OAI21X1_77 ( .A(i_add2[17]), .B(i_add1[17]), .C(_97_), .Y(_98_) );
INVX1 INVX1_169 ( .A(_98_), .Y(w_C_18_) );
INVX1 INVX1_170 ( .A(i_add2[18]), .Y(_99_) );
INVX1 INVX1_171 ( .A(i_add1[18]), .Y(_100_) );
NOR2X1 NOR2X1_95 ( .A(_99_), .B(_100_), .Y(_101_) );
INVX1 INVX1_172 ( .A(_101_), .Y(_102_) );
NOR2X1 NOR2X1_96 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_103_) );
INVX1 INVX1_173 ( .A(_103_), .Y(_104_) );
NOR2X1 NOR2X1_97 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_105_) );
INVX1 INVX1_174 ( .A(_105_), .Y(_106_) );
NAND3X1 NAND3X1_94 ( .A(_104_), .B(_106_), .C(_97_), .Y(_107_) );
AND2X2 AND2X2_79 ( .A(_107_), .B(_102_), .Y(_108_) );
INVX1 INVX1_175 ( .A(_108_), .Y(w_C_19_) );
AND2X2 AND2X2_80 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_109_) );
INVX1 INVX1_176 ( .A(_109_), .Y(_110_) );
NAND3X1 NAND3X1_95 ( .A(_102_), .B(_110_), .C(_107_), .Y(_111_) );
OAI21X1 OAI21X1_78 ( .A(i_add2[19]), .B(i_add1[19]), .C(_111_), .Y(_112_) );
INVX1 INVX1_177 ( .A(_112_), .Y(w_C_20_) );
INVX1 INVX1_178 ( .A(i_add2[20]), .Y(_113_) );
INVX1 INVX1_179 ( .A(i_add1[20]), .Y(_114_) );
NOR2X1 NOR2X1_98 ( .A(_113_), .B(_114_), .Y(_115_) );
INVX1 INVX1_180 ( .A(_115_), .Y(_116_) );
NOR2X1 NOR2X1_99 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_117_) );
INVX1 INVX1_181 ( .A(_117_), .Y(_118_) );
NOR2X1 NOR2X1_100 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_119_) );
INVX1 INVX1_182 ( .A(_119_), .Y(_120_) );
NAND3X1 NAND3X1_96 ( .A(_118_), .B(_120_), .C(_111_), .Y(_121_) );
AND2X2 AND2X2_81 ( .A(_121_), .B(_116_), .Y(_122_) );
INVX1 INVX1_183 ( .A(_122_), .Y(w_C_21_) );
AND2X2 AND2X2_82 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_123_) );
INVX1 INVX1_184 ( .A(_123_), .Y(_124_) );
NAND3X1 NAND3X1_97 ( .A(_116_), .B(_124_), .C(_121_), .Y(_125_) );
OAI21X1 OAI21X1_79 ( .A(i_add2[21]), .B(i_add1[21]), .C(_125_), .Y(_126_) );
INVX1 INVX1_185 ( .A(_126_), .Y(w_C_22_) );
INVX1 INVX1_186 ( .A(i_add2[22]), .Y(_127_) );
INVX1 INVX1_187 ( .A(i_add1[22]), .Y(_128_) );
NOR2X1 NOR2X1_101 ( .A(_127_), .B(_128_), .Y(_129_) );
INVX1 INVX1_188 ( .A(_129_), .Y(_130_) );
NOR2X1 NOR2X1_102 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_131_) );
INVX1 INVX1_189 ( .A(_131_), .Y(_132_) );
NOR2X1 NOR2X1_103 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_133_) );
INVX1 INVX1_190 ( .A(_133_), .Y(_134_) );
NAND3X1 NAND3X1_98 ( .A(_132_), .B(_134_), .C(_125_), .Y(_135_) );
AND2X2 AND2X2_83 ( .A(_135_), .B(_130_), .Y(_136_) );
INVX1 INVX1_191 ( .A(_136_), .Y(w_C_23_) );
AND2X2 AND2X2_84 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_137_) );
INVX1 INVX1_192 ( .A(_137_), .Y(_138_) );
NAND3X1 NAND3X1_99 ( .A(_130_), .B(_138_), .C(_135_), .Y(_139_) );
OAI21X1 OAI21X1_80 ( .A(i_add2[23]), .B(i_add1[23]), .C(_139_), .Y(_140_) );
INVX1 INVX1_193 ( .A(_140_), .Y(w_C_24_) );
INVX1 INVX1_194 ( .A(i_add2[24]), .Y(_141_) );
INVX1 INVX1_195 ( .A(i_add1[24]), .Y(_142_) );
NOR2X1 NOR2X1_104 ( .A(_141_), .B(_142_), .Y(_143_) );
INVX1 INVX1_196 ( .A(_143_), .Y(_144_) );
NOR2X1 NOR2X1_105 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_145_) );
INVX1 INVX1_197 ( .A(_145_), .Y(_146_) );
NOR2X1 NOR2X1_106 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_147_) );
INVX1 INVX1_198 ( .A(_147_), .Y(_148_) );
NAND3X1 NAND3X1_100 ( .A(_146_), .B(_148_), .C(_139_), .Y(_149_) );
AND2X2 AND2X2_85 ( .A(_149_), .B(_144_), .Y(_150_) );
INVX1 INVX1_199 ( .A(_150_), .Y(w_C_25_) );
AND2X2 AND2X2_86 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_151_) );
INVX1 INVX1_200 ( .A(_151_), .Y(_152_) );
NAND3X1 NAND3X1_101 ( .A(_144_), .B(_152_), .C(_149_), .Y(_153_) );
OAI21X1 OAI21X1_81 ( .A(i_add2[25]), .B(i_add1[25]), .C(_153_), .Y(_154_) );
INVX1 INVX1_201 ( .A(_154_), .Y(w_C_26_) );
INVX1 INVX1_202 ( .A(i_add2[26]), .Y(_155_) );
INVX1 INVX1_203 ( .A(i_add1[26]), .Y(_156_) );
NOR2X1 NOR2X1_107 ( .A(_155_), .B(_156_), .Y(_157_) );
INVX1 INVX1_204 ( .A(_157_), .Y(_158_) );
NOR2X1 NOR2X1_108 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_159_) );
INVX1 INVX1_205 ( .A(_159_), .Y(_160_) );
NOR2X1 NOR2X1_109 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_161_) );
BUFX2 BUFX2_53 ( .A(w_C_51_), .Y(_306__51_) );
BUFX2 BUFX2_54 ( .A(gnd), .Y(w_C_0_) );
endmodule
