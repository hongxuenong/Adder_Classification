module CSkipA_61bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [60:0] i_add_term1;
input [60:0] i_add_term2;
output [60:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

NOR2X1 NOR2X1_1 ( .A(_230_), .B(_235_), .Y(_36_) );
INVX1 INVX1_1 ( .A(_34_), .Y(_236_) );
NAND2X1 NAND2X1_1 ( .A(gnd), .B(_36_), .Y(_237_) );
OAI21X1 OAI21X1_1 ( .A(_36_), .B(_236_), .C(_237_), .Y(w_cout_12_) );
INVX1 INVX1_2 ( .A(i_add_term1[48]), .Y(_238_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[48]), .B(_238_), .Y(_239_) );
INVX1 INVX1_3 ( .A(i_add_term2[48]), .Y(_240_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term1[48]), .B(_240_), .Y(_241_) );
INVX1 INVX1_4 ( .A(i_add_term1[49]), .Y(_242_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[49]), .B(_242_), .Y(_243_) );
INVX1 INVX1_5 ( .A(i_add_term2[49]), .Y(_244_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term1[49]), .B(_244_), .Y(_245_) );
OAI22X1 OAI22X1_1 ( .A(_239_), .B(_241_), .C(_243_), .D(_245_), .Y(_246_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_247_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_248_) );
NOR2X1 NOR2X1_7 ( .A(_247_), .B(_248_), .Y(_249_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_250_) );
NAND2X1 NAND2X1_2 ( .A(_249_), .B(_250_), .Y(_251_) );
NOR2X1 NOR2X1_8 ( .A(_246_), .B(_251_), .Y(_39_) );
INVX1 INVX1_6 ( .A(_37_), .Y(_252_) );
NAND2X1 NAND2X1_3 ( .A(gnd), .B(_39_), .Y(_253_) );
OAI21X1 OAI21X1_2 ( .A(_39_), .B(_252_), .C(_253_), .Y(w_cout_13_) );
INVX1 INVX1_7 ( .A(i_add_term1[52]), .Y(_254_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[52]), .B(_254_), .Y(_255_) );
INVX1 INVX1_8 ( .A(i_add_term2[52]), .Y(_256_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term1[52]), .B(_256_), .Y(_257_) );
INVX1 INVX1_9 ( .A(i_add_term1[53]), .Y(_258_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[53]), .B(_258_), .Y(_259_) );
INVX1 INVX1_10 ( .A(i_add_term2[53]), .Y(_260_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term1[53]), .B(_260_), .Y(_261_) );
OAI22X1 OAI22X1_2 ( .A(_255_), .B(_257_), .C(_259_), .D(_261_), .Y(_262_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_263_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_264_) );
NOR2X1 NOR2X1_14 ( .A(_263_), .B(_264_), .Y(_265_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_266_) );
NAND2X1 NAND2X1_4 ( .A(_265_), .B(_266_), .Y(_267_) );
NOR2X1 NOR2X1_15 ( .A(_262_), .B(_267_), .Y(_42_) );
INVX1 INVX1_11 ( .A(_40_), .Y(_268_) );
NAND2X1 NAND2X1_5 ( .A(gnd), .B(_42_), .Y(_269_) );
OAI21X1 OAI21X1_3 ( .A(_42_), .B(_268_), .C(_269_), .Y(w_cout_14_) );
INVX1 INVX1_12 ( .A(i_add_term1[56]), .Y(_270_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[56]), .B(_270_), .Y(_271_) );
INVX1 INVX1_13 ( .A(i_add_term2[56]), .Y(_272_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term1[56]), .B(_272_), .Y(_273_) );
INVX1 INVX1_14 ( .A(i_add_term1[57]), .Y(_274_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[57]), .B(_274_), .Y(_275_) );
INVX1 INVX1_15 ( .A(i_add_term2[57]), .Y(_276_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term1[57]), .B(_276_), .Y(_277_) );
OAI22X1 OAI22X1_3 ( .A(_271_), .B(_273_), .C(_275_), .D(_277_), .Y(_278_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_279_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_280_) );
NOR2X1 NOR2X1_21 ( .A(_279_), .B(_280_), .Y(_281_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_282_) );
NAND2X1 NAND2X1_6 ( .A(_281_), .B(_282_), .Y(_283_) );
NOR2X1 NOR2X1_22 ( .A(_278_), .B(_283_), .Y(_45_) );
INVX1 INVX1_16 ( .A(_43_), .Y(_284_) );
NAND2X1 NAND2X1_7 ( .A(gnd), .B(_45_), .Y(_285_) );
OAI21X1 OAI21X1_4 ( .A(_45_), .B(_284_), .C(_285_), .Y(cskip1_inst_cin) );
INVX1 INVX1_17 ( .A(gnd), .Y(_289_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_290_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_291_) );
NAND3X1 NAND3X1_1 ( .A(_289_), .B(_291_), .C(_290_), .Y(_292_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_286_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_287_) );
OAI21X1 OAI21X1_5 ( .A(_286_), .B(_287_), .C(gnd), .Y(_288_) );
NAND2X1 NAND2X1_9 ( .A(_288_), .B(_292_), .Y(_0__0_) );
OAI21X1 OAI21X1_6 ( .A(_289_), .B(_286_), .C(_291_), .Y(_2__1_) );
INVX1 INVX1_18 ( .A(_2__1_), .Y(_296_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_297_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_298_) );
NAND3X1 NAND3X1_2 ( .A(_296_), .B(_298_), .C(_297_), .Y(_299_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_293_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_294_) );
OAI21X1 OAI21X1_7 ( .A(_293_), .B(_294_), .C(_2__1_), .Y(_295_) );
NAND2X1 NAND2X1_11 ( .A(_295_), .B(_299_), .Y(_0__1_) );
OAI21X1 OAI21X1_8 ( .A(_296_), .B(_293_), .C(_298_), .Y(_2__2_) );
INVX1 INVX1_19 ( .A(_2__2_), .Y(_303_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_304_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_305_) );
NAND3X1 NAND3X1_3 ( .A(_303_), .B(_305_), .C(_304_), .Y(_306_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_300_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_301_) );
OAI21X1 OAI21X1_9 ( .A(_300_), .B(_301_), .C(_2__2_), .Y(_302_) );
NAND2X1 NAND2X1_13 ( .A(_302_), .B(_306_), .Y(_0__2_) );
OAI21X1 OAI21X1_10 ( .A(_303_), .B(_300_), .C(_305_), .Y(_2__3_) );
INVX1 INVX1_20 ( .A(_2__3_), .Y(_310_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_311_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_312_) );
NAND3X1 NAND3X1_4 ( .A(_310_), .B(_312_), .C(_311_), .Y(_313_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_307_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_308_) );
OAI21X1 OAI21X1_11 ( .A(_307_), .B(_308_), .C(_2__3_), .Y(_309_) );
NAND2X1 NAND2X1_15 ( .A(_309_), .B(_313_), .Y(_0__3_) );
OAI21X1 OAI21X1_12 ( .A(_310_), .B(_307_), .C(_312_), .Y(_1_) );
INVX1 INVX1_21 ( .A(w_cout_1_), .Y(_317_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_318_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_319_) );
NAND3X1 NAND3X1_5 ( .A(_317_), .B(_319_), .C(_318_), .Y(_320_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_314_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_315_) );
OAI21X1 OAI21X1_13 ( .A(_314_), .B(_315_), .C(w_cout_1_), .Y(_316_) );
NAND2X1 NAND2X1_17 ( .A(_316_), .B(_320_), .Y(_0__4_) );
OAI21X1 OAI21X1_14 ( .A(_317_), .B(_314_), .C(_319_), .Y(_5__1_) );
INVX1 INVX1_22 ( .A(_5__1_), .Y(_324_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_325_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_326_) );
NAND3X1 NAND3X1_6 ( .A(_324_), .B(_326_), .C(_325_), .Y(_327_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_321_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_322_) );
OAI21X1 OAI21X1_15 ( .A(_321_), .B(_322_), .C(_5__1_), .Y(_323_) );
NAND2X1 NAND2X1_19 ( .A(_323_), .B(_327_), .Y(_0__5_) );
OAI21X1 OAI21X1_16 ( .A(_324_), .B(_321_), .C(_326_), .Y(_5__2_) );
INVX1 INVX1_23 ( .A(_5__2_), .Y(_331_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_332_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_333_) );
NAND3X1 NAND3X1_7 ( .A(_331_), .B(_333_), .C(_332_), .Y(_334_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_328_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_329_) );
OAI21X1 OAI21X1_17 ( .A(_328_), .B(_329_), .C(_5__2_), .Y(_330_) );
NAND2X1 NAND2X1_21 ( .A(_330_), .B(_334_), .Y(_0__6_) );
OAI21X1 OAI21X1_18 ( .A(_331_), .B(_328_), .C(_333_), .Y(_5__3_) );
INVX1 INVX1_24 ( .A(_5__3_), .Y(_338_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_339_) );
NAND2X1 NAND2X1_22 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_340_) );
NAND3X1 NAND3X1_8 ( .A(_338_), .B(_340_), .C(_339_), .Y(_341_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_335_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_336_) );
OAI21X1 OAI21X1_19 ( .A(_335_), .B(_336_), .C(_5__3_), .Y(_337_) );
NAND2X1 NAND2X1_23 ( .A(_337_), .B(_341_), .Y(_0__7_) );
OAI21X1 OAI21X1_20 ( .A(_338_), .B(_335_), .C(_340_), .Y(_4_) );
INVX1 INVX1_25 ( .A(w_cout_2_), .Y(_345_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_346_) );
NAND2X1 NAND2X1_24 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_347_) );
NAND3X1 NAND3X1_9 ( .A(_345_), .B(_347_), .C(_346_), .Y(_348_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_342_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_343_) );
OAI21X1 OAI21X1_21 ( .A(_342_), .B(_343_), .C(w_cout_2_), .Y(_344_) );
NAND2X1 NAND2X1_25 ( .A(_344_), .B(_348_), .Y(_0__8_) );
OAI21X1 OAI21X1_22 ( .A(_345_), .B(_342_), .C(_347_), .Y(_8__1_) );
INVX1 INVX1_26 ( .A(_8__1_), .Y(_352_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_353_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_354_) );
NAND3X1 NAND3X1_10 ( .A(_352_), .B(_354_), .C(_353_), .Y(_355_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_349_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_350_) );
OAI21X1 OAI21X1_23 ( .A(_349_), .B(_350_), .C(_8__1_), .Y(_351_) );
NAND2X1 NAND2X1_27 ( .A(_351_), .B(_355_), .Y(_0__9_) );
OAI21X1 OAI21X1_24 ( .A(_352_), .B(_349_), .C(_354_), .Y(_8__2_) );
INVX1 INVX1_27 ( .A(_8__2_), .Y(_359_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_360_) );
NAND2X1 NAND2X1_28 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_361_) );
NAND3X1 NAND3X1_11 ( .A(_359_), .B(_361_), .C(_360_), .Y(_362_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_356_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_357_) );
OAI21X1 OAI21X1_25 ( .A(_356_), .B(_357_), .C(_8__2_), .Y(_358_) );
NAND2X1 NAND2X1_29 ( .A(_358_), .B(_362_), .Y(_0__10_) );
OAI21X1 OAI21X1_26 ( .A(_359_), .B(_356_), .C(_361_), .Y(_8__3_) );
INVX1 INVX1_28 ( .A(_8__3_), .Y(_366_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_367_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_368_) );
NAND3X1 NAND3X1_12 ( .A(_366_), .B(_368_), .C(_367_), .Y(_369_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_363_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_364_) );
OAI21X1 OAI21X1_27 ( .A(_363_), .B(_364_), .C(_8__3_), .Y(_365_) );
NAND2X1 NAND2X1_31 ( .A(_365_), .B(_369_), .Y(_0__11_) );
OAI21X1 OAI21X1_28 ( .A(_366_), .B(_363_), .C(_368_), .Y(_7_) );
INVX1 INVX1_29 ( .A(w_cout_3_), .Y(_373_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_374_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_375_) );
NAND3X1 NAND3X1_13 ( .A(_373_), .B(_375_), .C(_374_), .Y(_376_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_370_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_371_) );
OAI21X1 OAI21X1_29 ( .A(_370_), .B(_371_), .C(w_cout_3_), .Y(_372_) );
NAND2X1 NAND2X1_33 ( .A(_372_), .B(_376_), .Y(_0__12_) );
OAI21X1 OAI21X1_30 ( .A(_373_), .B(_370_), .C(_375_), .Y(_11__1_) );
INVX1 INVX1_30 ( .A(_11__1_), .Y(_380_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_381_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_382_) );
NAND3X1 NAND3X1_14 ( .A(_380_), .B(_382_), .C(_381_), .Y(_383_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_377_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_378_) );
OAI21X1 OAI21X1_31 ( .A(_377_), .B(_378_), .C(_11__1_), .Y(_379_) );
NAND2X1 NAND2X1_35 ( .A(_379_), .B(_383_), .Y(_0__13_) );
OAI21X1 OAI21X1_32 ( .A(_380_), .B(_377_), .C(_382_), .Y(_11__2_) );
INVX1 INVX1_31 ( .A(_11__2_), .Y(_387_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_388_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_389_) );
NAND3X1 NAND3X1_15 ( .A(_387_), .B(_389_), .C(_388_), .Y(_390_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_384_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_385_) );
OAI21X1 OAI21X1_33 ( .A(_384_), .B(_385_), .C(_11__2_), .Y(_386_) );
NAND2X1 NAND2X1_37 ( .A(_386_), .B(_390_), .Y(_0__14_) );
OAI21X1 OAI21X1_34 ( .A(_387_), .B(_384_), .C(_389_), .Y(_11__3_) );
INVX1 INVX1_32 ( .A(_11__3_), .Y(_394_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_395_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_396_) );
NAND3X1 NAND3X1_16 ( .A(_394_), .B(_396_), .C(_395_), .Y(_397_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_391_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_392_) );
OAI21X1 OAI21X1_35 ( .A(_391_), .B(_392_), .C(_11__3_), .Y(_393_) );
NAND2X1 NAND2X1_39 ( .A(_393_), .B(_397_), .Y(_0__15_) );
OAI21X1 OAI21X1_36 ( .A(_394_), .B(_391_), .C(_396_), .Y(_10_) );
INVX1 INVX1_33 ( .A(w_cout_4_), .Y(_401_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_402_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_403_) );
NAND3X1 NAND3X1_17 ( .A(_401_), .B(_403_), .C(_402_), .Y(_404_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_398_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_399_) );
OAI21X1 OAI21X1_37 ( .A(_398_), .B(_399_), .C(w_cout_4_), .Y(_400_) );
NAND2X1 NAND2X1_41 ( .A(_400_), .B(_404_), .Y(_0__16_) );
OAI21X1 OAI21X1_38 ( .A(_401_), .B(_398_), .C(_403_), .Y(_14__1_) );
INVX1 INVX1_34 ( .A(_14__1_), .Y(_408_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_409_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_410_) );
NAND3X1 NAND3X1_18 ( .A(_408_), .B(_410_), .C(_409_), .Y(_411_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_405_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_406_) );
OAI21X1 OAI21X1_39 ( .A(_405_), .B(_406_), .C(_14__1_), .Y(_407_) );
NAND2X1 NAND2X1_43 ( .A(_407_), .B(_411_), .Y(_0__17_) );
OAI21X1 OAI21X1_40 ( .A(_408_), .B(_405_), .C(_410_), .Y(_14__2_) );
INVX1 INVX1_35 ( .A(_14__2_), .Y(_415_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_416_) );
NAND2X1 NAND2X1_44 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_417_) );
NAND3X1 NAND3X1_19 ( .A(_415_), .B(_417_), .C(_416_), .Y(_418_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_412_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_413_) );
OAI21X1 OAI21X1_41 ( .A(_412_), .B(_413_), .C(_14__2_), .Y(_414_) );
NAND2X1 NAND2X1_45 ( .A(_414_), .B(_418_), .Y(_0__18_) );
OAI21X1 OAI21X1_42 ( .A(_415_), .B(_412_), .C(_417_), .Y(_14__3_) );
INVX1 INVX1_36 ( .A(_14__3_), .Y(_422_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_423_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_424_) );
NAND3X1 NAND3X1_20 ( .A(_422_), .B(_424_), .C(_423_), .Y(_425_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_419_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_420_) );
OAI21X1 OAI21X1_43 ( .A(_419_), .B(_420_), .C(_14__3_), .Y(_421_) );
NAND2X1 NAND2X1_47 ( .A(_421_), .B(_425_), .Y(_0__19_) );
OAI21X1 OAI21X1_44 ( .A(_422_), .B(_419_), .C(_424_), .Y(_13_) );
INVX1 INVX1_37 ( .A(w_cout_5_), .Y(_429_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_430_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_431_) );
NAND3X1 NAND3X1_21 ( .A(_429_), .B(_431_), .C(_430_), .Y(_432_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_426_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_427_) );
OAI21X1 OAI21X1_45 ( .A(_426_), .B(_427_), .C(w_cout_5_), .Y(_428_) );
NAND2X1 NAND2X1_49 ( .A(_428_), .B(_432_), .Y(_0__20_) );
OAI21X1 OAI21X1_46 ( .A(_429_), .B(_426_), .C(_431_), .Y(_17__1_) );
INVX1 INVX1_38 ( .A(_17__1_), .Y(_436_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_437_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_438_) );
NAND3X1 NAND3X1_22 ( .A(_436_), .B(_438_), .C(_437_), .Y(_439_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_433_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_434_) );
OAI21X1 OAI21X1_47 ( .A(_433_), .B(_434_), .C(_17__1_), .Y(_435_) );
NAND2X1 NAND2X1_51 ( .A(_435_), .B(_439_), .Y(_0__21_) );
OAI21X1 OAI21X1_48 ( .A(_436_), .B(_433_), .C(_438_), .Y(_17__2_) );
INVX1 INVX1_39 ( .A(_17__2_), .Y(_443_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_444_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_445_) );
NAND3X1 NAND3X1_23 ( .A(_443_), .B(_445_), .C(_444_), .Y(_446_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_440_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_441_) );
OAI21X1 OAI21X1_49 ( .A(_440_), .B(_441_), .C(_17__2_), .Y(_442_) );
NAND2X1 NAND2X1_53 ( .A(_442_), .B(_446_), .Y(_0__22_) );
OAI21X1 OAI21X1_50 ( .A(_443_), .B(_440_), .C(_445_), .Y(_17__3_) );
INVX1 INVX1_40 ( .A(_17__3_), .Y(_450_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_451_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_452_) );
NAND3X1 NAND3X1_24 ( .A(_450_), .B(_452_), .C(_451_), .Y(_453_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_447_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_448_) );
OAI21X1 OAI21X1_51 ( .A(_447_), .B(_448_), .C(_17__3_), .Y(_449_) );
NAND2X1 NAND2X1_55 ( .A(_449_), .B(_453_), .Y(_0__23_) );
OAI21X1 OAI21X1_52 ( .A(_450_), .B(_447_), .C(_452_), .Y(_16_) );
INVX1 INVX1_41 ( .A(w_cout_6_), .Y(_457_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_458_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_459_) );
NAND3X1 NAND3X1_25 ( .A(_457_), .B(_459_), .C(_458_), .Y(_460_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_454_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_455_) );
OAI21X1 OAI21X1_53 ( .A(_454_), .B(_455_), .C(w_cout_6_), .Y(_456_) );
NAND2X1 NAND2X1_57 ( .A(_456_), .B(_460_), .Y(_0__24_) );
OAI21X1 OAI21X1_54 ( .A(_457_), .B(_454_), .C(_459_), .Y(_20__1_) );
INVX1 INVX1_42 ( .A(_20__1_), .Y(_464_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_465_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_466_) );
NAND3X1 NAND3X1_26 ( .A(_464_), .B(_466_), .C(_465_), .Y(_467_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_461_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_462_) );
OAI21X1 OAI21X1_55 ( .A(_461_), .B(_462_), .C(_20__1_), .Y(_463_) );
NAND2X1 NAND2X1_59 ( .A(_463_), .B(_467_), .Y(_0__25_) );
OAI21X1 OAI21X1_56 ( .A(_464_), .B(_461_), .C(_466_), .Y(_20__2_) );
INVX1 INVX1_43 ( .A(_20__2_), .Y(_471_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_472_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_473_) );
NAND3X1 NAND3X1_27 ( .A(_471_), .B(_473_), .C(_472_), .Y(_474_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_468_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_469_) );
OAI21X1 OAI21X1_57 ( .A(_468_), .B(_469_), .C(_20__2_), .Y(_470_) );
NAND2X1 NAND2X1_61 ( .A(_470_), .B(_474_), .Y(_0__26_) );
OAI21X1 OAI21X1_58 ( .A(_471_), .B(_468_), .C(_473_), .Y(_20__3_) );
INVX1 INVX1_44 ( .A(_20__3_), .Y(_478_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_479_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_480_) );
NAND3X1 NAND3X1_28 ( .A(_478_), .B(_480_), .C(_479_), .Y(_481_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_475_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_476_) );
OAI21X1 OAI21X1_59 ( .A(_475_), .B(_476_), .C(_20__3_), .Y(_477_) );
NAND2X1 NAND2X1_63 ( .A(_477_), .B(_481_), .Y(_0__27_) );
OAI21X1 OAI21X1_60 ( .A(_478_), .B(_475_), .C(_480_), .Y(_19_) );
INVX1 INVX1_45 ( .A(w_cout_7_), .Y(_485_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_486_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_487_) );
NAND3X1 NAND3X1_29 ( .A(_485_), .B(_487_), .C(_486_), .Y(_488_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_482_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_483_) );
OAI21X1 OAI21X1_61 ( .A(_482_), .B(_483_), .C(w_cout_7_), .Y(_484_) );
NAND2X1 NAND2X1_65 ( .A(_484_), .B(_488_), .Y(_0__28_) );
OAI21X1 OAI21X1_62 ( .A(_485_), .B(_482_), .C(_487_), .Y(_23__1_) );
INVX1 INVX1_46 ( .A(_23__1_), .Y(_492_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_493_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_494_) );
NAND3X1 NAND3X1_30 ( .A(_492_), .B(_494_), .C(_493_), .Y(_495_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_489_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_490_) );
OAI21X1 OAI21X1_63 ( .A(_489_), .B(_490_), .C(_23__1_), .Y(_491_) );
NAND2X1 NAND2X1_67 ( .A(_491_), .B(_495_), .Y(_0__29_) );
OAI21X1 OAI21X1_64 ( .A(_492_), .B(_489_), .C(_494_), .Y(_23__2_) );
INVX1 INVX1_47 ( .A(_23__2_), .Y(_499_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_500_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_501_) );
NAND3X1 NAND3X1_31 ( .A(_499_), .B(_501_), .C(_500_), .Y(_502_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_496_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_497_) );
OAI21X1 OAI21X1_65 ( .A(_496_), .B(_497_), .C(_23__2_), .Y(_498_) );
NAND2X1 NAND2X1_69 ( .A(_498_), .B(_502_), .Y(_0__30_) );
OAI21X1 OAI21X1_66 ( .A(_499_), .B(_496_), .C(_501_), .Y(_23__3_) );
INVX1 INVX1_48 ( .A(_23__3_), .Y(_506_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_507_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_508_) );
NAND3X1 NAND3X1_32 ( .A(_506_), .B(_508_), .C(_507_), .Y(_509_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_503_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_504_) );
OAI21X1 OAI21X1_67 ( .A(_503_), .B(_504_), .C(_23__3_), .Y(_505_) );
NAND2X1 NAND2X1_71 ( .A(_505_), .B(_509_), .Y(_0__31_) );
OAI21X1 OAI21X1_68 ( .A(_506_), .B(_503_), .C(_508_), .Y(_22_) );
INVX1 INVX1_49 ( .A(w_cout_8_), .Y(_513_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_514_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_515_) );
NAND3X1 NAND3X1_33 ( .A(_513_), .B(_515_), .C(_514_), .Y(_516_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_510_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_511_) );
OAI21X1 OAI21X1_69 ( .A(_510_), .B(_511_), .C(w_cout_8_), .Y(_512_) );
NAND2X1 NAND2X1_73 ( .A(_512_), .B(_516_), .Y(_0__32_) );
OAI21X1 OAI21X1_70 ( .A(_513_), .B(_510_), .C(_515_), .Y(_26__1_) );
INVX1 INVX1_50 ( .A(_26__1_), .Y(_520_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_521_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_522_) );
NAND3X1 NAND3X1_34 ( .A(_520_), .B(_522_), .C(_521_), .Y(_523_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_517_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_518_) );
OAI21X1 OAI21X1_71 ( .A(_517_), .B(_518_), .C(_26__1_), .Y(_519_) );
NAND2X1 NAND2X1_75 ( .A(_519_), .B(_523_), .Y(_0__33_) );
OAI21X1 OAI21X1_72 ( .A(_520_), .B(_517_), .C(_522_), .Y(_26__2_) );
INVX1 INVX1_51 ( .A(_26__2_), .Y(_527_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_528_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_529_) );
NAND3X1 NAND3X1_35 ( .A(_527_), .B(_529_), .C(_528_), .Y(_530_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_524_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_525_) );
OAI21X1 OAI21X1_73 ( .A(_524_), .B(_525_), .C(_26__2_), .Y(_526_) );
NAND2X1 NAND2X1_77 ( .A(_526_), .B(_530_), .Y(_0__34_) );
OAI21X1 OAI21X1_74 ( .A(_527_), .B(_524_), .C(_529_), .Y(_26__3_) );
INVX1 INVX1_52 ( .A(_26__3_), .Y(_534_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_535_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_536_) );
NAND3X1 NAND3X1_36 ( .A(_534_), .B(_536_), .C(_535_), .Y(_537_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_531_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_532_) );
OAI21X1 OAI21X1_75 ( .A(_531_), .B(_532_), .C(_26__3_), .Y(_533_) );
NAND2X1 NAND2X1_79 ( .A(_533_), .B(_537_), .Y(_0__35_) );
OAI21X1 OAI21X1_76 ( .A(_534_), .B(_531_), .C(_536_), .Y(_25_) );
INVX1 INVX1_53 ( .A(w_cout_9_), .Y(_541_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_542_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_543_) );
NAND3X1 NAND3X1_37 ( .A(_541_), .B(_543_), .C(_542_), .Y(_544_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_538_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_539_) );
OAI21X1 OAI21X1_77 ( .A(_538_), .B(_539_), .C(w_cout_9_), .Y(_540_) );
NAND2X1 NAND2X1_81 ( .A(_540_), .B(_544_), .Y(_0__36_) );
OAI21X1 OAI21X1_78 ( .A(_541_), .B(_538_), .C(_543_), .Y(_29__1_) );
INVX1 INVX1_54 ( .A(_29__1_), .Y(_548_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_549_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_550_) );
NAND3X1 NAND3X1_38 ( .A(_548_), .B(_550_), .C(_549_), .Y(_551_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_545_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_546_) );
OAI21X1 OAI21X1_79 ( .A(_545_), .B(_546_), .C(_29__1_), .Y(_547_) );
NAND2X1 NAND2X1_83 ( .A(_547_), .B(_551_), .Y(_0__37_) );
OAI21X1 OAI21X1_80 ( .A(_548_), .B(_545_), .C(_550_), .Y(_29__2_) );
INVX1 INVX1_55 ( .A(_29__2_), .Y(_555_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_556_) );
NAND2X1 NAND2X1_84 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_557_) );
NAND3X1 NAND3X1_39 ( .A(_555_), .B(_557_), .C(_556_), .Y(_558_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_552_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_553_) );
OAI21X1 OAI21X1_81 ( .A(_552_), .B(_553_), .C(_29__2_), .Y(_554_) );
NAND2X1 NAND2X1_85 ( .A(_554_), .B(_558_), .Y(_0__38_) );
OAI21X1 OAI21X1_82 ( .A(_555_), .B(_552_), .C(_557_), .Y(_29__3_) );
INVX1 INVX1_56 ( .A(_29__3_), .Y(_562_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_563_) );
NAND2X1 NAND2X1_86 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_564_) );
NAND3X1 NAND3X1_40 ( .A(_562_), .B(_564_), .C(_563_), .Y(_565_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_559_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_560_) );
OAI21X1 OAI21X1_83 ( .A(_559_), .B(_560_), .C(_29__3_), .Y(_561_) );
NAND2X1 NAND2X1_87 ( .A(_561_), .B(_565_), .Y(_0__39_) );
OAI21X1 OAI21X1_84 ( .A(_562_), .B(_559_), .C(_564_), .Y(_28_) );
INVX1 INVX1_57 ( .A(w_cout_10_), .Y(_569_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_570_) );
NAND2X1 NAND2X1_88 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_571_) );
NAND3X1 NAND3X1_41 ( .A(_569_), .B(_571_), .C(_570_), .Y(_572_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_566_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_567_) );
OAI21X1 OAI21X1_85 ( .A(_566_), .B(_567_), .C(w_cout_10_), .Y(_568_) );
NAND2X1 NAND2X1_89 ( .A(_568_), .B(_572_), .Y(_0__40_) );
OAI21X1 OAI21X1_86 ( .A(_569_), .B(_566_), .C(_571_), .Y(_32__1_) );
INVX1 INVX1_58 ( .A(_32__1_), .Y(_576_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_577_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_578_) );
NAND3X1 NAND3X1_42 ( .A(_576_), .B(_578_), .C(_577_), .Y(_579_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_573_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_574_) );
OAI21X1 OAI21X1_87 ( .A(_573_), .B(_574_), .C(_32__1_), .Y(_575_) );
NAND2X1 NAND2X1_91 ( .A(_575_), .B(_579_), .Y(_0__41_) );
OAI21X1 OAI21X1_88 ( .A(_576_), .B(_573_), .C(_578_), .Y(_32__2_) );
INVX1 INVX1_59 ( .A(_32__2_), .Y(_583_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_584_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_585_) );
NAND3X1 NAND3X1_43 ( .A(_583_), .B(_585_), .C(_584_), .Y(_586_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_580_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_581_) );
OAI21X1 OAI21X1_89 ( .A(_580_), .B(_581_), .C(_32__2_), .Y(_582_) );
NAND2X1 NAND2X1_93 ( .A(_582_), .B(_586_), .Y(_0__42_) );
OAI21X1 OAI21X1_90 ( .A(_583_), .B(_580_), .C(_585_), .Y(_32__3_) );
INVX1 INVX1_60 ( .A(_32__3_), .Y(_590_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_591_) );
NAND2X1 NAND2X1_94 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_592_) );
NAND3X1 NAND3X1_44 ( .A(_590_), .B(_592_), .C(_591_), .Y(_593_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_587_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_588_) );
OAI21X1 OAI21X1_91 ( .A(_587_), .B(_588_), .C(_32__3_), .Y(_589_) );
NAND2X1 NAND2X1_95 ( .A(_589_), .B(_593_), .Y(_0__43_) );
OAI21X1 OAI21X1_92 ( .A(_590_), .B(_587_), .C(_592_), .Y(_31_) );
INVX1 INVX1_61 ( .A(w_cout_11_), .Y(_597_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_598_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_599_) );
NAND3X1 NAND3X1_45 ( .A(_597_), .B(_599_), .C(_598_), .Y(_600_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_594_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_595_) );
OAI21X1 OAI21X1_93 ( .A(_594_), .B(_595_), .C(w_cout_11_), .Y(_596_) );
NAND2X1 NAND2X1_97 ( .A(_596_), .B(_600_), .Y(_0__44_) );
OAI21X1 OAI21X1_94 ( .A(_597_), .B(_594_), .C(_599_), .Y(_35__1_) );
INVX1 INVX1_62 ( .A(_35__1_), .Y(_604_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_605_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_606_) );
NAND3X1 NAND3X1_46 ( .A(_604_), .B(_606_), .C(_605_), .Y(_607_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_601_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_602_) );
OAI21X1 OAI21X1_95 ( .A(_601_), .B(_602_), .C(_35__1_), .Y(_603_) );
NAND2X1 NAND2X1_99 ( .A(_603_), .B(_607_), .Y(_0__45_) );
OAI21X1 OAI21X1_96 ( .A(_604_), .B(_601_), .C(_606_), .Y(_35__2_) );
INVX1 INVX1_63 ( .A(_35__2_), .Y(_611_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_612_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_613_) );
NAND3X1 NAND3X1_47 ( .A(_611_), .B(_613_), .C(_612_), .Y(_614_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_608_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_609_) );
OAI21X1 OAI21X1_97 ( .A(_608_), .B(_609_), .C(_35__2_), .Y(_610_) );
NAND2X1 NAND2X1_101 ( .A(_610_), .B(_614_), .Y(_0__46_) );
OAI21X1 OAI21X1_98 ( .A(_611_), .B(_608_), .C(_613_), .Y(_35__3_) );
INVX1 INVX1_64 ( .A(_35__3_), .Y(_618_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_619_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_620_) );
NAND3X1 NAND3X1_48 ( .A(_618_), .B(_620_), .C(_619_), .Y(_621_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_615_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_616_) );
OAI21X1 OAI21X1_99 ( .A(_615_), .B(_616_), .C(_35__3_), .Y(_617_) );
NAND2X1 NAND2X1_103 ( .A(_617_), .B(_621_), .Y(_0__47_) );
OAI21X1 OAI21X1_100 ( .A(_618_), .B(_615_), .C(_620_), .Y(_34_) );
INVX1 INVX1_65 ( .A(w_cout_12_), .Y(_625_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_626_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_627_) );
NAND3X1 NAND3X1_49 ( .A(_625_), .B(_627_), .C(_626_), .Y(_628_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_622_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_623_) );
OAI21X1 OAI21X1_101 ( .A(_622_), .B(_623_), .C(w_cout_12_), .Y(_624_) );
NAND2X1 NAND2X1_105 ( .A(_624_), .B(_628_), .Y(_0__48_) );
OAI21X1 OAI21X1_102 ( .A(_625_), .B(_622_), .C(_627_), .Y(_38__1_) );
INVX1 INVX1_66 ( .A(_38__1_), .Y(_632_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_633_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_634_) );
NAND3X1 NAND3X1_50 ( .A(_632_), .B(_634_), .C(_633_), .Y(_635_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_629_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_630_) );
OAI21X1 OAI21X1_103 ( .A(_629_), .B(_630_), .C(_38__1_), .Y(_631_) );
NAND2X1 NAND2X1_107 ( .A(_631_), .B(_635_), .Y(_0__49_) );
OAI21X1 OAI21X1_104 ( .A(_632_), .B(_629_), .C(_634_), .Y(_38__2_) );
INVX1 INVX1_67 ( .A(_38__2_), .Y(_639_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_640_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_641_) );
NAND3X1 NAND3X1_51 ( .A(_639_), .B(_641_), .C(_640_), .Y(_642_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_636_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_637_) );
OAI21X1 OAI21X1_105 ( .A(_636_), .B(_637_), .C(_38__2_), .Y(_638_) );
NAND2X1 NAND2X1_109 ( .A(_638_), .B(_642_), .Y(_0__50_) );
OAI21X1 OAI21X1_106 ( .A(_639_), .B(_636_), .C(_641_), .Y(_38__3_) );
INVX1 INVX1_68 ( .A(_38__3_), .Y(_646_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_647_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_648_) );
NAND3X1 NAND3X1_52 ( .A(_646_), .B(_648_), .C(_647_), .Y(_649_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_643_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_644_) );
OAI21X1 OAI21X1_107 ( .A(_643_), .B(_644_), .C(_38__3_), .Y(_645_) );
NAND2X1 NAND2X1_111 ( .A(_645_), .B(_649_), .Y(_0__51_) );
OAI21X1 OAI21X1_108 ( .A(_646_), .B(_643_), .C(_648_), .Y(_37_) );
INVX1 INVX1_69 ( .A(w_cout_13_), .Y(_653_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_654_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_655_) );
NAND3X1 NAND3X1_53 ( .A(_653_), .B(_655_), .C(_654_), .Y(_656_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_650_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_651_) );
OAI21X1 OAI21X1_109 ( .A(_650_), .B(_651_), .C(w_cout_13_), .Y(_652_) );
NAND2X1 NAND2X1_113 ( .A(_652_), .B(_656_), .Y(_0__52_) );
OAI21X1 OAI21X1_110 ( .A(_653_), .B(_650_), .C(_655_), .Y(_41__1_) );
INVX1 INVX1_70 ( .A(_41__1_), .Y(_660_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_661_) );
NAND2X1 NAND2X1_114 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_662_) );
NAND3X1 NAND3X1_54 ( .A(_660_), .B(_662_), .C(_661_), .Y(_663_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_657_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_658_) );
OAI21X1 OAI21X1_111 ( .A(_657_), .B(_658_), .C(_41__1_), .Y(_659_) );
NAND2X1 NAND2X1_115 ( .A(_659_), .B(_663_), .Y(_0__53_) );
OAI21X1 OAI21X1_112 ( .A(_660_), .B(_657_), .C(_662_), .Y(_41__2_) );
INVX1 INVX1_71 ( .A(_41__2_), .Y(_667_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_668_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_669_) );
NAND3X1 NAND3X1_55 ( .A(_667_), .B(_669_), .C(_668_), .Y(_670_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_664_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_665_) );
OAI21X1 OAI21X1_113 ( .A(_664_), .B(_665_), .C(_41__2_), .Y(_666_) );
NAND2X1 NAND2X1_117 ( .A(_666_), .B(_670_), .Y(_0__54_) );
OAI21X1 OAI21X1_114 ( .A(_667_), .B(_664_), .C(_669_), .Y(_41__3_) );
INVX1 INVX1_72 ( .A(_41__3_), .Y(_674_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_675_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_676_) );
NAND3X1 NAND3X1_56 ( .A(_674_), .B(_676_), .C(_675_), .Y(_677_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_671_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_672_) );
OAI21X1 OAI21X1_115 ( .A(_671_), .B(_672_), .C(_41__3_), .Y(_673_) );
NAND2X1 NAND2X1_119 ( .A(_673_), .B(_677_), .Y(_0__55_) );
OAI21X1 OAI21X1_116 ( .A(_674_), .B(_671_), .C(_676_), .Y(_40_) );
INVX1 INVX1_73 ( .A(w_cout_14_), .Y(_681_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_682_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_683_) );
NAND3X1 NAND3X1_57 ( .A(_681_), .B(_683_), .C(_682_), .Y(_684_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_678_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_679_) );
OAI21X1 OAI21X1_117 ( .A(_678_), .B(_679_), .C(w_cout_14_), .Y(_680_) );
NAND2X1 NAND2X1_121 ( .A(_680_), .B(_684_), .Y(_0__56_) );
OAI21X1 OAI21X1_118 ( .A(_681_), .B(_678_), .C(_683_), .Y(_44__1_) );
INVX1 INVX1_74 ( .A(_44__1_), .Y(_688_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_689_) );
NAND2X1 NAND2X1_122 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_690_) );
NAND3X1 NAND3X1_58 ( .A(_688_), .B(_690_), .C(_689_), .Y(_691_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_685_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_686_) );
OAI21X1 OAI21X1_119 ( .A(_685_), .B(_686_), .C(_44__1_), .Y(_687_) );
NAND2X1 NAND2X1_123 ( .A(_687_), .B(_691_), .Y(_0__57_) );
OAI21X1 OAI21X1_120 ( .A(_688_), .B(_685_), .C(_690_), .Y(_44__2_) );
INVX1 INVX1_75 ( .A(_44__2_), .Y(_695_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_696_) );
NAND2X1 NAND2X1_124 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_697_) );
NAND3X1 NAND3X1_59 ( .A(_695_), .B(_697_), .C(_696_), .Y(_698_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_692_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_693_) );
OAI21X1 OAI21X1_121 ( .A(_692_), .B(_693_), .C(_44__2_), .Y(_694_) );
NAND2X1 NAND2X1_125 ( .A(_694_), .B(_698_), .Y(_0__58_) );
OAI21X1 OAI21X1_122 ( .A(_695_), .B(_692_), .C(_697_), .Y(_44__3_) );
INVX1 INVX1_76 ( .A(_44__3_), .Y(_702_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_703_) );
NAND2X1 NAND2X1_126 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_704_) );
NAND3X1 NAND3X1_60 ( .A(_702_), .B(_704_), .C(_703_), .Y(_705_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_699_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_700_) );
OAI21X1 OAI21X1_123 ( .A(_699_), .B(_700_), .C(_44__3_), .Y(_701_) );
NAND2X1 NAND2X1_127 ( .A(_701_), .B(_705_), .Y(_0__59_) );
OAI21X1 OAI21X1_124 ( .A(_702_), .B(_699_), .C(_704_), .Y(_43_) );
INVX1 INVX1_77 ( .A(cskip1_inst_cin), .Y(_709_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_710_) );
NAND2X1 NAND2X1_128 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_711_) );
NAND3X1 NAND3X1_61 ( .A(_709_), .B(_711_), .C(_710_), .Y(_712_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_706_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_707_) );
OAI21X1 OAI21X1_125 ( .A(_706_), .B(_707_), .C(cskip1_inst_cin), .Y(_708_) );
NAND2X1 NAND2X1_129 ( .A(_708_), .B(_712_), .Y(cskip1_inst_sum) );
OAI21X1 OAI21X1_126 ( .A(_709_), .B(_706_), .C(_711_), .Y(cskip1_inst_rca0_w_CARRY_1_) );
INVX1 INVX1_78 ( .A(cskip1_inst_rca0_w_CARRY_1_), .Y(_714_) );
NAND2X1 NAND2X1_130 ( .A(gnd), .B(gnd), .Y(_715_) );
NOR2X1 NOR2X1_84 ( .A(gnd), .B(gnd), .Y(_713_) );
OAI21X1 OAI21X1_127 ( .A(_714_), .B(_713_), .C(_715_), .Y(cskip1_inst_rca0_w_CARRY_2_) );
INVX1 INVX1_79 ( .A(cskip1_inst_rca0_w_CARRY_2_), .Y(_717_) );
NAND2X1 NAND2X1_131 ( .A(gnd), .B(gnd), .Y(_718_) );
NOR2X1 NOR2X1_85 ( .A(gnd), .B(gnd), .Y(_716_) );
OAI21X1 OAI21X1_128 ( .A(_717_), .B(_716_), .C(_718_), .Y(cskip1_inst_rca0_w_CARRY_3_) );
INVX1 INVX1_80 ( .A(cskip1_inst_rca0_w_CARRY_3_), .Y(_720_) );
NAND2X1 NAND2X1_132 ( .A(gnd), .B(gnd), .Y(_721_) );
NOR2X1 NOR2X1_86 ( .A(gnd), .B(gnd), .Y(_719_) );
OAI21X1 OAI21X1_129 ( .A(_720_), .B(_719_), .C(_721_), .Y(cskip1_inst_cout0) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_722_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_723_) );
NOR2X1 NOR2X1_88 ( .A(_722_), .B(_723_), .Y(cskip1_inst_skip0_P) );
INVX1 INVX1_81 ( .A(cskip1_inst_cout0), .Y(_724_) );
NAND2X1 NAND2X1_133 ( .A(gnd), .B(cskip1_inst_skip0_P), .Y(_725_) );
OAI21X1 OAI21X1_130 ( .A(cskip1_inst_skip0_P), .B(_724_), .C(_725_), .Y(w_cout_16_) );
BUFX2 BUFX2_1 ( .A(w_cout_16_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .A(_0__54_), .Y(sum[54]) );
BUFX2 BUFX2_57 ( .A(_0__55_), .Y(sum[55]) );
BUFX2 BUFX2_58 ( .A(_0__56_), .Y(sum[56]) );
BUFX2 BUFX2_59 ( .A(_0__57_), .Y(sum[57]) );
BUFX2 BUFX2_60 ( .A(_0__58_), .Y(sum[58]) );
BUFX2 BUFX2_61 ( .A(_0__59_), .Y(sum[59]) );
BUFX2 BUFX2_62 ( .A(cskip1_inst_sum), .Y(sum[60]) );
INVX1 INVX1_82 ( .A(i_add_term1[0]), .Y(_46_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[0]), .B(_46_), .Y(_47_) );
INVX1 INVX1_83 ( .A(i_add_term2[0]), .Y(_48_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term1[0]), .B(_48_), .Y(_49_) );
INVX1 INVX1_84 ( .A(i_add_term1[1]), .Y(_50_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[1]), .B(_50_), .Y(_51_) );
INVX1 INVX1_85 ( .A(i_add_term2[1]), .Y(_52_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term1[1]), .B(_52_), .Y(_53_) );
OAI22X1 OAI22X1_4 ( .A(_47_), .B(_49_), .C(_51_), .D(_53_), .Y(_54_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_55_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_56_) );
NOR2X1 NOR2X1_94 ( .A(_55_), .B(_56_), .Y(_57_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_58_) );
NAND2X1 NAND2X1_134 ( .A(_57_), .B(_58_), .Y(_59_) );
NOR2X1 NOR2X1_95 ( .A(_54_), .B(_59_), .Y(_3_) );
INVX1 INVX1_86 ( .A(_1_), .Y(_60_) );
NAND2X1 NAND2X1_135 ( .A(gnd), .B(_3_), .Y(_61_) );
OAI21X1 OAI21X1_131 ( .A(_3_), .B(_60_), .C(_61_), .Y(w_cout_1_) );
INVX1 INVX1_87 ( .A(i_add_term1[4]), .Y(_62_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[4]), .B(_62_), .Y(_63_) );
INVX1 INVX1_88 ( .A(i_add_term2[4]), .Y(_64_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term1[4]), .B(_64_), .Y(_65_) );
INVX1 INVX1_89 ( .A(i_add_term1[5]), .Y(_66_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[5]), .B(_66_), .Y(_67_) );
INVX1 INVX1_90 ( .A(i_add_term2[5]), .Y(_68_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term1[5]), .B(_68_), .Y(_69_) );
OAI22X1 OAI22X1_5 ( .A(_63_), .B(_65_), .C(_67_), .D(_69_), .Y(_70_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_71_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_72_) );
NOR2X1 NOR2X1_101 ( .A(_71_), .B(_72_), .Y(_73_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_74_) );
NAND2X1 NAND2X1_136 ( .A(_73_), .B(_74_), .Y(_75_) );
NOR2X1 NOR2X1_102 ( .A(_70_), .B(_75_), .Y(_6_) );
INVX1 INVX1_91 ( .A(_4_), .Y(_76_) );
NAND2X1 NAND2X1_137 ( .A(gnd), .B(_6_), .Y(_77_) );
OAI21X1 OAI21X1_132 ( .A(_6_), .B(_76_), .C(_77_), .Y(w_cout_2_) );
INVX1 INVX1_92 ( .A(i_add_term1[8]), .Y(_78_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[8]), .B(_78_), .Y(_79_) );
INVX1 INVX1_93 ( .A(i_add_term2[8]), .Y(_80_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term1[8]), .B(_80_), .Y(_81_) );
INVX1 INVX1_94 ( .A(i_add_term1[9]), .Y(_82_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[9]), .B(_82_), .Y(_83_) );
INVX1 INVX1_95 ( .A(i_add_term2[9]), .Y(_84_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term1[9]), .B(_84_), .Y(_85_) );
OAI22X1 OAI22X1_6 ( .A(_79_), .B(_81_), .C(_83_), .D(_85_), .Y(_86_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_87_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_88_) );
NOR2X1 NOR2X1_108 ( .A(_87_), .B(_88_), .Y(_89_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_90_) );
NAND2X1 NAND2X1_138 ( .A(_89_), .B(_90_), .Y(_91_) );
NOR2X1 NOR2X1_109 ( .A(_86_), .B(_91_), .Y(_9_) );
INVX1 INVX1_96 ( .A(_7_), .Y(_92_) );
NAND2X1 NAND2X1_139 ( .A(gnd), .B(_9_), .Y(_93_) );
OAI21X1 OAI21X1_133 ( .A(_9_), .B(_92_), .C(_93_), .Y(w_cout_3_) );
INVX1 INVX1_97 ( .A(i_add_term1[12]), .Y(_94_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term2[12]), .B(_94_), .Y(_95_) );
INVX1 INVX1_98 ( .A(i_add_term2[12]), .Y(_96_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term1[12]), .B(_96_), .Y(_97_) );
INVX1 INVX1_99 ( .A(i_add_term1[13]), .Y(_98_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term2[13]), .B(_98_), .Y(_99_) );
INVX1 INVX1_100 ( .A(i_add_term2[13]), .Y(_100_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term1[13]), .B(_100_), .Y(_101_) );
OAI22X1 OAI22X1_7 ( .A(_95_), .B(_97_), .C(_99_), .D(_101_), .Y(_102_) );
NOR2X1 NOR2X1_114 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_103_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_104_) );
NOR2X1 NOR2X1_115 ( .A(_103_), .B(_104_), .Y(_105_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_106_) );
NAND2X1 NAND2X1_140 ( .A(_105_), .B(_106_), .Y(_107_) );
NOR2X1 NOR2X1_116 ( .A(_102_), .B(_107_), .Y(_12_) );
INVX1 INVX1_101 ( .A(_10_), .Y(_108_) );
NAND2X1 NAND2X1_141 ( .A(gnd), .B(_12_), .Y(_109_) );
OAI21X1 OAI21X1_134 ( .A(_12_), .B(_108_), .C(_109_), .Y(w_cout_4_) );
INVX1 INVX1_102 ( .A(i_add_term1[16]), .Y(_110_) );
NOR2X1 NOR2X1_117 ( .A(i_add_term2[16]), .B(_110_), .Y(_111_) );
INVX1 INVX1_103 ( .A(i_add_term2[16]), .Y(_112_) );
NOR2X1 NOR2X1_118 ( .A(i_add_term1[16]), .B(_112_), .Y(_113_) );
INVX1 INVX1_104 ( .A(i_add_term1[17]), .Y(_114_) );
NOR2X1 NOR2X1_119 ( .A(i_add_term2[17]), .B(_114_), .Y(_115_) );
INVX1 INVX1_105 ( .A(i_add_term2[17]), .Y(_116_) );
NOR2X1 NOR2X1_120 ( .A(i_add_term1[17]), .B(_116_), .Y(_117_) );
OAI22X1 OAI22X1_8 ( .A(_111_), .B(_113_), .C(_115_), .D(_117_), .Y(_118_) );
NOR2X1 NOR2X1_121 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_119_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_120_) );
NOR2X1 NOR2X1_122 ( .A(_119_), .B(_120_), .Y(_121_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_122_) );
NAND2X1 NAND2X1_142 ( .A(_121_), .B(_122_), .Y(_123_) );
NOR2X1 NOR2X1_123 ( .A(_118_), .B(_123_), .Y(_15_) );
INVX1 INVX1_106 ( .A(_13_), .Y(_124_) );
NAND2X1 NAND2X1_143 ( .A(gnd), .B(_15_), .Y(_125_) );
OAI21X1 OAI21X1_135 ( .A(_15_), .B(_124_), .C(_125_), .Y(w_cout_5_) );
INVX1 INVX1_107 ( .A(i_add_term1[20]), .Y(_126_) );
NOR2X1 NOR2X1_124 ( .A(i_add_term2[20]), .B(_126_), .Y(_127_) );
INVX1 INVX1_108 ( .A(i_add_term2[20]), .Y(_128_) );
NOR2X1 NOR2X1_125 ( .A(i_add_term1[20]), .B(_128_), .Y(_129_) );
INVX1 INVX1_109 ( .A(i_add_term1[21]), .Y(_130_) );
NOR2X1 NOR2X1_126 ( .A(i_add_term2[21]), .B(_130_), .Y(_131_) );
INVX1 INVX1_110 ( .A(i_add_term2[21]), .Y(_132_) );
NOR2X1 NOR2X1_127 ( .A(i_add_term1[21]), .B(_132_), .Y(_133_) );
OAI22X1 OAI22X1_9 ( .A(_127_), .B(_129_), .C(_131_), .D(_133_), .Y(_134_) );
NOR2X1 NOR2X1_128 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_135_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_136_) );
NOR2X1 NOR2X1_129 ( .A(_135_), .B(_136_), .Y(_137_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_138_) );
NAND2X1 NAND2X1_144 ( .A(_137_), .B(_138_), .Y(_139_) );
NOR2X1 NOR2X1_130 ( .A(_134_), .B(_139_), .Y(_18_) );
INVX1 INVX1_111 ( .A(_16_), .Y(_140_) );
NAND2X1 NAND2X1_145 ( .A(gnd), .B(_18_), .Y(_141_) );
OAI21X1 OAI21X1_136 ( .A(_18_), .B(_140_), .C(_141_), .Y(w_cout_6_) );
INVX1 INVX1_112 ( .A(i_add_term1[24]), .Y(_142_) );
NOR2X1 NOR2X1_131 ( .A(i_add_term2[24]), .B(_142_), .Y(_143_) );
INVX1 INVX1_113 ( .A(i_add_term2[24]), .Y(_144_) );
NOR2X1 NOR2X1_132 ( .A(i_add_term1[24]), .B(_144_), .Y(_145_) );
INVX1 INVX1_114 ( .A(i_add_term1[25]), .Y(_146_) );
NOR2X1 NOR2X1_133 ( .A(i_add_term2[25]), .B(_146_), .Y(_147_) );
INVX1 INVX1_115 ( .A(i_add_term2[25]), .Y(_148_) );
NOR2X1 NOR2X1_134 ( .A(i_add_term1[25]), .B(_148_), .Y(_149_) );
OAI22X1 OAI22X1_10 ( .A(_143_), .B(_145_), .C(_147_), .D(_149_), .Y(_150_) );
NOR2X1 NOR2X1_135 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_151_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_152_) );
NOR2X1 NOR2X1_136 ( .A(_151_), .B(_152_), .Y(_153_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_154_) );
NAND2X1 NAND2X1_146 ( .A(_153_), .B(_154_), .Y(_155_) );
NOR2X1 NOR2X1_137 ( .A(_150_), .B(_155_), .Y(_21_) );
INVX1 INVX1_116 ( .A(_19_), .Y(_156_) );
NAND2X1 NAND2X1_147 ( .A(gnd), .B(_21_), .Y(_157_) );
OAI21X1 OAI21X1_137 ( .A(_21_), .B(_156_), .C(_157_), .Y(w_cout_7_) );
INVX1 INVX1_117 ( .A(i_add_term1[28]), .Y(_158_) );
NOR2X1 NOR2X1_138 ( .A(i_add_term2[28]), .B(_158_), .Y(_159_) );
INVX1 INVX1_118 ( .A(i_add_term2[28]), .Y(_160_) );
NOR2X1 NOR2X1_139 ( .A(i_add_term1[28]), .B(_160_), .Y(_161_) );
INVX1 INVX1_119 ( .A(i_add_term1[29]), .Y(_162_) );
NOR2X1 NOR2X1_140 ( .A(i_add_term2[29]), .B(_162_), .Y(_163_) );
INVX1 INVX1_120 ( .A(i_add_term2[29]), .Y(_164_) );
NOR2X1 NOR2X1_141 ( .A(i_add_term1[29]), .B(_164_), .Y(_165_) );
OAI22X1 OAI22X1_11 ( .A(_159_), .B(_161_), .C(_163_), .D(_165_), .Y(_166_) );
NOR2X1 NOR2X1_142 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_167_) );
AND2X2 AND2X2_73 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_168_) );
NOR2X1 NOR2X1_143 ( .A(_167_), .B(_168_), .Y(_169_) );
XOR2X1 XOR2X1_11 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_170_) );
NAND2X1 NAND2X1_148 ( .A(_169_), .B(_170_), .Y(_171_) );
NOR2X1 NOR2X1_144 ( .A(_166_), .B(_171_), .Y(_24_) );
INVX1 INVX1_121 ( .A(_22_), .Y(_172_) );
NAND2X1 NAND2X1_149 ( .A(gnd), .B(_24_), .Y(_173_) );
OAI21X1 OAI21X1_138 ( .A(_24_), .B(_172_), .C(_173_), .Y(w_cout_8_) );
INVX1 INVX1_122 ( .A(i_add_term1[32]), .Y(_174_) );
NOR2X1 NOR2X1_145 ( .A(i_add_term2[32]), .B(_174_), .Y(_175_) );
INVX1 INVX1_123 ( .A(i_add_term2[32]), .Y(_176_) );
NOR2X1 NOR2X1_146 ( .A(i_add_term1[32]), .B(_176_), .Y(_177_) );
INVX1 INVX1_124 ( .A(i_add_term1[33]), .Y(_178_) );
NOR2X1 NOR2X1_147 ( .A(i_add_term2[33]), .B(_178_), .Y(_179_) );
INVX1 INVX1_125 ( .A(i_add_term2[33]), .Y(_180_) );
NOR2X1 NOR2X1_148 ( .A(i_add_term1[33]), .B(_180_), .Y(_181_) );
OAI22X1 OAI22X1_12 ( .A(_175_), .B(_177_), .C(_179_), .D(_181_), .Y(_182_) );
NOR2X1 NOR2X1_149 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_183_) );
AND2X2 AND2X2_74 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_184_) );
NOR2X1 NOR2X1_150 ( .A(_183_), .B(_184_), .Y(_185_) );
XOR2X1 XOR2X1_12 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_186_) );
NAND2X1 NAND2X1_150 ( .A(_185_), .B(_186_), .Y(_187_) );
NOR2X1 NOR2X1_151 ( .A(_182_), .B(_187_), .Y(_27_) );
INVX1 INVX1_126 ( .A(_25_), .Y(_188_) );
NAND2X1 NAND2X1_151 ( .A(gnd), .B(_27_), .Y(_189_) );
OAI21X1 OAI21X1_139 ( .A(_27_), .B(_188_), .C(_189_), .Y(w_cout_9_) );
INVX1 INVX1_127 ( .A(i_add_term1[36]), .Y(_190_) );
NOR2X1 NOR2X1_152 ( .A(i_add_term2[36]), .B(_190_), .Y(_191_) );
INVX1 INVX1_128 ( .A(i_add_term2[36]), .Y(_192_) );
NOR2X1 NOR2X1_153 ( .A(i_add_term1[36]), .B(_192_), .Y(_193_) );
INVX1 INVX1_129 ( .A(i_add_term1[37]), .Y(_194_) );
NOR2X1 NOR2X1_154 ( .A(i_add_term2[37]), .B(_194_), .Y(_195_) );
INVX1 INVX1_130 ( .A(i_add_term2[37]), .Y(_196_) );
NOR2X1 NOR2X1_155 ( .A(i_add_term1[37]), .B(_196_), .Y(_197_) );
OAI22X1 OAI22X1_13 ( .A(_191_), .B(_193_), .C(_195_), .D(_197_), .Y(_198_) );
NOR2X1 NOR2X1_156 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_199_) );
AND2X2 AND2X2_75 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_200_) );
NOR2X1 NOR2X1_157 ( .A(_199_), .B(_200_), .Y(_201_) );
XOR2X1 XOR2X1_13 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_202_) );
NAND2X1 NAND2X1_152 ( .A(_201_), .B(_202_), .Y(_203_) );
NOR2X1 NOR2X1_158 ( .A(_198_), .B(_203_), .Y(_30_) );
INVX1 INVX1_131 ( .A(_28_), .Y(_204_) );
NAND2X1 NAND2X1_153 ( .A(gnd), .B(_30_), .Y(_205_) );
OAI21X1 OAI21X1_140 ( .A(_30_), .B(_204_), .C(_205_), .Y(w_cout_10_) );
INVX1 INVX1_132 ( .A(i_add_term1[40]), .Y(_206_) );
NOR2X1 NOR2X1_159 ( .A(i_add_term2[40]), .B(_206_), .Y(_207_) );
INVX1 INVX1_133 ( .A(i_add_term2[40]), .Y(_208_) );
NOR2X1 NOR2X1_160 ( .A(i_add_term1[40]), .B(_208_), .Y(_209_) );
INVX1 INVX1_134 ( .A(i_add_term1[41]), .Y(_210_) );
NOR2X1 NOR2X1_161 ( .A(i_add_term2[41]), .B(_210_), .Y(_211_) );
INVX1 INVX1_135 ( .A(i_add_term2[41]), .Y(_212_) );
NOR2X1 NOR2X1_162 ( .A(i_add_term1[41]), .B(_212_), .Y(_213_) );
OAI22X1 OAI22X1_14 ( .A(_207_), .B(_209_), .C(_211_), .D(_213_), .Y(_214_) );
NOR2X1 NOR2X1_163 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_215_) );
AND2X2 AND2X2_76 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_216_) );
NOR2X1 NOR2X1_164 ( .A(_215_), .B(_216_), .Y(_217_) );
XOR2X1 XOR2X1_14 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_218_) );
NAND2X1 NAND2X1_154 ( .A(_217_), .B(_218_), .Y(_219_) );
NOR2X1 NOR2X1_165 ( .A(_214_), .B(_219_), .Y(_33_) );
INVX1 INVX1_136 ( .A(_31_), .Y(_220_) );
NAND2X1 NAND2X1_155 ( .A(gnd), .B(_33_), .Y(_221_) );
OAI21X1 OAI21X1_141 ( .A(_33_), .B(_220_), .C(_221_), .Y(w_cout_11_) );
INVX1 INVX1_137 ( .A(i_add_term1[44]), .Y(_222_) );
NOR2X1 NOR2X1_166 ( .A(i_add_term2[44]), .B(_222_), .Y(_223_) );
INVX1 INVX1_138 ( .A(i_add_term2[44]), .Y(_224_) );
NOR2X1 NOR2X1_167 ( .A(i_add_term1[44]), .B(_224_), .Y(_225_) );
INVX1 INVX1_139 ( .A(i_add_term1[45]), .Y(_226_) );
NOR2X1 NOR2X1_168 ( .A(i_add_term2[45]), .B(_226_), .Y(_227_) );
INVX1 INVX1_140 ( .A(i_add_term2[45]), .Y(_228_) );
NOR2X1 NOR2X1_169 ( .A(i_add_term1[45]), .B(_228_), .Y(_229_) );
OAI22X1 OAI22X1_15 ( .A(_223_), .B(_225_), .C(_227_), .D(_229_), .Y(_230_) );
NOR2X1 NOR2X1_170 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_231_) );
AND2X2 AND2X2_77 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_232_) );
NOR2X1 NOR2X1_171 ( .A(_231_), .B(_232_), .Y(_233_) );
XOR2X1 XOR2X1_15 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_234_) );
NAND2X1 NAND2X1_156 ( .A(_233_), .B(_234_), .Y(_235_) );
BUFX2 BUFX2_63 ( .A(cskip1_inst_sum), .Y(_0__60_) );
BUFX2 BUFX2_64 ( .A(gnd), .Y(_2__0_) );
BUFX2 BUFX2_65 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_66 ( .A(w_cout_1_), .Y(_5__0_) );
BUFX2 BUFX2_67 ( .A(_4_), .Y(_5__4_) );
BUFX2 BUFX2_68 ( .A(w_cout_2_), .Y(_8__0_) );
BUFX2 BUFX2_69 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_70 ( .A(w_cout_3_), .Y(_11__0_) );
BUFX2 BUFX2_71 ( .A(_10_), .Y(_11__4_) );
BUFX2 BUFX2_72 ( .A(w_cout_4_), .Y(_14__0_) );
BUFX2 BUFX2_73 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_74 ( .A(w_cout_5_), .Y(_17__0_) );
BUFX2 BUFX2_75 ( .A(_16_), .Y(_17__4_) );
BUFX2 BUFX2_76 ( .A(w_cout_6_), .Y(_20__0_) );
BUFX2 BUFX2_77 ( .A(_19_), .Y(_20__4_) );
BUFX2 BUFX2_78 ( .A(w_cout_7_), .Y(_23__0_) );
BUFX2 BUFX2_79 ( .A(_22_), .Y(_23__4_) );
BUFX2 BUFX2_80 ( .A(w_cout_8_), .Y(_26__0_) );
BUFX2 BUFX2_81 ( .A(_25_), .Y(_26__4_) );
BUFX2 BUFX2_82 ( .A(w_cout_9_), .Y(_29__0_) );
BUFX2 BUFX2_83 ( .A(_28_), .Y(_29__4_) );
BUFX2 BUFX2_84 ( .A(w_cout_10_), .Y(_32__0_) );
BUFX2 BUFX2_85 ( .A(_31_), .Y(_32__4_) );
BUFX2 BUFX2_86 ( .A(w_cout_11_), .Y(_35__0_) );
BUFX2 BUFX2_87 ( .A(_34_), .Y(_35__4_) );
BUFX2 BUFX2_88 ( .A(w_cout_12_), .Y(_38__0_) );
BUFX2 BUFX2_89 ( .A(_37_), .Y(_38__4_) );
BUFX2 BUFX2_90 ( .A(w_cout_13_), .Y(_41__0_) );
BUFX2 BUFX2_91 ( .A(_40_), .Y(_41__4_) );
BUFX2 BUFX2_92 ( .A(w_cout_14_), .Y(_44__0_) );
BUFX2 BUFX2_93 ( .A(_43_), .Y(_44__4_) );
BUFX2 BUFX2_94 ( .A(cskip1_inst_cin), .Y(cskip1_inst_rca0_w_CARRY_0_) );
BUFX2 BUFX2_95 ( .A(cskip1_inst_cout0), .Y(cskip1_inst_rca0_w_CARRY_4_) );
BUFX2 BUFX2_96 ( .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_97 ( .A(cskip1_inst_cin), .Y(w_cout_15_) );
endmodule
