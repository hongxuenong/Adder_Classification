module csa_6bit ( gnd, vdd, i_add_term1, i_add_term2, sum, cout);

input gnd, vdd;
output cout;
input [5:0] i_add_term1;
input [5:0] i_add_term2;
output [5:0] sum;

NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_27_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_27_), .C(_26_), .Y(_28_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_22_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_23_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_23_), .C(vdd), .Y(_24_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_28_), .Y(csa_inst_rca0_1_fa0_o_sum) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_22_), .C(_27_), .Y(csa_inst_rca0_1_c) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_1_c), .Y(_32_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_33_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_34_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_34_), .C(_33_), .Y(_35_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_29_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_30_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_30_), .C(csa_inst_rca0_1_c), .Y(_31_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_35_), .Y(csa_inst_rca0_1_fa31_o_sum) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_29_), .C(_34_), .Y(csa_inst_cout0_1) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_39_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_40_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_41_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_41_), .C(_40_), .Y(_42_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_36_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_37_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_37_), .C(gnd), .Y(_38_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_42_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_36_), .C(_41_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_i_carry), .Y(_46_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_47_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_48_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_48_), .C(_47_), .Y(_49_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_43_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_44_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_44_), .C(rca_inst_fa3_i_carry), .Y(_45_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_49_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_43_), .C(_48_), .Y(csa_inst_cin) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_carry), .Y(_53_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_54_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_55_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_55_), .C(_54_), .Y(_56_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_50_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_51_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_51_), .C(rca_inst_fa0_o_carry), .Y(_52_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_56_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_50_), .C(_55_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_carry), .Y(_60_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_61_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_62_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_62_), .C(_61_), .Y(_63_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_57_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_58_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_58_), .C(rca_inst_fa_1__o_carry), .Y(_59_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_63_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_57_), .C(_62_), .Y(rca_inst_fa3_i_carry) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(cout) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_1__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_1__5_), .Y(sum[5]) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cout0_0), .Y(_2_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cout0_1), .B(csa_inst_cin), .Y(_3_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .B(_2_), .C(_3_), .Y(_0_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_0_fa0_o_sum), .Y(_6_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_1_fa0_o_sum), .B(csa_inst_cin), .Y(_7_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .B(_6_), .C(_7_), .Y(_1__4_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_0_fa31_o_sum), .Y(_4_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .B(csa_inst_rca0_1_fa31_o_sum), .Y(_5_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .B(_4_), .C(_5_), .Y(_1__5_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_11_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_12_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_13_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_13_), .C(_12_), .Y(_14_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_8_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_9_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_9_), .C(gnd), .Y(_10_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_14_), .Y(csa_inst_rca0_0_fa0_o_sum) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_8_), .C(_13_), .Y(csa_inst_rca0_0_c) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_0_c), .Y(_18_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_19_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_20_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_20_), .C(_19_), .Y(_21_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_15_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_16_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_16_), .C(csa_inst_rca0_0_c), .Y(_17_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_21_), .Y(csa_inst_rca0_0_fa31_o_sum) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_15_), .C(_20_), .Y(csa_inst_cout0_0) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_25_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_26_) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_sum), .Y(_1__0_) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_sum), .Y(_1__1_) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_2__o_sum), .Y(_1__2_) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_o_sum), .Y(_1__3_) );
endmodule
