module cla_29bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add1[19], i_add1[20], i_add1[21], i_add1[22], i_add1[23], i_add1[24], i_add1[25], i_add1[26], i_add1[27], i_add1[28], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], i_add2[19], i_add2[20], i_add2[21], i_add2[22], i_add2[23], i_add2[24], i_add2[25], i_add2[26], i_add2[27], i_add2[28], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21], o_result[22], o_result[23], o_result[24], o_result[25], o_result[26], o_result[27], o_result[28], o_result[29]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add1[19];
input i_add1[20];
input i_add1[21];
input i_add1[22];
input i_add1[23];
input i_add1[24];
input i_add1[25];
input i_add1[26];
input i_add1[27];
input i_add1[28];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
input i_add2[19];
input i_add2[20];
input i_add2[21];
input i_add2[22];
input i_add2[23];
input i_add2[24];
input i_add2[25];
input i_add2[26];
input i_add2[27];
input i_add2[28];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];
output o_result[22];
output o_result[23];
output o_result[24];
output o_result[25];
output o_result[26];
output o_result[27];
output o_result[28];
output o_result[29];

NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_148_) );
INVX1 INVX1_1 ( .A(_148_), .Y(w_C_1_) );
NAND2X1 NAND2X1_2 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_149_) );
NAND2X1 NAND2X1_3 ( .A(_148_), .B(_149_), .Y(_150_) );
OAI21X1 OAI21X1_1 ( .A(i_add2[1]), .B(i_add1[1]), .C(_150_), .Y(_151_) );
INVX1 INVX1_2 ( .A(_151_), .Y(w_C_2_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_152_) );
OR2X2 OR2X2_1 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_153_) );
OR2X2 OR2X2_2 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_154_) );
NAND3X1 NAND3X1_1 ( .A(_153_), .B(_154_), .C(_150_), .Y(_155_) );
NAND2X1 NAND2X1_5 ( .A(_152_), .B(_155_), .Y(w_C_3_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_156_) );
NAND3X1 NAND3X1_2 ( .A(_152_), .B(_156_), .C(_155_), .Y(_0_) );
OAI21X1 OAI21X1_2 ( .A(i_add2[3]), .B(i_add1[3]), .C(_0_), .Y(_1_) );
INVX1 INVX1_3 ( .A(_1_), .Y(w_C_4_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_2_) );
OR2X2 OR2X2_3 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_3_) );
OR2X2 OR2X2_4 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_4_) );
NAND3X1 NAND3X1_3 ( .A(_3_), .B(_4_), .C(_0_), .Y(_5_) );
NAND2X1 NAND2X1_8 ( .A(_2_), .B(_5_), .Y(w_C_5_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_6_) );
NAND3X1 NAND3X1_4 ( .A(_2_), .B(_6_), .C(_5_), .Y(_7_) );
OAI21X1 OAI21X1_3 ( .A(i_add2[5]), .B(i_add1[5]), .C(_7_), .Y(_8_) );
INVX1 INVX1_4 ( .A(_8_), .Y(w_C_6_) );
INVX1 INVX1_5 ( .A(i_add2[6]), .Y(_9_) );
INVX1 INVX1_6 ( .A(i_add1[6]), .Y(_10_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_11_) );
INVX1 INVX1_7 ( .A(_11_), .Y(_12_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_13_) );
INVX1 INVX1_8 ( .A(_13_), .Y(_14_) );
NAND3X1 NAND3X1_5 ( .A(_12_), .B(_14_), .C(_7_), .Y(_15_) );
OAI21X1 OAI21X1_4 ( .A(_9_), .B(_10_), .C(_15_), .Y(w_C_7_) );
NOR2X1 NOR2X1_3 ( .A(_9_), .B(_10_), .Y(_16_) );
INVX1 INVX1_9 ( .A(_16_), .Y(_17_) );
AND2X2 AND2X2_1 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_18_) );
INVX1 INVX1_10 ( .A(_18_), .Y(_19_) );
NAND3X1 NAND3X1_6 ( .A(_17_), .B(_19_), .C(_15_), .Y(_20_) );
OAI21X1 OAI21X1_5 ( .A(i_add2[7]), .B(i_add1[7]), .C(_20_), .Y(_21_) );
INVX1 INVX1_11 ( .A(_21_), .Y(w_C_8_) );
INVX1 INVX1_12 ( .A(i_add2[8]), .Y(_22_) );
INVX1 INVX1_13 ( .A(i_add1[8]), .Y(_23_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_24_) );
INVX1 INVX1_14 ( .A(_24_), .Y(_25_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_26_) );
INVX1 INVX1_15 ( .A(_26_), .Y(_27_) );
NAND3X1 NAND3X1_7 ( .A(_25_), .B(_27_), .C(_20_), .Y(_28_) );
OAI21X1 OAI21X1_6 ( .A(_22_), .B(_23_), .C(_28_), .Y(w_C_9_) );
NOR2X1 NOR2X1_6 ( .A(_22_), .B(_23_), .Y(_29_) );
INVX1 INVX1_16 ( .A(_29_), .Y(_30_) );
AND2X2 AND2X2_2 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_31_) );
INVX1 INVX1_17 ( .A(_31_), .Y(_32_) );
NAND3X1 NAND3X1_8 ( .A(_30_), .B(_32_), .C(_28_), .Y(_33_) );
OAI21X1 OAI21X1_7 ( .A(i_add2[9]), .B(i_add1[9]), .C(_33_), .Y(_34_) );
INVX1 INVX1_18 ( .A(_34_), .Y(w_C_10_) );
INVX1 INVX1_19 ( .A(i_add2[10]), .Y(_35_) );
INVX1 INVX1_20 ( .A(i_add1[10]), .Y(_36_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_37_) );
INVX1 INVX1_21 ( .A(_37_), .Y(_38_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_39_) );
INVX1 INVX1_22 ( .A(_39_), .Y(_40_) );
NAND3X1 NAND3X1_9 ( .A(_38_), .B(_40_), .C(_33_), .Y(_41_) );
OAI21X1 OAI21X1_8 ( .A(_35_), .B(_36_), .C(_41_), .Y(w_C_11_) );
NOR2X1 NOR2X1_9 ( .A(_35_), .B(_36_), .Y(_42_) );
INVX1 INVX1_23 ( .A(_42_), .Y(_43_) );
AND2X2 AND2X2_3 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_44_) );
INVX1 INVX1_24 ( .A(_44_), .Y(_45_) );
NAND3X1 NAND3X1_10 ( .A(_43_), .B(_45_), .C(_41_), .Y(_46_) );
OAI21X1 OAI21X1_9 ( .A(i_add2[11]), .B(i_add1[11]), .C(_46_), .Y(_47_) );
INVX1 INVX1_25 ( .A(_47_), .Y(w_C_12_) );
INVX1 INVX1_26 ( .A(i_add2[12]), .Y(_48_) );
INVX1 INVX1_27 ( .A(i_add1[12]), .Y(_49_) );
NOR2X1 NOR2X1_10 ( .A(_48_), .B(_49_), .Y(_50_) );
INVX1 INVX1_28 ( .A(_50_), .Y(_51_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_52_) );
INVX1 INVX1_29 ( .A(_52_), .Y(_53_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_54_) );
INVX1 INVX1_30 ( .A(_54_), .Y(_55_) );
NAND3X1 NAND3X1_11 ( .A(_53_), .B(_55_), .C(_46_), .Y(_56_) );
AND2X2 AND2X2_4 ( .A(_56_), .B(_51_), .Y(_57_) );
INVX1 INVX1_31 ( .A(_57_), .Y(w_C_13_) );
AND2X2 AND2X2_5 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_58_) );
INVX1 INVX1_32 ( .A(_58_), .Y(_59_) );
NAND3X1 NAND3X1_12 ( .A(_51_), .B(_59_), .C(_56_), .Y(_60_) );
OAI21X1 OAI21X1_10 ( .A(i_add2[13]), .B(i_add1[13]), .C(_60_), .Y(_61_) );
INVX1 INVX1_33 ( .A(_61_), .Y(w_C_14_) );
INVX1 INVX1_34 ( .A(i_add2[14]), .Y(_62_) );
INVX1 INVX1_35 ( .A(i_add1[14]), .Y(_63_) );
NOR2X1 NOR2X1_13 ( .A(_62_), .B(_63_), .Y(_64_) );
INVX1 INVX1_36 ( .A(_64_), .Y(_65_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_66_) );
INVX1 INVX1_37 ( .A(_66_), .Y(_67_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_68_) );
INVX1 INVX1_38 ( .A(_68_), .Y(_69_) );
NAND3X1 NAND3X1_13 ( .A(_67_), .B(_69_), .C(_60_), .Y(_70_) );
AND2X2 AND2X2_6 ( .A(_70_), .B(_65_), .Y(_71_) );
INVX1 INVX1_39 ( .A(_71_), .Y(w_C_15_) );
AND2X2 AND2X2_7 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_72_) );
INVX1 INVX1_40 ( .A(_72_), .Y(_73_) );
NAND3X1 NAND3X1_14 ( .A(_65_), .B(_73_), .C(_70_), .Y(_74_) );
OAI21X1 OAI21X1_11 ( .A(i_add2[15]), .B(i_add1[15]), .C(_74_), .Y(_75_) );
INVX1 INVX1_41 ( .A(_75_), .Y(w_C_16_) );
INVX1 INVX1_42 ( .A(i_add2[16]), .Y(_76_) );
INVX1 INVX1_43 ( .A(i_add1[16]), .Y(_77_) );
NOR2X1 NOR2X1_16 ( .A(_76_), .B(_77_), .Y(_78_) );
INVX1 INVX1_44 ( .A(_78_), .Y(_79_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_80_) );
INVX1 INVX1_45 ( .A(_80_), .Y(_81_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_82_) );
INVX1 INVX1_46 ( .A(_82_), .Y(_83_) );
NAND3X1 NAND3X1_15 ( .A(_81_), .B(_83_), .C(_74_), .Y(_84_) );
AND2X2 AND2X2_8 ( .A(_84_), .B(_79_), .Y(_85_) );
INVX1 INVX1_47 ( .A(_85_), .Y(w_C_17_) );
AND2X2 AND2X2_9 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_86_) );
INVX1 INVX1_48 ( .A(_86_), .Y(_87_) );
NAND3X1 NAND3X1_16 ( .A(_79_), .B(_87_), .C(_84_), .Y(_88_) );
OAI21X1 OAI21X1_12 ( .A(i_add2[17]), .B(i_add1[17]), .C(_88_), .Y(_89_) );
INVX1 INVX1_49 ( .A(_89_), .Y(w_C_18_) );
INVX1 INVX1_50 ( .A(i_add2[18]), .Y(_90_) );
INVX1 INVX1_51 ( .A(i_add1[18]), .Y(_91_) );
NOR2X1 NOR2X1_19 ( .A(_90_), .B(_91_), .Y(_92_) );
INVX1 INVX1_52 ( .A(_92_), .Y(_93_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_94_) );
INVX1 INVX1_53 ( .A(_94_), .Y(_95_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_96_) );
INVX1 INVX1_54 ( .A(_96_), .Y(_97_) );
NAND3X1 NAND3X1_17 ( .A(_95_), .B(_97_), .C(_88_), .Y(_98_) );
AND2X2 AND2X2_10 ( .A(_98_), .B(_93_), .Y(_99_) );
INVX1 INVX1_55 ( .A(_99_), .Y(w_C_19_) );
AND2X2 AND2X2_11 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_100_) );
INVX1 INVX1_56 ( .A(_100_), .Y(_101_) );
NAND3X1 NAND3X1_18 ( .A(_93_), .B(_101_), .C(_98_), .Y(_102_) );
OAI21X1 OAI21X1_13 ( .A(i_add2[19]), .B(i_add1[19]), .C(_102_), .Y(_103_) );
INVX1 INVX1_57 ( .A(_103_), .Y(w_C_20_) );
INVX1 INVX1_58 ( .A(i_add2[20]), .Y(_104_) );
INVX1 INVX1_59 ( .A(i_add1[20]), .Y(_105_) );
NOR2X1 NOR2X1_22 ( .A(_104_), .B(_105_), .Y(_106_) );
INVX1 INVX1_60 ( .A(_106_), .Y(_107_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_108_) );
INVX1 INVX1_61 ( .A(_108_), .Y(_109_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_110_) );
INVX1 INVX1_62 ( .A(_110_), .Y(_111_) );
NAND3X1 NAND3X1_19 ( .A(_109_), .B(_111_), .C(_102_), .Y(_112_) );
AND2X2 AND2X2_12 ( .A(_112_), .B(_107_), .Y(_113_) );
INVX1 INVX1_63 ( .A(_113_), .Y(w_C_21_) );
AND2X2 AND2X2_13 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_114_) );
INVX1 INVX1_64 ( .A(_114_), .Y(_115_) );
NAND3X1 NAND3X1_20 ( .A(_107_), .B(_115_), .C(_112_), .Y(_116_) );
OAI21X1 OAI21X1_14 ( .A(i_add2[21]), .B(i_add1[21]), .C(_116_), .Y(_117_) );
INVX1 INVX1_65 ( .A(_117_), .Y(w_C_22_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_118_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_119_) );
OAI21X1 OAI21X1_15 ( .A(_119_), .B(_117_), .C(_118_), .Y(w_C_23_) );
OR2X2 OR2X2_5 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_120_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_121_) );
INVX1 INVX1_66 ( .A(_121_), .Y(_122_) );
INVX1 INVX1_67 ( .A(_119_), .Y(_123_) );
NAND3X1 NAND3X1_21 ( .A(_122_), .B(_123_), .C(_116_), .Y(_124_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_125_) );
NAND3X1 NAND3X1_22 ( .A(_118_), .B(_125_), .C(_124_), .Y(_126_) );
AND2X2 AND2X2_14 ( .A(_126_), .B(_120_), .Y(w_C_24_) );
INVX1 INVX1_68 ( .A(i_add2[24]), .Y(_127_) );
INVX1 INVX1_69 ( .A(i_add1[24]), .Y(_128_) );
NAND2X1 NAND2X1_12 ( .A(_127_), .B(_128_), .Y(_129_) );
NAND3X1 NAND3X1_23 ( .A(_120_), .B(_129_), .C(_126_), .Y(_130_) );
OAI21X1 OAI21X1_16 ( .A(_127_), .B(_128_), .C(_130_), .Y(w_C_25_) );
INVX1 INVX1_70 ( .A(i_add2[25]), .Y(_131_) );
INVX1 INVX1_71 ( .A(i_add1[25]), .Y(_132_) );
NAND2X1 NAND2X1_13 ( .A(_131_), .B(_132_), .Y(_133_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_134_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_135_) );
NAND3X1 NAND3X1_24 ( .A(_134_), .B(_135_), .C(_130_), .Y(_136_) );
AND2X2 AND2X2_15 ( .A(_136_), .B(_133_), .Y(w_C_26_) );
INVX1 INVX1_72 ( .A(i_add2[26]), .Y(_137_) );
INVX1 INVX1_73 ( .A(i_add1[26]), .Y(_138_) );
NAND2X1 NAND2X1_16 ( .A(_137_), .B(_138_), .Y(_139_) );
NAND3X1 NAND3X1_25 ( .A(_133_), .B(_139_), .C(_136_), .Y(_140_) );
OAI21X1 OAI21X1_17 ( .A(_137_), .B(_138_), .C(_140_), .Y(w_C_27_) );
OR2X2 OR2X2_6 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_141_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_142_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_143_) );
NAND3X1 NAND3X1_26 ( .A(_142_), .B(_143_), .C(_140_), .Y(_144_) );
AND2X2 AND2X2_16 ( .A(_144_), .B(_141_), .Y(w_C_28_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_145_) );
OR2X2 OR2X2_7 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_146_) );
NAND3X1 NAND3X1_27 ( .A(_141_), .B(_146_), .C(_144_), .Y(_147_) );
NAND2X1 NAND2X1_20 ( .A(_145_), .B(_147_), .Y(w_C_29_) );
BUFX2 BUFX2_1 ( .A(_157__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_157__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_157__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_157__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_157__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_157__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_157__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_157__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_157__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_157__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_157__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_157__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_157__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_157__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_157__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_157__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_157__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_157__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_157__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_157__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_157__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_157__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_157__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_157__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_157__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_157__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_157__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_157__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_157__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(w_C_29_), .Y(o_result[29]) );
INVX1 INVX1_74 ( .A(w_C_4_), .Y(_161_) );
OR2X2 OR2X2_8 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_162_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_163_) );
NAND3X1 NAND3X1_28 ( .A(_161_), .B(_163_), .C(_162_), .Y(_164_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_158_) );
AND2X2 AND2X2_17 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_159_) );
OAI21X1 OAI21X1_18 ( .A(_158_), .B(_159_), .C(w_C_4_), .Y(_160_) );
NAND2X1 NAND2X1_22 ( .A(_160_), .B(_164_), .Y(_157__4_) );
INVX1 INVX1_75 ( .A(w_C_5_), .Y(_168_) );
OR2X2 OR2X2_9 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_169_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_170_) );
NAND3X1 NAND3X1_29 ( .A(_168_), .B(_170_), .C(_169_), .Y(_171_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_165_) );
AND2X2 AND2X2_18 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_166_) );
OAI21X1 OAI21X1_19 ( .A(_165_), .B(_166_), .C(w_C_5_), .Y(_167_) );
NAND2X1 NAND2X1_24 ( .A(_167_), .B(_171_), .Y(_157__5_) );
INVX1 INVX1_76 ( .A(w_C_6_), .Y(_175_) );
OR2X2 OR2X2_10 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_176_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_177_) );
NAND3X1 NAND3X1_30 ( .A(_175_), .B(_177_), .C(_176_), .Y(_178_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_172_) );
AND2X2 AND2X2_19 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_173_) );
OAI21X1 OAI21X1_20 ( .A(_172_), .B(_173_), .C(w_C_6_), .Y(_174_) );
NAND2X1 NAND2X1_26 ( .A(_174_), .B(_178_), .Y(_157__6_) );
INVX1 INVX1_77 ( .A(w_C_7_), .Y(_182_) );
OR2X2 OR2X2_11 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_183_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_184_) );
NAND3X1 NAND3X1_31 ( .A(_182_), .B(_184_), .C(_183_), .Y(_185_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_179_) );
AND2X2 AND2X2_20 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_180_) );
OAI21X1 OAI21X1_21 ( .A(_179_), .B(_180_), .C(w_C_7_), .Y(_181_) );
NAND2X1 NAND2X1_28 ( .A(_181_), .B(_185_), .Y(_157__7_) );
INVX1 INVX1_78 ( .A(w_C_8_), .Y(_189_) );
OR2X2 OR2X2_12 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_190_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_191_) );
NAND3X1 NAND3X1_32 ( .A(_189_), .B(_191_), .C(_190_), .Y(_192_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_186_) );
AND2X2 AND2X2_21 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_187_) );
OAI21X1 OAI21X1_22 ( .A(_186_), .B(_187_), .C(w_C_8_), .Y(_188_) );
NAND2X1 NAND2X1_30 ( .A(_188_), .B(_192_), .Y(_157__8_) );
INVX1 INVX1_79 ( .A(w_C_9_), .Y(_196_) );
OR2X2 OR2X2_13 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_197_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_198_) );
NAND3X1 NAND3X1_33 ( .A(_196_), .B(_198_), .C(_197_), .Y(_199_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_193_) );
AND2X2 AND2X2_22 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_194_) );
OAI21X1 OAI21X1_23 ( .A(_193_), .B(_194_), .C(w_C_9_), .Y(_195_) );
NAND2X1 NAND2X1_32 ( .A(_195_), .B(_199_), .Y(_157__9_) );
INVX1 INVX1_80 ( .A(w_C_10_), .Y(_203_) );
OR2X2 OR2X2_14 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_204_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_205_) );
NAND3X1 NAND3X1_34 ( .A(_203_), .B(_205_), .C(_204_), .Y(_206_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_200_) );
AND2X2 AND2X2_23 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_201_) );
OAI21X1 OAI21X1_24 ( .A(_200_), .B(_201_), .C(w_C_10_), .Y(_202_) );
NAND2X1 NAND2X1_34 ( .A(_202_), .B(_206_), .Y(_157__10_) );
INVX1 INVX1_81 ( .A(w_C_11_), .Y(_210_) );
OR2X2 OR2X2_15 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_211_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_212_) );
NAND3X1 NAND3X1_35 ( .A(_210_), .B(_212_), .C(_211_), .Y(_213_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_207_) );
AND2X2 AND2X2_24 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_208_) );
OAI21X1 OAI21X1_25 ( .A(_207_), .B(_208_), .C(w_C_11_), .Y(_209_) );
NAND2X1 NAND2X1_36 ( .A(_209_), .B(_213_), .Y(_157__11_) );
INVX1 INVX1_82 ( .A(w_C_12_), .Y(_217_) );
OR2X2 OR2X2_16 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_218_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_219_) );
NAND3X1 NAND3X1_36 ( .A(_217_), .B(_219_), .C(_218_), .Y(_220_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_214_) );
AND2X2 AND2X2_25 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_215_) );
OAI21X1 OAI21X1_26 ( .A(_214_), .B(_215_), .C(w_C_12_), .Y(_216_) );
NAND2X1 NAND2X1_38 ( .A(_216_), .B(_220_), .Y(_157__12_) );
INVX1 INVX1_83 ( .A(w_C_13_), .Y(_224_) );
OR2X2 OR2X2_17 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_225_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_226_) );
NAND3X1 NAND3X1_37 ( .A(_224_), .B(_226_), .C(_225_), .Y(_227_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_221_) );
AND2X2 AND2X2_26 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_222_) );
OAI21X1 OAI21X1_27 ( .A(_221_), .B(_222_), .C(w_C_13_), .Y(_223_) );
NAND2X1 NAND2X1_40 ( .A(_223_), .B(_227_), .Y(_157__13_) );
INVX1 INVX1_84 ( .A(w_C_14_), .Y(_231_) );
OR2X2 OR2X2_18 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_232_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_233_) );
NAND3X1 NAND3X1_38 ( .A(_231_), .B(_233_), .C(_232_), .Y(_234_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_228_) );
AND2X2 AND2X2_27 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_229_) );
OAI21X1 OAI21X1_28 ( .A(_228_), .B(_229_), .C(w_C_14_), .Y(_230_) );
NAND2X1 NAND2X1_42 ( .A(_230_), .B(_234_), .Y(_157__14_) );
INVX1 INVX1_85 ( .A(w_C_15_), .Y(_238_) );
OR2X2 OR2X2_19 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_239_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_240_) );
NAND3X1 NAND3X1_39 ( .A(_238_), .B(_240_), .C(_239_), .Y(_241_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_235_) );
AND2X2 AND2X2_28 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_236_) );
OAI21X1 OAI21X1_29 ( .A(_235_), .B(_236_), .C(w_C_15_), .Y(_237_) );
NAND2X1 NAND2X1_44 ( .A(_237_), .B(_241_), .Y(_157__15_) );
INVX1 INVX1_86 ( .A(w_C_16_), .Y(_245_) );
OR2X2 OR2X2_20 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_246_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_247_) );
NAND3X1 NAND3X1_40 ( .A(_245_), .B(_247_), .C(_246_), .Y(_248_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_242_) );
AND2X2 AND2X2_29 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_243_) );
OAI21X1 OAI21X1_30 ( .A(_242_), .B(_243_), .C(w_C_16_), .Y(_244_) );
NAND2X1 NAND2X1_46 ( .A(_244_), .B(_248_), .Y(_157__16_) );
INVX1 INVX1_87 ( .A(w_C_17_), .Y(_252_) );
OR2X2 OR2X2_21 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_253_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_254_) );
NAND3X1 NAND3X1_41 ( .A(_252_), .B(_254_), .C(_253_), .Y(_255_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_249_) );
AND2X2 AND2X2_30 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_250_) );
OAI21X1 OAI21X1_31 ( .A(_249_), .B(_250_), .C(w_C_17_), .Y(_251_) );
NAND2X1 NAND2X1_48 ( .A(_251_), .B(_255_), .Y(_157__17_) );
INVX1 INVX1_88 ( .A(w_C_18_), .Y(_259_) );
OR2X2 OR2X2_22 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_260_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_261_) );
NAND3X1 NAND3X1_42 ( .A(_259_), .B(_261_), .C(_260_), .Y(_262_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_256_) );
AND2X2 AND2X2_31 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_257_) );
OAI21X1 OAI21X1_32 ( .A(_256_), .B(_257_), .C(w_C_18_), .Y(_258_) );
NAND2X1 NAND2X1_50 ( .A(_258_), .B(_262_), .Y(_157__18_) );
INVX1 INVX1_89 ( .A(w_C_19_), .Y(_266_) );
OR2X2 OR2X2_23 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_267_) );
NAND2X1 NAND2X1_51 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_268_) );
NAND3X1 NAND3X1_43 ( .A(_266_), .B(_268_), .C(_267_), .Y(_269_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_263_) );
AND2X2 AND2X2_32 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_264_) );
OAI21X1 OAI21X1_33 ( .A(_263_), .B(_264_), .C(w_C_19_), .Y(_265_) );
NAND2X1 NAND2X1_52 ( .A(_265_), .B(_269_), .Y(_157__19_) );
INVX1 INVX1_90 ( .A(w_C_20_), .Y(_273_) );
OR2X2 OR2X2_24 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_274_) );
NAND2X1 NAND2X1_53 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_275_) );
NAND3X1 NAND3X1_44 ( .A(_273_), .B(_275_), .C(_274_), .Y(_276_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_270_) );
AND2X2 AND2X2_33 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_271_) );
OAI21X1 OAI21X1_34 ( .A(_270_), .B(_271_), .C(w_C_20_), .Y(_272_) );
NAND2X1 NAND2X1_54 ( .A(_272_), .B(_276_), .Y(_157__20_) );
INVX1 INVX1_91 ( .A(w_C_21_), .Y(_280_) );
OR2X2 OR2X2_25 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_281_) );
NAND2X1 NAND2X1_55 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_282_) );
NAND3X1 NAND3X1_45 ( .A(_280_), .B(_282_), .C(_281_), .Y(_283_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_277_) );
AND2X2 AND2X2_34 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_278_) );
OAI21X1 OAI21X1_35 ( .A(_277_), .B(_278_), .C(w_C_21_), .Y(_279_) );
NAND2X1 NAND2X1_56 ( .A(_279_), .B(_283_), .Y(_157__21_) );
INVX1 INVX1_92 ( .A(w_C_22_), .Y(_287_) );
OR2X2 OR2X2_26 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_288_) );
NAND2X1 NAND2X1_57 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_289_) );
NAND3X1 NAND3X1_46 ( .A(_287_), .B(_289_), .C(_288_), .Y(_290_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_284_) );
AND2X2 AND2X2_35 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_285_) );
OAI21X1 OAI21X1_36 ( .A(_284_), .B(_285_), .C(w_C_22_), .Y(_286_) );
NAND2X1 NAND2X1_58 ( .A(_286_), .B(_290_), .Y(_157__22_) );
INVX1 INVX1_93 ( .A(w_C_23_), .Y(_294_) );
OR2X2 OR2X2_27 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_295_) );
NAND2X1 NAND2X1_59 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_296_) );
NAND3X1 NAND3X1_47 ( .A(_294_), .B(_296_), .C(_295_), .Y(_297_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_291_) );
AND2X2 AND2X2_36 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_292_) );
OAI21X1 OAI21X1_37 ( .A(_291_), .B(_292_), .C(w_C_23_), .Y(_293_) );
NAND2X1 NAND2X1_60 ( .A(_293_), .B(_297_), .Y(_157__23_) );
INVX1 INVX1_94 ( .A(w_C_24_), .Y(_301_) );
OR2X2 OR2X2_28 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_302_) );
NAND2X1 NAND2X1_61 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_303_) );
NAND3X1 NAND3X1_48 ( .A(_301_), .B(_303_), .C(_302_), .Y(_304_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_298_) );
AND2X2 AND2X2_37 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_299_) );
OAI21X1 OAI21X1_38 ( .A(_298_), .B(_299_), .C(w_C_24_), .Y(_300_) );
NAND2X1 NAND2X1_62 ( .A(_300_), .B(_304_), .Y(_157__24_) );
INVX1 INVX1_95 ( .A(w_C_25_), .Y(_308_) );
OR2X2 OR2X2_29 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_309_) );
NAND2X1 NAND2X1_63 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_310_) );
NAND3X1 NAND3X1_49 ( .A(_308_), .B(_310_), .C(_309_), .Y(_311_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_305_) );
AND2X2 AND2X2_38 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_306_) );
OAI21X1 OAI21X1_39 ( .A(_305_), .B(_306_), .C(w_C_25_), .Y(_307_) );
NAND2X1 NAND2X1_64 ( .A(_307_), .B(_311_), .Y(_157__25_) );
INVX1 INVX1_96 ( .A(w_C_26_), .Y(_315_) );
OR2X2 OR2X2_30 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_316_) );
NAND2X1 NAND2X1_65 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_317_) );
NAND3X1 NAND3X1_50 ( .A(_315_), .B(_317_), .C(_316_), .Y(_318_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_312_) );
AND2X2 AND2X2_39 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_313_) );
OAI21X1 OAI21X1_40 ( .A(_312_), .B(_313_), .C(w_C_26_), .Y(_314_) );
NAND2X1 NAND2X1_66 ( .A(_314_), .B(_318_), .Y(_157__26_) );
INVX1 INVX1_97 ( .A(w_C_27_), .Y(_322_) );
OR2X2 OR2X2_31 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_323_) );
NAND2X1 NAND2X1_67 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_324_) );
NAND3X1 NAND3X1_51 ( .A(_322_), .B(_324_), .C(_323_), .Y(_325_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_319_) );
AND2X2 AND2X2_40 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_320_) );
OAI21X1 OAI21X1_41 ( .A(_319_), .B(_320_), .C(w_C_27_), .Y(_321_) );
NAND2X1 NAND2X1_68 ( .A(_321_), .B(_325_), .Y(_157__27_) );
INVX1 INVX1_98 ( .A(w_C_28_), .Y(_329_) );
OR2X2 OR2X2_32 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_330_) );
NAND2X1 NAND2X1_69 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_331_) );
NAND3X1 NAND3X1_52 ( .A(_329_), .B(_331_), .C(_330_), .Y(_332_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_326_) );
AND2X2 AND2X2_41 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_327_) );
OAI21X1 OAI21X1_42 ( .A(_326_), .B(_327_), .C(w_C_28_), .Y(_328_) );
NAND2X1 NAND2X1_70 ( .A(_328_), .B(_332_), .Y(_157__28_) );
INVX1 INVX1_99 ( .A(1'b0), .Y(_336_) );
OR2X2 OR2X2_33 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_337_) );
NAND2X1 NAND2X1_71 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_338_) );
NAND3X1 NAND3X1_53 ( .A(_336_), .B(_338_), .C(_337_), .Y(_339_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_333_) );
AND2X2 AND2X2_42 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_334_) );
OAI21X1 OAI21X1_43 ( .A(_333_), .B(_334_), .C(1'b0), .Y(_335_) );
NAND2X1 NAND2X1_72 ( .A(_335_), .B(_339_), .Y(_157__0_) );
INVX1 INVX1_100 ( .A(w_C_1_), .Y(_343_) );
OR2X2 OR2X2_34 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_344_) );
NAND2X1 NAND2X1_73 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_345_) );
NAND3X1 NAND3X1_54 ( .A(_343_), .B(_345_), .C(_344_), .Y(_346_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_340_) );
AND2X2 AND2X2_43 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_341_) );
OAI21X1 OAI21X1_44 ( .A(_340_), .B(_341_), .C(w_C_1_), .Y(_342_) );
NAND2X1 NAND2X1_74 ( .A(_342_), .B(_346_), .Y(_157__1_) );
INVX1 INVX1_101 ( .A(w_C_2_), .Y(_350_) );
OR2X2 OR2X2_35 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_351_) );
NAND2X1 NAND2X1_75 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_352_) );
NAND3X1 NAND3X1_55 ( .A(_350_), .B(_352_), .C(_351_), .Y(_353_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_347_) );
AND2X2 AND2X2_44 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_348_) );
OAI21X1 OAI21X1_45 ( .A(_347_), .B(_348_), .C(w_C_2_), .Y(_349_) );
NAND2X1 NAND2X1_76 ( .A(_349_), .B(_353_), .Y(_157__2_) );
INVX1 INVX1_102 ( .A(w_C_3_), .Y(_357_) );
OR2X2 OR2X2_36 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_358_) );
NAND2X1 NAND2X1_77 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_359_) );
NAND3X1 NAND3X1_56 ( .A(_357_), .B(_359_), .C(_358_), .Y(_360_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_354_) );
AND2X2 AND2X2_45 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_355_) );
OAI21X1 OAI21X1_46 ( .A(_354_), .B(_355_), .C(w_C_3_), .Y(_356_) );
NAND2X1 NAND2X1_78 ( .A(_356_), .B(_360_), .Y(_157__3_) );
BUFX2 BUFX2_31 ( .A(w_C_29_), .Y(_157__29_) );
BUFX2 BUFX2_32 ( .A(1'b0), .Y(w_C_0_) );
endmodule
