module CSkipA_62bit ( gnd, vdd, i_add_term1, i_add_term2, sum, cout);

input gnd, vdd;
output cout;
input [61:0] i_add_term1;
input [61:0] i_add_term2;
output [61:0] sum;

NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_215_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_216_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_216_), .Y(_217_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_218_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_218_), .Y(_219_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_219_), .Y(_12_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(_220_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_12_), .Y(_221_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_220_), .C(_221_), .Y(w_cout_4_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .Y(_225_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_226_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_227_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_227_), .C(_226_), .Y(_228_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_222_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_223_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_223_), .C(w_cout_4_), .Y(_224_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_228_), .Y(_0__16_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_222_), .C(_227_), .Y(_14__1_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_14__3_), .Y(_232_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_233_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_234_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_234_), .C(_233_), .Y(_235_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_229_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_230_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_230_), .C(_14__3_), .Y(_231_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_235_), .Y(_0__19_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_229_), .C(_234_), .Y(_13_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_14__1_), .Y(_239_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_240_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_241_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_241_), .C(_240_), .Y(_242_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_236_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_237_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_237_), .C(_14__1_), .Y(_238_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_238_), .B(_242_), .Y(_0__17_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_236_), .C(_241_), .Y(_14__2_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_14__2_), .Y(_246_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_247_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_248_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_248_), .C(_247_), .Y(_249_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_243_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_244_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_244_), .C(_14__2_), .Y(_245_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_249_), .Y(_0__18_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_243_), .C(_248_), .Y(_14__3_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[16]), .Y(_250_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(_250_), .Y(_251_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .Y(_252_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[16]), .B(_252_), .Y(_253_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[17]), .Y(_254_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(_254_), .Y(_255_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .Y(_256_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[17]), .B(_256_), .Y(_257_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_253_), .C(_255_), .D(_257_), .Y(_258_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_259_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_260_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_260_), .Y(_261_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_262_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_262_), .Y(_263_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_263_), .Y(_15_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_264_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_15_), .Y(_265_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_264_), .C(_265_), .Y(w_cout_5_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .Y(_269_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_270_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_271_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_271_), .C(_270_), .Y(_272_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_266_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_267_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_267_), .C(w_cout_5_), .Y(_268_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_272_), .Y(_0__20_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_266_), .C(_271_), .Y(_17__1_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_17__3_), .Y(_276_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_277_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_278_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_278_), .C(_277_), .Y(_279_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_273_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_274_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_274_), .C(_17__3_), .Y(_275_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_279_), .Y(_0__23_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_273_), .C(_278_), .Y(_16_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_17__1_), .Y(_283_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_284_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_285_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_283_), .B(_285_), .C(_284_), .Y(_286_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_280_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_281_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_281_), .C(_17__1_), .Y(_282_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_286_), .Y(_0__21_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_283_), .B(_280_), .C(_285_), .Y(_17__2_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_17__2_), .Y(_290_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_291_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_292_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_292_), .C(_291_), .Y(_293_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_287_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_288_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_287_), .B(_288_), .C(_17__2_), .Y(_289_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_293_), .Y(_0__22_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_287_), .C(_292_), .Y(_17__3_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[20]), .Y(_294_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(_294_), .Y(_295_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .Y(_296_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[20]), .B(_296_), .Y(_297_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[21]), .Y(_298_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(_298_), .Y(_299_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .Y(_300_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[21]), .B(_300_), .Y(_301_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_297_), .C(_299_), .D(_301_), .Y(_302_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_303_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_304_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_304_), .Y(_305_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_306_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_306_), .Y(_307_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_307_), .Y(_18_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_308_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_18_), .Y(_309_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_308_), .C(_309_), .Y(w_cout_6_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .Y(_313_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_314_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_315_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_315_), .C(_314_), .Y(_316_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_310_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_311_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_311_), .C(w_cout_6_), .Y(_312_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_316_), .Y(_0__24_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_310_), .C(_315_), .Y(_20__1_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_20__3_), .Y(_320_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_321_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_322_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_322_), .C(_321_), .Y(_323_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_317_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_318_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_318_), .C(_20__3_), .Y(_319_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_323_), .Y(_0__27_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_317_), .C(_322_), .Y(_19_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_20__1_), .Y(_327_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_328_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_329_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_329_), .C(_328_), .Y(_330_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_324_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_325_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_325_), .C(_20__1_), .Y(_326_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_330_), .Y(_0__25_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_324_), .C(_329_), .Y(_20__2_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_20__2_), .Y(_334_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_335_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_336_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_336_), .C(_335_), .Y(_337_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_331_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_332_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_332_), .C(_20__2_), .Y(_333_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_337_), .Y(_0__26_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_331_), .C(_336_), .Y(_20__3_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[24]), .Y(_338_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(_338_), .Y(_339_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .Y(_340_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[24]), .B(_340_), .Y(_341_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[25]), .Y(_342_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(_342_), .Y(_343_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .Y(_344_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[25]), .B(_344_), .Y(_345_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_341_), .C(_343_), .D(_345_), .Y(_346_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_347_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_348_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_348_), .Y(_349_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_350_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_350_), .Y(_351_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_351_), .Y(_21_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_352_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_21_), .Y(_353_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_352_), .C(_353_), .Y(w_cout_7_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .Y(_357_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_358_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_359_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_359_), .C(_358_), .Y(_360_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_354_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_355_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_355_), .C(w_cout_7_), .Y(_356_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_360_), .Y(_0__28_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_354_), .C(_359_), .Y(_23__1_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_23__3_), .Y(_364_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_365_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_366_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_366_), .C(_365_), .Y(_367_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_361_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_362_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_362_), .C(_23__3_), .Y(_363_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_367_), .Y(_0__31_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_361_), .C(_366_), .Y(_22_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_23__1_), .Y(_371_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_372_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_373_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_373_), .C(_372_), .Y(_374_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_368_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_369_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_369_), .C(_23__1_), .Y(_370_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_374_), .Y(_0__29_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_368_), .C(_373_), .Y(_23__2_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_23__2_), .Y(_378_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_379_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_380_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_380_), .C(_379_), .Y(_381_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_375_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_376_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_376_), .C(_23__2_), .Y(_377_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_381_), .Y(_0__30_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_375_), .C(_380_), .Y(_23__3_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[28]), .Y(_382_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(_382_), .Y(_383_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .Y(_384_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[28]), .B(_384_), .Y(_385_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[29]), .Y(_386_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(_386_), .Y(_387_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .Y(_388_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[29]), .B(_388_), .Y(_389_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_385_), .C(_387_), .D(_389_), .Y(_390_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_391_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_392_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_392_), .Y(_393_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_394_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_394_), .Y(_395_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_395_), .Y(_24_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_396_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_24_), .Y(_397_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_396_), .C(_397_), .Y(w_cout_8_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .Y(_401_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_402_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_403_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_403_), .C(_402_), .Y(_404_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_398_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_399_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_399_), .C(w_cout_8_), .Y(_400_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_400_), .B(_404_), .Y(_0__32_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_398_), .C(_403_), .Y(_26__1_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_26__3_), .Y(_408_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_409_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_410_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_410_), .C(_409_), .Y(_411_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_405_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_406_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_406_), .C(_26__3_), .Y(_407_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_411_), .Y(_0__35_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_405_), .C(_410_), .Y(_25_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_26__1_), .Y(_415_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_416_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_417_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_415_), .B(_417_), .C(_416_), .Y(_418_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_412_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_413_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_413_), .C(_26__1_), .Y(_414_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_414_), .B(_418_), .Y(_0__33_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_415_), .B(_412_), .C(_417_), .Y(_26__2_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_26__2_), .Y(_422_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_423_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_424_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_422_), .B(_424_), .C(_423_), .Y(_425_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_419_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_420_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_420_), .C(_26__2_), .Y(_421_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_425_), .Y(_0__34_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_422_), .B(_419_), .C(_424_), .Y(_26__3_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[32]), .Y(_426_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(_426_), .Y(_427_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .Y(_428_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[32]), .B(_428_), .Y(_429_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[33]), .Y(_430_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(_430_), .Y(_431_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .Y(_432_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[33]), .B(_432_), .Y(_433_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_427_), .B(_429_), .C(_431_), .D(_433_), .Y(_434_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_435_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_436_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_436_), .Y(_437_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_438_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_438_), .Y(_439_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_439_), .Y(_27_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(_440_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_27_), .Y(_441_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_440_), .C(_441_), .Y(w_cout_9_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .Y(_445_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_446_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_447_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_445_), .B(_447_), .C(_446_), .Y(_448_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_442_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_443_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_443_), .C(w_cout_9_), .Y(_444_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_448_), .Y(_0__36_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_445_), .B(_442_), .C(_447_), .Y(_29__1_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_29__3_), .Y(_452_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_453_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_454_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_454_), .C(_453_), .Y(_455_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_449_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_450_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_450_), .C(_29__3_), .Y(_451_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_455_), .Y(_0__39_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_449_), .C(_454_), .Y(_28_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_29__1_), .Y(_459_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_460_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_461_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_461_), .C(_460_), .Y(_462_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_456_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_457_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_456_), .B(_457_), .C(_29__1_), .Y(_458_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_462_), .Y(_0__37_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_456_), .C(_461_), .Y(_29__2_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_29__2_), .Y(_466_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_467_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_468_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_466_), .B(_468_), .C(_467_), .Y(_469_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_463_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_464_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_464_), .C(_29__2_), .Y(_465_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_469_), .Y(_0__38_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_466_), .B(_463_), .C(_468_), .Y(_29__3_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[36]), .Y(_470_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(_470_), .Y(_471_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .Y(_472_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[36]), .B(_472_), .Y(_473_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[37]), .Y(_474_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(_474_), .Y(_475_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .Y(_476_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[37]), .B(_476_), .Y(_477_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_473_), .C(_475_), .D(_477_), .Y(_478_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_479_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_480_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_480_), .Y(_481_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_482_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_482_), .Y(_483_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_483_), .Y(_30_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_28_), .Y(_484_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_30_), .Y(_485_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_484_), .C(_485_), .Y(w_cout_10_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .Y(_489_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_490_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_491_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_491_), .C(_490_), .Y(_492_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_486_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_487_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_487_), .C(w_cout_10_), .Y(_488_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_492_), .Y(_0__40_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_486_), .C(_491_), .Y(_32__1_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_32__3_), .Y(_496_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_497_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_498_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_498_), .C(_497_), .Y(_499_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_493_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_494_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_494_), .C(_32__3_), .Y(_495_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_495_), .B(_499_), .Y(_0__43_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_493_), .C(_498_), .Y(_31_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_32__1_), .Y(_503_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_504_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_505_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_505_), .C(_504_), .Y(_506_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_500_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_501_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_501_), .C(_32__1_), .Y(_502_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_502_), .B(_506_), .Y(_0__41_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_500_), .C(_505_), .Y(_32__2_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_32__2_), .Y(_510_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_511_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_512_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_512_), .C(_511_), .Y(_513_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_507_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_508_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_508_), .C(_32__2_), .Y(_509_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_513_), .Y(_0__42_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_507_), .C(_512_), .Y(_32__3_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[40]), .Y(_514_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(_514_), .Y(_515_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .Y(_516_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[40]), .B(_516_), .Y(_517_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[41]), .Y(_518_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(_518_), .Y(_519_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .Y(_520_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[41]), .B(_520_), .Y(_521_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_517_), .C(_519_), .D(_521_), .Y(_522_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_523_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_524_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_524_), .Y(_525_) );
XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_526_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_525_), .B(_526_), .Y(_527_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_522_), .B(_527_), .Y(_33_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_31_), .Y(_528_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_33_), .Y(_529_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_528_), .C(_529_), .Y(w_cout_11_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .Y(_533_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_534_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_535_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_535_), .C(_534_), .Y(_536_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_530_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_531_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_531_), .C(w_cout_11_), .Y(_532_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_532_), .B(_536_), .Y(_0__44_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_530_), .C(_535_), .Y(_35__1_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_35__3_), .Y(_540_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_541_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_542_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_542_), .C(_541_), .Y(_543_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_537_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_538_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_538_), .C(_35__3_), .Y(_539_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_539_), .B(_543_), .Y(_0__47_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_537_), .C(_542_), .Y(_34_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_35__1_), .Y(_547_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_548_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_549_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_549_), .C(_548_), .Y(_550_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_544_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_545_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_545_), .C(_35__1_), .Y(_546_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_546_), .B(_550_), .Y(_0__45_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_544_), .C(_549_), .Y(_35__2_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_35__2_), .Y(_554_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_555_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_556_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_556_), .C(_555_), .Y(_557_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_551_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_552_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_551_), .B(_552_), .C(_35__2_), .Y(_553_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_553_), .B(_557_), .Y(_0__46_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_551_), .C(_556_), .Y(_35__3_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[44]), .Y(_558_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(_558_), .Y(_559_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .Y(_560_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[44]), .B(_560_), .Y(_561_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[45]), .Y(_562_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(_562_), .Y(_563_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .Y(_564_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[45]), .B(_564_), .Y(_565_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_561_), .C(_563_), .D(_565_), .Y(_566_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_567_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_568_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_567_), .B(_568_), .Y(_569_) );
XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_570_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_569_), .B(_570_), .Y(_571_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_571_), .Y(_36_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(_34_), .Y(_572_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_36_), .Y(_573_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_572_), .C(_573_), .Y(w_cout_12_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .Y(_577_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_578_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_579_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_579_), .C(_578_), .Y(_580_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_574_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_575_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_574_), .B(_575_), .C(w_cout_12_), .Y(_576_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_576_), .B(_580_), .Y(_0__48_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_574_), .C(_579_), .Y(_38__1_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_38__3_), .Y(_584_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_585_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_586_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_586_), .C(_585_), .Y(_587_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_581_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_582_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_581_), .B(_582_), .C(_38__3_), .Y(_583_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_583_), .B(_587_), .Y(_0__51_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_581_), .C(_586_), .Y(_37_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_38__1_), .Y(_591_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_592_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_593_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_593_), .C(_592_), .Y(_594_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_588_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_589_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_588_), .B(_589_), .C(_38__1_), .Y(_590_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_590_), .B(_594_), .Y(_0__49_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_588_), .C(_593_), .Y(_38__2_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_38__2_), .Y(_598_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_599_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_600_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_598_), .B(_600_), .C(_599_), .Y(_601_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_595_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_596_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_595_), .B(_596_), .C(_38__2_), .Y(_597_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_597_), .B(_601_), .Y(_0__50_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_598_), .B(_595_), .C(_600_), .Y(_38__3_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[48]), .Y(_602_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(_602_), .Y(_603_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .Y(_604_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[48]), .B(_604_), .Y(_605_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[49]), .Y(_606_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(_606_), .Y(_607_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .Y(_608_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[49]), .B(_608_), .Y(_609_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_603_), .B(_605_), .C(_607_), .D(_609_), .Y(_610_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_611_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_612_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_612_), .Y(_613_) );
XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_614_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_613_), .B(_614_), .Y(_615_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_615_), .Y(_39_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_37_), .Y(_616_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_39_), .Y(_617_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_616_), .C(_617_), .Y(w_cout_13_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(w_cout_13_), .Y(_621_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_622_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_623_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_623_), .C(_622_), .Y(_624_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_618_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_619_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_618_), .B(_619_), .C(w_cout_13_), .Y(_620_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_624_), .Y(_0__52_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_618_), .C(_623_), .Y(_41__1_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(_41__3_), .Y(_628_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_629_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_630_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_630_), .C(_629_), .Y(_631_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_625_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_626_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_625_), .B(_626_), .C(_41__3_), .Y(_627_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(_631_), .Y(_0__55_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_625_), .C(_630_), .Y(_40_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_41__1_), .Y(_635_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_636_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_637_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_637_), .C(_636_), .Y(_638_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_632_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_633_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_632_), .B(_633_), .C(_41__1_), .Y(_634_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_634_), .B(_638_), .Y(_0__53_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_632_), .C(_637_), .Y(_41__2_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_41__2_), .Y(_642_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_643_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_644_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_642_), .B(_644_), .C(_643_), .Y(_645_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_639_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_640_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_640_), .C(_41__2_), .Y(_641_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_641_), .B(_645_), .Y(_0__54_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_642_), .B(_639_), .C(_644_), .Y(_41__3_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[52]), .Y(_646_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(_646_), .Y(_647_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .Y(_648_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[52]), .B(_648_), .Y(_649_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[53]), .Y(_650_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(_650_), .Y(_651_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .Y(_652_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[53]), .B(_652_), .Y(_653_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_647_), .B(_649_), .C(_651_), .D(_653_), .Y(_654_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_655_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_656_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_656_), .Y(_657_) );
XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_658_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_657_), .B(_658_), .Y(_659_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_659_), .Y(_42_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(_40_), .Y(_660_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_42_), .Y(_661_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_660_), .C(_661_), .Y(w_cout_14_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(w_cout_14_), .Y(_665_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_666_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_667_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_665_), .B(_667_), .C(_666_), .Y(_668_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_662_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_663_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_663_), .C(w_cout_14_), .Y(_664_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_668_), .Y(_0__56_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_665_), .B(_662_), .C(_667_), .Y(_44__1_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(_44__3_), .Y(_672_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_673_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_674_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_672_), .B(_674_), .C(_673_), .Y(_675_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_669_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_670_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_669_), .B(_670_), .C(_44__3_), .Y(_671_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_671_), .B(_675_), .Y(_0__59_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_672_), .B(_669_), .C(_674_), .Y(_43_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_44__1_), .Y(_679_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_680_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_681_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_679_), .B(_681_), .C(_680_), .Y(_682_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_676_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_677_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_676_), .B(_677_), .C(_44__1_), .Y(_678_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_682_), .Y(_0__57_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_679_), .B(_676_), .C(_681_), .Y(_44__2_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_44__2_), .Y(_686_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_687_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_688_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_686_), .B(_688_), .C(_687_), .Y(_689_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_683_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_684_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_683_), .B(_684_), .C(_44__2_), .Y(_685_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_689_), .Y(_0__58_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_686_), .B(_683_), .C(_688_), .Y(_44__3_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[56]), .Y(_690_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(_690_), .Y(_691_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .Y(_692_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[56]), .B(_692_), .Y(_693_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[57]), .Y(_694_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(_694_), .Y(_695_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .Y(_696_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[57]), .B(_696_), .Y(_697_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_691_), .B(_693_), .C(_695_), .D(_697_), .Y(_698_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_699_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_700_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_700_), .Y(_701_) );
XOR2X1 XOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_702_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_701_), .B(_702_), .Y(_703_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_703_), .Y(_45_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(_704_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_45_), .Y(_705_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_704_), .C(_705_), .Y(cskip2_inst_cin) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_cin), .Y(_709_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_710_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_711_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_711_), .C(_710_), .Y(_712_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_706_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_707_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_707_), .C(cskip2_inst_cin), .Y(_708_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_708_), .B(_712_), .Y(cskip2_inst_rca0_fa0_o_sum) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_706_), .C(_711_), .Y(cskip2_inst_rca0_c) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_rca0_c), .Y(_716_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_717_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_718_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_716_), .B(_718_), .C(_717_), .Y(_719_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_713_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_714_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_714_), .C(cskip2_inst_rca0_c), .Y(_715_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(_719_), .Y(cskip2_inst_rca0_fa31_o_sum) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_716_), .B(_713_), .C(_718_), .Y(cskip2_inst_cout0) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[61]), .Y(_724_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[61]), .B(_724_), .Y(_725_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[61]), .Y(_726_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[61]), .B(_726_), .Y(_727_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[60]), .Y(_720_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[60]), .B(_720_), .Y(_721_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[60]), .Y(_722_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[60]), .B(_722_), .Y(_723_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(_727_), .C(_721_), .D(_723_), .Y(cskip2_inst_skip0_P) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_cout0), .Y(_728_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(cskip2_inst_skip0_P), .Y(_729_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_skip0_P), .B(_728_), .C(_729_), .Y(w_cout_16_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(w_cout_16_), .Y(cout) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_0__54_), .Y(sum[54]) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_0__55_), .Y(sum[55]) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_0__56_), .Y(sum[56]) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_0__57_), .Y(sum[57]) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(_0__58_), .Y(sum[58]) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(_0__59_), .Y(sum[59]) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_rca0_fa0_o_sum), .Y(sum[60]) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_rca0_fa31_o_sum), .Y(sum[61]) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_49_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_50_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_51_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_51_), .C(_50_), .Y(_52_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_46_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_47_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_47_), .C(gnd), .Y(_48_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_52_), .Y(_0__0_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_46_), .C(_51_), .Y(_2__1_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_2__3_), .Y(_56_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_57_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_58_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_58_), .C(_57_), .Y(_59_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_53_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_54_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_54_), .C(_2__3_), .Y(_55_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_59_), .Y(_0__3_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_53_), .C(_58_), .Y(_1_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(_2__1_), .Y(_63_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_64_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_65_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_65_), .C(_64_), .Y(_66_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_60_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_61_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_61_), .C(_2__1_), .Y(_62_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_66_), .Y(_0__1_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_60_), .C(_65_), .Y(_2__2_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_2__2_), .Y(_70_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_71_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_72_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_72_), .C(_71_), .Y(_73_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_67_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_68_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_68_), .C(_2__2_), .Y(_69_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_73_), .Y(_0__2_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_67_), .C(_72_), .Y(_2__3_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .Y(_74_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(_74_), .Y(_75_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .Y(_76_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .B(_76_), .Y(_77_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .Y(_78_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(_78_), .Y(_79_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .Y(_80_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .B(_80_), .Y(_81_) );
OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_77_), .C(_79_), .D(_81_), .Y(_82_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_83_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_84_) );
NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_84_), .Y(_85_) );
XOR2X1 XOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_86_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_86_), .Y(_87_) );
NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_87_), .Y(_3_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_88_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_3_), .Y(_89_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_88_), .C(_89_), .Y(w_cout_1_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .Y(_93_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_94_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_95_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_95_), .C(_94_), .Y(_96_) );
NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_90_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_91_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_91_), .C(w_cout_1_), .Y(_92_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_96_), .Y(_0__4_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_90_), .C(_95_), .Y(_5__1_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(_5__3_), .Y(_100_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_101_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_102_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_102_), .C(_101_), .Y(_103_) );
NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_97_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_98_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_98_), .C(_5__3_), .Y(_99_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_103_), .Y(_0__7_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_97_), .C(_102_), .Y(_4_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(_5__1_), .Y(_107_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_108_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_109_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_109_), .C(_108_), .Y(_110_) );
NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_104_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_105_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_105_), .C(_5__1_), .Y(_106_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_106_), .B(_110_), .Y(_0__5_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_104_), .C(_109_), .Y(_5__2_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(_5__2_), .Y(_114_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_115_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_116_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_116_), .C(_115_), .Y(_117_) );
NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_111_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_112_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_112_), .C(_5__2_), .Y(_113_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_117_), .Y(_0__6_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_111_), .C(_116_), .Y(_5__3_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[4]), .Y(_118_) );
NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(_118_), .Y(_119_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .Y(_120_) );
NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[4]), .B(_120_), .Y(_121_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[5]), .Y(_122_) );
NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(_122_), .Y(_123_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .Y(_124_) );
NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[5]), .B(_124_), .Y(_125_) );
OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_121_), .C(_123_), .D(_125_), .Y(_126_) );
NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_127_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_128_) );
NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_128_), .Y(_129_) );
XOR2X1 XOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_130_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_129_), .B(_130_), .Y(_131_) );
NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_131_), .Y(_6_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(_132_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_6_), .Y(_133_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_132_), .C(_133_), .Y(w_cout_2_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .Y(_137_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_138_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_139_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(_139_), .C(_138_), .Y(_140_) );
NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_134_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_135_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_135_), .C(w_cout_2_), .Y(_136_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_140_), .Y(_0__8_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(_134_), .C(_139_), .Y(_8__1_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(_8__3_), .Y(_144_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_145_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_146_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_146_), .C(_145_), .Y(_147_) );
NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_141_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_142_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_142_), .C(_8__3_), .Y(_143_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_147_), .Y(_0__11_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_141_), .C(_146_), .Y(_7_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(_8__1_), .Y(_151_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_152_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_153_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_153_), .C(_152_), .Y(_154_) );
NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_148_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_149_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_149_), .C(_8__1_), .Y(_150_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_154_), .Y(_0__9_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_148_), .C(_153_), .Y(_8__2_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(_8__2_), .Y(_158_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_159_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_160_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_160_), .C(_159_), .Y(_161_) );
NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_155_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_156_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_156_), .C(_8__2_), .Y(_157_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_161_), .Y(_0__10_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_155_), .C(_160_), .Y(_8__3_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[8]), .Y(_162_) );
NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(_162_), .Y(_163_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .Y(_164_) );
NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[8]), .B(_164_), .Y(_165_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[9]), .Y(_166_) );
NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(_166_), .Y(_167_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .Y(_168_) );
NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[9]), .B(_168_), .Y(_169_) );
OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_165_), .C(_167_), .D(_169_), .Y(_170_) );
NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_171_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_172_) );
NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_172_), .Y(_173_) );
XOR2X1 XOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_174_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(_174_), .Y(_175_) );
NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_175_), .Y(_9_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_176_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_9_), .Y(_177_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_176_), .C(_177_), .Y(w_cout_3_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .Y(_181_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_182_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_183_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_183_), .C(_182_), .Y(_184_) );
NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_178_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_179_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_179_), .C(w_cout_3_), .Y(_180_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_184_), .Y(_0__12_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_178_), .C(_183_), .Y(_11__1_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(_11__3_), .Y(_188_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_189_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_190_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_190_), .C(_189_), .Y(_191_) );
NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_185_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_186_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_186_), .C(_11__3_), .Y(_187_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(_191_), .Y(_0__15_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_185_), .C(_190_), .Y(_10_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(_11__1_), .Y(_195_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_196_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_197_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_197_), .C(_196_), .Y(_198_) );
NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_192_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_193_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(_193_), .C(_11__1_), .Y(_194_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_198_), .Y(_0__13_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_192_), .C(_197_), .Y(_11__2_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(_11__2_), .Y(_202_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_203_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_204_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_204_), .C(_203_), .Y(_205_) );
NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_199_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_200_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_200_), .C(_11__2_), .Y(_201_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_205_), .Y(_0__14_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_199_), .C(_204_), .Y(_11__3_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[12]), .Y(_206_) );
NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(_206_), .Y(_207_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .Y(_208_) );
NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[12]), .B(_208_), .Y(_209_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[13]), .Y(_210_) );
NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(_210_), .Y(_211_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .Y(_212_) );
NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[13]), .B(_212_), .Y(_213_) );
OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_209_), .C(_211_), .D(_213_), .Y(_214_) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_rca0_fa0_o_sum), .Y(_0__60_) );
BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_rca0_fa31_o_sum), .Y(_0__61_) );
BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_67 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_cin), .Y(w_cout_15_) );
endmodule
