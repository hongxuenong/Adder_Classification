magic
tech scmos
magscale 1 2
timestamp 1586568500
<< metal1 >>
rect 616 1606 622 1614
rect 630 1606 636 1614
rect 644 1606 650 1614
rect 658 1606 664 1614
rect 749 1537 764 1543
rect 813 1517 828 1523
rect 164 1497 179 1503
rect 189 1497 204 1503
rect 493 1497 563 1503
rect 861 1503 867 1523
rect 861 1497 876 1503
rect 1213 1497 1251 1503
rect 1261 1497 1299 1503
rect 1485 1497 1500 1503
rect 1581 1497 1667 1503
rect 205 1477 220 1483
rect 205 1457 211 1477
rect 333 1477 348 1483
rect 333 1457 339 1477
rect 644 1477 668 1483
rect 676 1477 684 1483
rect 692 1477 723 1483
rect 893 1477 908 1483
rect 1037 1477 1059 1483
rect 1133 1477 1155 1483
rect 1165 1477 1203 1483
rect 660 1457 707 1463
rect 1197 1457 1203 1477
rect 1581 1477 1587 1497
rect 1940 1497 1955 1503
rect 2141 1503 2147 1523
rect 2109 1497 2147 1503
rect 2173 1497 2211 1503
rect 1725 1477 1747 1483
rect 1965 1477 1980 1483
rect 2013 1483 2019 1496
rect 2013 1477 2051 1483
rect 2020 1457 2035 1463
rect 148 1436 150 1444
rect 637 1437 684 1443
rect 1576 1406 1582 1414
rect 1590 1406 1596 1414
rect 1604 1406 1610 1414
rect 1618 1406 1624 1414
rect 973 1363 979 1383
rect 1274 1376 1276 1384
rect 973 1357 995 1363
rect 1508 1357 1523 1363
rect 52 1317 83 1323
rect 237 1323 243 1343
rect 733 1337 771 1343
rect 813 1337 835 1343
rect 1005 1337 1020 1343
rect 1197 1343 1203 1356
rect 1181 1337 1203 1343
rect 212 1317 243 1323
rect 493 1317 531 1323
rect 1389 1323 1395 1343
rect 1501 1337 1516 1343
rect 1389 1317 1420 1323
rect 1501 1317 1507 1337
rect 1524 1337 1539 1343
rect 1741 1343 1747 1363
rect 1709 1337 1747 1343
rect 1757 1317 1795 1323
rect 1805 1317 1843 1323
rect 1988 1317 2003 1323
rect 2212 1317 2227 1323
rect 100 1297 115 1303
rect 1677 1297 1692 1303
rect 1260 1284 1268 1288
rect 973 1277 988 1283
rect 1492 1276 1494 1284
rect 1565 1277 1667 1283
rect 616 1206 622 1214
rect 630 1206 636 1214
rect 644 1206 650 1214
rect 658 1206 664 1214
rect 781 1117 819 1123
rect 1037 1117 1052 1123
rect 1085 1117 1100 1123
rect 1549 1117 1612 1123
rect 1732 1116 1740 1124
rect 589 1097 675 1103
rect 973 1097 1011 1103
rect 1117 1097 1155 1103
rect 1165 1097 1203 1103
rect 1716 1097 1731 1103
rect 1940 1097 1971 1103
rect 2045 1103 2051 1123
rect 2045 1097 2083 1103
rect 460 1092 468 1096
rect 61 1077 76 1083
rect 93 1077 124 1083
rect 173 1077 195 1083
rect 253 1077 275 1083
rect 445 1077 467 1083
rect 445 1057 451 1077
rect 765 1077 787 1083
rect 909 1077 924 1083
rect 1037 1077 1059 1083
rect 1069 1077 1107 1083
rect 1101 1057 1107 1077
rect 1293 1077 1308 1083
rect 1396 1077 1427 1083
rect 1556 1077 1619 1083
rect 1693 1077 1715 1083
rect 1869 1077 1900 1083
rect 1933 1077 1948 1083
rect 2228 1057 2236 1063
rect 538 1036 540 1044
rect 1380 1036 1382 1044
rect 1540 1036 1542 1044
rect 1576 1006 1582 1014
rect 1590 1006 1596 1014
rect 1604 1006 1610 1014
rect 1618 1006 1624 1014
rect 282 976 284 984
rect 708 976 710 984
rect 1204 976 1206 984
rect 2237 957 2252 963
rect 509 937 547 943
rect 621 937 691 943
rect 733 937 764 943
rect 925 937 956 943
rect 996 937 1011 943
rect 1117 937 1139 943
rect 1149 937 1187 943
rect 1309 937 1331 943
rect 1629 937 1667 943
rect 1876 937 1891 943
rect 1965 937 1996 943
rect 420 917 435 923
rect 493 917 508 923
rect 541 917 595 923
rect 1053 917 1091 923
rect 1236 917 1251 923
rect 1332 917 1347 923
rect 1533 917 1635 923
rect 1668 917 1683 923
rect 452 897 467 903
rect 756 897 771 903
rect 1437 897 1452 903
rect 1709 897 1724 903
rect 1741 897 1763 903
rect 2077 897 2092 903
rect 2109 897 2131 903
rect 716 884 724 888
rect 1116 877 1139 883
rect 1133 857 1139 877
rect 2100 877 2115 883
rect 1530 836 1532 844
rect 1684 836 1686 844
rect 2052 836 2054 844
rect 616 806 622 814
rect 630 806 636 814
rect 644 806 650 814
rect 658 806 664 814
rect 61 737 76 743
rect 1021 737 1036 743
rect 500 717 515 723
rect 557 717 595 723
rect 1076 717 1091 723
rect 1524 716 1532 724
rect 589 697 659 703
rect 340 677 355 683
rect 388 677 419 683
rect 653 677 659 697
rect 1101 697 1116 703
rect 1533 697 1619 703
rect 1821 703 1827 723
rect 1837 717 1875 723
rect 2084 716 2092 724
rect 1789 697 1827 703
rect 1901 697 1939 703
rect 1956 697 1971 703
rect 2068 697 2083 703
rect 1245 677 1267 683
rect 1325 677 1347 683
rect 1396 677 1427 683
rect 2221 677 2236 683
rect 1476 636 1478 644
rect 1576 606 1582 614
rect 1590 606 1596 614
rect 1604 606 1610 614
rect 1618 606 1624 614
rect 893 557 908 563
rect 404 537 419 543
rect 797 537 828 543
rect 861 537 876 543
rect 1172 537 1187 543
rect 1229 537 1267 543
rect 1565 537 1628 543
rect 1949 537 1971 543
rect 2013 537 2051 543
rect 2093 537 2108 543
rect 269 517 307 523
rect 461 517 499 523
rect 573 517 588 523
rect 1485 517 1523 523
rect 109 497 147 503
rect 228 497 236 503
rect 500 496 508 504
rect 1485 497 1491 517
rect 2045 517 2076 523
rect 2180 477 2211 483
rect 730 436 732 444
rect 1284 436 1286 444
rect 616 406 622 414
rect 630 406 636 414
rect 644 406 650 414
rect 658 406 664 414
rect 1140 376 1142 384
rect 2180 337 2195 343
rect 1292 332 1300 336
rect 2092 332 2100 336
rect 45 297 60 303
rect 93 303 99 323
rect 628 317 691 323
rect 765 317 787 323
rect 932 316 940 324
rect 1037 317 1059 323
rect 1549 317 1596 323
rect 1620 317 1635 323
rect 1052 304 1060 308
rect 93 297 131 303
rect 189 297 227 303
rect 621 297 707 303
rect 141 277 163 283
rect 269 277 284 283
rect 349 277 371 283
rect 573 277 611 283
rect 621 277 627 297
rect 1197 297 1212 303
rect 573 257 579 277
rect 756 277 771 283
rect 1533 277 1555 283
rect 1684 277 1715 283
rect 1917 283 1923 303
rect 2077 303 2083 323
rect 2013 297 2051 303
rect 2077 297 2092 303
rect 1892 277 1923 283
rect 1956 277 1971 283
rect 2221 277 2236 283
rect 84 236 86 244
rect 749 237 755 263
rect 1565 257 1612 263
rect 1901 257 1916 263
rect 2237 257 2252 263
rect 1386 236 1388 244
rect 2106 236 2108 244
rect 1576 206 1582 214
rect 1590 206 1596 214
rect 1604 206 1610 214
rect 1618 206 1624 214
rect 141 143 147 163
rect 1172 157 1196 163
rect 141 137 179 143
rect 301 137 332 143
rect 580 137 611 143
rect 1117 137 1132 143
rect 1229 143 1235 163
rect 1220 137 1235 143
rect 1732 137 1740 143
rect 1780 137 1811 143
rect 1116 124 1124 128
rect 45 117 83 123
rect 93 117 131 123
rect 484 117 499 123
rect 804 117 835 123
rect 1012 117 1027 123
rect 1165 117 1180 123
rect 1309 117 1324 123
rect 1380 117 1395 123
rect 1565 117 1651 123
rect 1869 117 1900 123
rect 2196 117 2211 123
rect 196 97 211 103
rect 349 97 387 103
rect 797 97 803 116
rect 1901 97 1907 116
rect 2068 97 2083 103
rect 221 77 275 83
rect 1837 77 1852 83
rect 2237 77 2252 83
rect 616 6 622 14
rect 630 6 636 14
rect 644 6 650 14
rect 658 6 664 14
<< m2contact >>
rect 622 1606 630 1614
rect 636 1606 644 1614
rect 650 1606 658 1614
rect 588 1576 596 1584
rect 1324 1576 1332 1584
rect 1532 1576 1540 1584
rect 1868 1576 1876 1584
rect 428 1556 436 1564
rect 956 1556 964 1564
rect 1820 1556 1828 1564
rect 284 1536 292 1544
rect 412 1536 420 1544
rect 764 1536 772 1544
rect 940 1536 948 1544
rect 1836 1536 1844 1544
rect 2076 1536 2084 1544
rect 156 1516 164 1524
rect 380 1516 388 1524
rect 444 1516 452 1524
rect 508 1516 516 1524
rect 636 1516 644 1524
rect 828 1516 836 1524
rect 44 1496 52 1504
rect 156 1496 164 1504
rect 204 1496 212 1504
rect 236 1496 244 1504
rect 428 1496 436 1504
rect 780 1496 788 1504
rect 844 1496 852 1504
rect 972 1516 980 1524
rect 988 1516 996 1524
rect 1052 1516 1060 1524
rect 1132 1516 1140 1524
rect 1180 1516 1188 1524
rect 1276 1516 1284 1524
rect 1436 1516 1444 1524
rect 1548 1516 1556 1524
rect 1644 1516 1652 1524
rect 1724 1516 1732 1524
rect 1788 1516 1796 1524
rect 1804 1516 1812 1524
rect 1932 1516 1940 1524
rect 2124 1516 2132 1524
rect 876 1496 884 1504
rect 956 1496 964 1504
rect 1020 1496 1028 1504
rect 1100 1496 1108 1504
rect 1356 1496 1364 1504
rect 1500 1496 1508 1504
rect 1564 1496 1572 1504
rect 76 1476 84 1484
rect 124 1476 132 1484
rect 60 1456 68 1464
rect 220 1476 228 1484
rect 316 1476 324 1484
rect 348 1476 356 1484
rect 540 1476 548 1484
rect 604 1476 612 1484
rect 636 1476 644 1484
rect 668 1476 676 1484
rect 684 1476 692 1484
rect 764 1476 772 1484
rect 828 1476 836 1484
rect 908 1476 916 1484
rect 1084 1476 1092 1484
rect 652 1456 660 1464
rect 908 1456 916 1464
rect 1068 1456 1076 1464
rect 1228 1476 1236 1484
rect 1340 1476 1348 1484
rect 1404 1476 1412 1484
rect 1676 1496 1684 1504
rect 1756 1496 1764 1504
rect 1820 1496 1828 1504
rect 1900 1496 1908 1504
rect 1932 1496 1940 1504
rect 2012 1496 2020 1504
rect 1692 1476 1700 1484
rect 1916 1476 1924 1484
rect 1980 1476 1988 1484
rect 1996 1476 2004 1484
rect 2092 1476 2100 1484
rect 2188 1476 2196 1484
rect 1708 1456 1716 1464
rect 1980 1456 1988 1464
rect 2012 1456 2020 1464
rect 2220 1456 2228 1464
rect 108 1436 116 1444
rect 140 1436 148 1444
rect 268 1436 276 1444
rect 380 1436 388 1444
rect 684 1436 692 1444
rect 988 1436 996 1444
rect 1388 1436 1396 1444
rect 1436 1436 1444 1444
rect 1788 1436 1796 1444
rect 2140 1436 2148 1444
rect 1582 1406 1590 1414
rect 1596 1406 1604 1414
rect 1610 1406 1618 1414
rect 2092 1396 2100 1404
rect 284 1356 292 1364
rect 316 1356 324 1364
rect 348 1356 356 1364
rect 364 1356 372 1364
rect 572 1356 580 1364
rect 588 1356 596 1364
rect 716 1356 724 1364
rect 924 1356 932 1364
rect 940 1356 948 1364
rect 1068 1376 1076 1384
rect 1276 1376 1284 1384
rect 1340 1376 1348 1384
rect 1868 1376 1876 1384
rect 1980 1376 1988 1384
rect 2204 1376 2212 1384
rect 1196 1356 1204 1364
rect 1308 1356 1316 1364
rect 1324 1356 1332 1364
rect 1468 1356 1476 1364
rect 1500 1356 1508 1364
rect 92 1336 100 1344
rect 220 1336 228 1344
rect 44 1316 52 1324
rect 140 1316 148 1324
rect 188 1316 196 1324
rect 204 1316 212 1324
rect 300 1336 308 1344
rect 428 1336 436 1344
rect 444 1336 452 1344
rect 508 1336 516 1344
rect 540 1336 548 1344
rect 652 1336 660 1344
rect 908 1336 916 1344
rect 1020 1336 1028 1344
rect 1212 1336 1220 1344
rect 1244 1336 1252 1344
rect 1292 1336 1300 1344
rect 252 1316 260 1324
rect 332 1316 340 1324
rect 396 1316 404 1324
rect 412 1316 420 1324
rect 460 1316 468 1324
rect 668 1316 676 1324
rect 748 1316 756 1324
rect 780 1316 788 1324
rect 972 1316 980 1324
rect 1036 1316 1044 1324
rect 1100 1316 1108 1324
rect 1372 1316 1380 1324
rect 1404 1336 1412 1344
rect 1420 1316 1428 1324
rect 1436 1316 1444 1324
rect 1516 1336 1524 1344
rect 1692 1336 1700 1344
rect 2092 1356 2100 1364
rect 1772 1336 1780 1344
rect 1932 1336 1940 1344
rect 1948 1336 1956 1344
rect 2044 1336 2052 1344
rect 2124 1336 2132 1344
rect 2156 1336 2164 1344
rect 2172 1336 2180 1344
rect 1644 1316 1652 1324
rect 1900 1316 1908 1324
rect 1916 1316 1924 1324
rect 1980 1316 1988 1324
rect 2028 1316 2036 1324
rect 2060 1316 2068 1324
rect 2076 1316 2084 1324
rect 2140 1316 2148 1324
rect 2204 1316 2212 1324
rect 60 1296 68 1304
rect 92 1296 100 1304
rect 156 1296 164 1304
rect 172 1296 180 1304
rect 284 1296 292 1304
rect 380 1296 388 1304
rect 556 1296 564 1304
rect 700 1296 708 1304
rect 812 1296 820 1304
rect 860 1296 868 1304
rect 1068 1296 1076 1304
rect 1084 1296 1092 1304
rect 1148 1296 1156 1304
rect 1164 1296 1172 1304
rect 1340 1296 1348 1304
rect 1452 1296 1460 1304
rect 1628 1296 1636 1304
rect 1692 1296 1700 1304
rect 1724 1296 1732 1304
rect 1820 1296 1828 1304
rect 1980 1296 1988 1304
rect 2108 1296 2116 1304
rect 2204 1296 2212 1304
rect 12 1276 20 1284
rect 124 1276 132 1284
rect 844 1276 852 1284
rect 988 1276 996 1284
rect 1116 1276 1124 1284
rect 1260 1276 1268 1284
rect 1484 1276 1492 1284
rect 1884 1276 1892 1284
rect 2252 1276 2260 1284
rect 748 1236 756 1244
rect 876 1236 884 1244
rect 1100 1236 1108 1244
rect 1884 1236 1892 1244
rect 622 1206 630 1214
rect 636 1206 644 1214
rect 650 1206 658 1214
rect 860 1176 868 1184
rect 1228 1176 1236 1184
rect 1484 1176 1492 1184
rect 1820 1176 1828 1184
rect 2156 1176 2164 1184
rect 348 1156 356 1164
rect 1676 1156 1684 1164
rect 364 1136 372 1144
rect 396 1136 404 1144
rect 844 1136 852 1144
rect 1804 1136 1812 1144
rect 1836 1136 1844 1144
rect 2140 1136 2148 1144
rect 2172 1136 2180 1144
rect 172 1116 180 1124
rect 220 1116 228 1124
rect 252 1116 260 1124
rect 316 1116 324 1124
rect 332 1116 340 1124
rect 524 1116 532 1124
rect 700 1116 708 1124
rect 716 1116 724 1124
rect 876 1116 884 1124
rect 1052 1116 1060 1124
rect 1100 1116 1108 1124
rect 1180 1116 1188 1124
rect 1388 1116 1396 1124
rect 1500 1116 1508 1124
rect 1612 1116 1620 1124
rect 1692 1116 1700 1124
rect 1724 1116 1732 1124
rect 1756 1116 1764 1124
rect 1772 1116 1780 1124
rect 1900 1116 1908 1124
rect 1916 1116 1924 1124
rect 12 1096 20 1104
rect 108 1096 116 1104
rect 140 1096 148 1104
rect 284 1096 292 1104
rect 348 1096 356 1104
rect 460 1096 468 1104
rect 748 1096 756 1104
rect 828 1096 836 1104
rect 940 1096 948 1104
rect 1276 1096 1284 1104
rect 1340 1096 1348 1104
rect 1628 1096 1636 1104
rect 1708 1096 1716 1104
rect 1788 1096 1796 1104
rect 1932 1096 1940 1104
rect 1980 1096 1988 1104
rect 2012 1096 2020 1104
rect 2060 1116 2068 1124
rect 2108 1116 2116 1124
rect 2124 1096 2132 1104
rect 44 1080 52 1088
rect 76 1076 84 1084
rect 124 1076 132 1084
rect 428 1076 436 1084
rect 476 1080 484 1088
rect 76 1056 84 1064
rect 204 1056 212 1064
rect 236 1056 244 1064
rect 316 1056 324 1064
rect 556 1076 564 1084
rect 652 1076 660 1084
rect 924 1076 932 1084
rect 988 1076 996 1084
rect 572 1056 580 1064
rect 796 1056 804 1064
rect 1132 1076 1140 1084
rect 1308 1076 1316 1084
rect 1356 1076 1364 1084
rect 1388 1076 1396 1084
rect 1468 1076 1476 1084
rect 1516 1076 1524 1084
rect 1548 1076 1556 1084
rect 1900 1076 1908 1084
rect 1948 1076 1956 1084
rect 1996 1076 2004 1084
rect 2076 1076 2084 1084
rect 2092 1076 2100 1084
rect 2204 1076 2212 1084
rect 1308 1056 1316 1064
rect 1404 1056 1412 1064
rect 1676 1056 1684 1064
rect 1884 1056 1892 1064
rect 1948 1056 1956 1064
rect 2220 1056 2228 1064
rect 2236 1056 2244 1064
rect 508 1036 516 1044
rect 540 1036 548 1044
rect 700 1036 708 1044
rect 716 1036 724 1044
rect 876 1036 884 1044
rect 1052 1036 1060 1044
rect 1244 1036 1252 1044
rect 1324 1036 1332 1044
rect 1372 1036 1380 1044
rect 1452 1036 1460 1044
rect 1532 1036 1540 1044
rect 1660 1036 1668 1044
rect 2044 1036 2052 1044
rect 1582 1006 1590 1014
rect 1596 1006 1604 1014
rect 1610 1006 1618 1014
rect 1996 996 2004 1004
rect 284 976 292 984
rect 700 976 708 984
rect 1196 976 1204 984
rect 1484 976 1492 984
rect 2012 976 2020 984
rect 140 956 148 964
rect 204 956 212 964
rect 396 956 404 964
rect 444 956 452 964
rect 460 956 468 964
rect 556 956 564 964
rect 748 956 756 964
rect 940 956 948 964
rect 988 956 996 964
rect 1292 956 1300 964
rect 1612 956 1620 964
rect 1724 956 1732 964
rect 1868 956 1876 964
rect 1980 956 1988 964
rect 1996 956 2004 964
rect 2092 956 2100 964
rect 2252 956 2260 964
rect 60 936 68 944
rect 92 936 100 944
rect 156 936 164 944
rect 172 936 180 944
rect 220 936 228 944
rect 300 936 308 944
rect 412 936 420 944
rect 572 936 580 944
rect 764 936 772 944
rect 796 936 804 944
rect 956 936 964 944
rect 972 936 980 944
rect 988 936 996 944
rect 1068 936 1076 944
rect 1276 936 1284 944
rect 1452 936 1460 944
rect 1548 936 1556 944
rect 1740 936 1748 944
rect 1852 936 1860 944
rect 1868 936 1876 944
rect 1996 936 2004 944
rect 2028 936 2036 944
rect 2220 936 2228 944
rect 44 916 52 924
rect 76 916 84 924
rect 348 916 356 924
rect 412 916 420 924
rect 508 916 516 924
rect 524 916 532 924
rect 780 916 788 924
rect 844 916 852 924
rect 956 916 964 924
rect 1020 916 1028 924
rect 1228 916 1236 924
rect 1260 916 1268 924
rect 1324 916 1332 924
rect 1356 916 1364 924
rect 1404 916 1412 924
rect 1644 916 1652 924
rect 1660 916 1668 924
rect 1772 916 1780 924
rect 1900 916 1908 924
rect 1932 916 1940 924
rect 1948 916 1956 924
rect 2044 916 2052 924
rect 2140 916 2148 924
rect 108 896 116 904
rect 124 896 132 904
rect 188 896 196 904
rect 268 896 276 904
rect 364 896 372 904
rect 380 896 388 904
rect 444 896 452 904
rect 620 896 628 904
rect 748 896 756 904
rect 812 896 820 904
rect 828 896 836 904
rect 876 896 884 904
rect 1164 896 1172 904
rect 1212 896 1220 904
rect 1228 896 1236 904
rect 1308 896 1316 904
rect 1372 896 1380 904
rect 1388 896 1396 904
rect 1452 896 1460 904
rect 1484 896 1492 904
rect 1500 896 1508 904
rect 1724 896 1732 904
rect 2092 896 2100 904
rect 12 876 20 884
rect 252 876 260 884
rect 332 876 340 884
rect 716 876 724 884
rect 860 876 868 884
rect 892 876 900 884
rect 348 856 356 864
rect 1420 876 1428 884
rect 1788 876 1796 884
rect 1820 876 1828 884
rect 2092 876 2100 884
rect 2156 876 2164 884
rect 2188 876 2196 884
rect 1532 836 1540 844
rect 1676 836 1684 844
rect 1804 836 1812 844
rect 2044 836 2052 844
rect 2140 836 2148 844
rect 622 806 630 814
rect 636 806 644 814
rect 650 806 658 814
rect 956 776 964 784
rect 2172 776 2180 784
rect 156 756 164 764
rect 764 756 772 764
rect 828 756 836 764
rect 1164 756 1172 764
rect 76 736 84 744
rect 140 736 148 744
rect 444 736 452 744
rect 524 736 532 744
rect 812 736 820 744
rect 956 736 964 744
rect 1036 736 1044 744
rect 1148 736 1156 744
rect 1996 736 2004 744
rect 108 716 116 724
rect 172 716 180 724
rect 188 716 196 724
rect 236 716 244 724
rect 380 716 388 724
rect 460 716 468 724
rect 492 716 500 724
rect 700 716 708 724
rect 716 716 724 724
rect 780 716 788 724
rect 844 716 852 724
rect 860 716 868 724
rect 1068 716 1076 724
rect 1180 716 1188 724
rect 1196 716 1204 724
rect 1260 716 1268 724
rect 1292 716 1300 724
rect 1340 716 1348 724
rect 1484 716 1492 724
rect 1500 716 1508 724
rect 1532 716 1540 724
rect 1724 716 1732 724
rect 1804 716 1812 724
rect 92 696 100 704
rect 156 696 164 704
rect 252 696 260 704
rect 268 696 276 704
rect 300 696 308 704
rect 316 696 324 704
rect 364 696 372 704
rect 540 696 548 704
rect 28 676 36 684
rect 76 676 84 684
rect 220 676 228 684
rect 284 676 292 684
rect 332 676 340 684
rect 380 676 388 684
rect 492 676 500 684
rect 668 696 676 704
rect 684 696 692 704
rect 828 696 836 704
rect 924 696 932 704
rect 1116 696 1124 704
rect 1164 696 1172 704
rect 1228 696 1236 704
rect 1372 696 1380 704
rect 1404 696 1412 704
rect 1644 696 1652 704
rect 1676 696 1684 704
rect 2012 716 2020 724
rect 2076 716 2084 724
rect 2108 716 2116 724
rect 2156 716 2164 724
rect 1884 696 1892 704
rect 1948 696 1956 704
rect 2060 696 2068 704
rect 2204 696 2212 704
rect 748 676 756 684
rect 876 676 884 684
rect 892 676 900 684
rect 908 676 916 684
rect 940 676 948 684
rect 988 676 996 684
rect 1036 676 1044 684
rect 1116 676 1124 684
rect 1388 676 1396 684
rect 1452 676 1460 684
rect 1548 676 1556 684
rect 1660 676 1668 684
rect 1692 676 1700 684
rect 1756 676 1764 684
rect 1772 676 1780 684
rect 1852 676 1860 684
rect 1916 676 1924 684
rect 2044 676 2052 684
rect 2060 676 2068 684
rect 2124 676 2132 684
rect 2236 676 2244 684
rect 12 656 20 664
rect 332 656 340 664
rect 396 656 404 664
rect 572 656 580 664
rect 764 656 772 664
rect 972 656 980 664
rect 1276 656 1284 664
rect 1436 656 1444 664
rect 1708 656 1716 664
rect 1948 656 1956 664
rect 2028 656 2036 664
rect 188 636 196 644
rect 460 636 468 644
rect 716 636 724 644
rect 1068 636 1076 644
rect 1196 636 1204 644
rect 1292 636 1300 644
rect 1468 636 1476 644
rect 1724 636 1732 644
rect 2156 636 2164 644
rect 1582 606 1590 614
rect 1596 606 1604 614
rect 1610 606 1618 614
rect 204 576 212 584
rect 236 576 244 584
rect 764 576 772 584
rect 828 576 836 584
rect 972 576 980 584
rect 1324 576 1332 584
rect 1388 576 1396 584
rect 172 556 180 564
rect 188 556 196 564
rect 220 556 228 564
rect 380 556 388 564
rect 396 556 404 564
rect 812 556 820 564
rect 876 556 884 564
rect 908 556 916 564
rect 988 556 996 564
rect 1196 556 1204 564
rect 1212 556 1220 564
rect 1548 556 1556 564
rect 1804 556 1812 564
rect 1820 556 1828 564
rect 1932 556 1940 564
rect 2060 556 2068 564
rect 2076 556 2084 564
rect 60 536 68 544
rect 124 536 132 544
rect 284 536 292 544
rect 332 532 340 540
rect 348 536 356 544
rect 396 536 404 544
rect 428 532 436 540
rect 476 536 484 544
rect 588 536 596 544
rect 748 536 756 544
rect 828 536 836 544
rect 876 536 884 544
rect 924 536 932 544
rect 1004 536 1012 544
rect 1164 536 1172 544
rect 1372 536 1380 544
rect 1436 536 1444 544
rect 1452 536 1460 544
rect 1532 536 1540 544
rect 1628 536 1636 544
rect 1788 536 1796 544
rect 1852 536 1860 544
rect 2108 536 2116 544
rect 44 516 52 524
rect 76 516 84 524
rect 92 516 100 524
rect 364 516 372 524
rect 588 516 596 524
rect 604 516 612 524
rect 620 516 628 524
rect 732 516 740 524
rect 908 516 916 524
rect 940 516 948 524
rect 1084 516 1092 524
rect 1132 516 1140 524
rect 1148 516 1156 524
rect 1244 516 1252 524
rect 1276 516 1284 524
rect 1356 516 1364 524
rect 1420 516 1428 524
rect 156 496 164 504
rect 220 496 228 504
rect 236 496 244 504
rect 492 496 500 504
rect 524 496 532 504
rect 636 496 644 504
rect 700 496 708 504
rect 828 496 836 504
rect 1100 496 1108 504
rect 1116 496 1124 504
rect 1228 496 1236 504
rect 1308 496 1316 504
rect 1644 516 1652 524
rect 1660 516 1668 524
rect 1708 516 1716 524
rect 1868 516 1876 524
rect 1996 516 2004 524
rect 2028 516 2036 524
rect 2076 516 2084 524
rect 2124 516 2132 524
rect 2140 516 2148 524
rect 2188 516 2196 524
rect 1500 496 1508 504
rect 1676 496 1684 504
rect 1692 496 1700 504
rect 1900 496 1908 504
rect 1916 496 1924 504
rect 1964 496 1972 504
rect 2156 496 2164 504
rect 2172 496 2180 504
rect 12 476 20 484
rect 1036 476 1044 484
rect 1068 476 1076 484
rect 1724 476 1732 484
rect 1756 476 1764 484
rect 2172 476 2180 484
rect 1708 456 1716 464
rect 2188 456 2196 464
rect 540 436 548 444
rect 732 436 740 444
rect 1084 436 1092 444
rect 1276 436 1284 444
rect 1468 436 1476 444
rect 1836 436 1844 444
rect 622 406 630 414
rect 636 406 644 414
rect 650 406 658 414
rect 556 376 564 384
rect 1132 376 1140 384
rect 2156 376 2164 384
rect 444 356 452 364
rect 492 356 500 364
rect 796 356 804 364
rect 1068 356 1076 364
rect 1804 356 1812 364
rect 1852 356 1860 364
rect 460 336 468 344
rect 812 336 820 344
rect 844 336 852 344
rect 1084 336 1092 344
rect 1292 336 1300 344
rect 1756 336 1764 344
rect 1820 336 1828 344
rect 2076 336 2084 344
rect 2092 336 2100 344
rect 2172 336 2180 344
rect 60 296 68 304
rect 108 316 116 324
rect 156 316 164 324
rect 348 316 356 324
rect 412 316 420 324
rect 428 316 436 324
rect 588 316 596 324
rect 620 316 628 324
rect 908 316 916 324
rect 940 316 948 324
rect 1004 316 1012 324
rect 1164 316 1172 324
rect 1212 316 1220 324
rect 1356 316 1364 324
rect 1372 316 1380 324
rect 1468 316 1476 324
rect 1484 316 1492 324
rect 1596 316 1604 324
rect 1612 316 1620 324
rect 1772 316 1780 324
rect 1788 316 1796 324
rect 300 296 308 304
rect 316 296 324 304
rect 380 296 388 304
rect 396 296 404 304
rect 444 296 452 304
rect 60 276 68 284
rect 204 276 212 284
rect 252 280 260 288
rect 284 276 292 284
rect 524 276 532 284
rect 716 296 724 304
rect 796 296 804 304
rect 940 296 948 304
rect 1052 296 1060 304
rect 1068 296 1076 304
rect 1132 296 1140 304
rect 1212 296 1220 304
rect 1324 296 1332 304
rect 1436 296 1444 304
rect 1516 296 1524 304
rect 1660 296 1668 304
rect 1692 296 1700 304
rect 1804 296 1812 304
rect 284 256 292 264
rect 332 256 340 264
rect 540 256 548 264
rect 732 276 740 284
rect 748 276 756 284
rect 876 276 884 284
rect 956 276 964 284
rect 972 276 980 284
rect 1116 276 1124 284
rect 1244 276 1252 284
rect 1260 276 1268 284
rect 1308 276 1316 284
rect 1404 276 1412 284
rect 1420 276 1428 284
rect 1484 276 1492 284
rect 1644 276 1652 284
rect 1676 276 1684 284
rect 1740 276 1748 284
rect 1884 276 1892 284
rect 1980 296 1988 304
rect 2140 316 2148 324
rect 2092 296 2100 304
rect 1948 276 1956 284
rect 2028 276 2036 284
rect 2060 276 2068 284
rect 2124 276 2132 284
rect 2172 276 2180 284
rect 2236 276 2244 284
rect 76 236 84 244
rect 620 236 628 244
rect 892 256 900 264
rect 1020 256 1028 264
rect 1180 256 1188 264
rect 1228 256 1236 264
rect 1612 256 1620 264
rect 1724 256 1732 264
rect 1916 256 1924 264
rect 1948 256 1956 264
rect 2252 256 2260 264
rect 860 236 868 244
rect 1004 236 1012 244
rect 1292 236 1300 244
rect 1356 236 1364 244
rect 1388 236 1396 244
rect 1468 236 1476 244
rect 1932 236 1940 244
rect 2108 236 2116 244
rect 1020 216 1028 224
rect 1582 206 1590 214
rect 1596 206 1604 214
rect 1610 206 1618 214
rect 380 176 388 184
rect 444 176 452 184
rect 524 176 532 184
rect 908 176 916 184
rect 1068 176 1076 184
rect 1148 176 1156 184
rect 1276 176 1284 184
rect 1676 176 1684 184
rect 1772 176 1780 184
rect 108 136 116 144
rect 316 156 324 164
rect 508 156 516 164
rect 588 156 596 164
rect 876 156 884 164
rect 892 156 900 164
rect 1132 156 1140 164
rect 1164 156 1172 164
rect 188 136 196 144
rect 332 136 340 144
rect 364 136 372 144
rect 428 136 436 144
rect 476 136 484 144
rect 572 136 580 144
rect 684 136 692 144
rect 748 136 756 144
rect 844 136 852 144
rect 956 136 964 144
rect 1132 136 1140 144
rect 1212 136 1220 144
rect 1292 156 1300 164
rect 1660 156 1668 164
rect 1788 156 1796 164
rect 1900 156 1908 164
rect 2044 156 2052 164
rect 2092 156 2100 164
rect 2108 156 2116 164
rect 1244 136 1252 144
rect 1372 136 1380 144
rect 1532 136 1540 144
rect 1580 136 1588 144
rect 1724 136 1732 144
rect 1740 136 1748 144
rect 1772 136 1780 144
rect 1852 136 1860 144
rect 1948 136 1956 144
rect 2060 136 2068 144
rect 2188 136 2196 144
rect 236 116 244 124
rect 412 116 420 124
rect 476 116 484 124
rect 556 116 564 124
rect 620 116 628 124
rect 700 116 708 124
rect 732 116 740 124
rect 764 116 772 124
rect 780 116 788 124
rect 796 116 804 124
rect 860 116 868 124
rect 940 116 948 124
rect 1004 116 1012 124
rect 1100 116 1108 124
rect 1116 116 1124 124
rect 1180 116 1188 124
rect 1324 116 1332 124
rect 1340 116 1348 124
rect 1356 116 1364 124
rect 1372 116 1380 124
rect 1436 116 1444 124
rect 1484 116 1492 124
rect 1708 116 1716 124
rect 1900 116 1908 124
rect 1932 116 1940 124
rect 1996 116 2004 124
rect 2156 116 2164 124
rect 2172 116 2180 124
rect 2188 116 2196 124
rect 60 96 68 104
rect 156 96 164 104
rect 188 96 196 104
rect 252 96 260 104
rect 332 96 340 104
rect 444 96 452 104
rect 524 96 532 104
rect 812 96 820 104
rect 1180 96 1188 104
rect 1324 96 1332 104
rect 1532 96 1540 104
rect 1772 96 1780 104
rect 1884 96 1892 104
rect 2012 96 2020 104
rect 2028 96 2036 104
rect 2060 96 2068 104
rect 2124 96 2132 104
rect 2140 96 2148 104
rect 12 76 20 84
rect 348 76 356 84
rect 1852 76 1860 84
rect 1980 76 1988 84
rect 2252 76 2260 84
rect 1996 56 2004 64
rect 972 36 980 44
rect 1420 36 1428 44
rect 1468 36 1476 44
rect 1516 36 1524 44
rect 622 6 630 14
rect 636 6 644 14
rect 650 6 658 14
<< metal2 >>
rect 45 1324 51 1496
rect 61 1464 67 1496
rect 77 1484 83 1536
rect 157 1524 163 1536
rect 157 1504 163 1516
rect 237 1504 243 1536
rect 125 1484 131 1496
rect 93 1344 99 1356
rect 13 1284 19 1296
rect 109 1283 115 1436
rect 141 1324 147 1436
rect 141 1304 147 1316
rect 157 1304 163 1336
rect 205 1324 211 1496
rect 221 1484 227 1496
rect 317 1484 323 1516
rect 269 1323 275 1436
rect 260 1317 275 1323
rect 109 1277 124 1283
rect 189 1244 195 1316
rect 317 1304 323 1356
rect 333 1324 339 1516
rect 349 1484 355 1643
rect 397 1524 403 1643
rect 573 1637 595 1643
rect 669 1637 691 1643
rect 589 1584 595 1637
rect 616 1606 622 1614
rect 630 1606 636 1614
rect 644 1606 650 1614
rect 658 1606 664 1614
rect 429 1524 435 1556
rect 349 1383 355 1476
rect 381 1444 387 1496
rect 349 1377 371 1383
rect 365 1364 371 1377
rect 365 1344 371 1356
rect 381 1304 387 1436
rect 445 1364 451 1516
rect 637 1484 643 1516
rect 685 1484 691 1637
rect 717 1484 723 1643
rect 973 1604 979 1643
rect 957 1544 963 1556
rect 1181 1524 1187 1536
rect 781 1484 787 1496
rect 877 1484 883 1496
rect 941 1483 947 1516
rect 989 1504 995 1516
rect 1005 1483 1011 1496
rect 1021 1484 1027 1496
rect 941 1477 1011 1483
rect 413 1324 419 1356
rect 429 1344 435 1356
rect 541 1344 547 1476
rect 397 1304 403 1316
rect 413 1304 419 1316
rect 509 1304 515 1336
rect 557 1304 563 1436
rect 589 1364 595 1436
rect 653 1364 659 1456
rect 653 1344 659 1356
rect 669 1324 675 1476
rect 109 1104 115 1136
rect 13 1084 19 1096
rect 77 1084 83 1096
rect 45 1044 51 1080
rect 77 1064 83 1076
rect 77 1004 83 1056
rect 109 1044 115 1096
rect 125 1084 131 1096
rect 141 1084 147 1096
rect 141 964 147 1056
rect 157 944 163 1236
rect 616 1206 622 1214
rect 630 1206 636 1214
rect 644 1206 650 1214
rect 658 1206 664 1214
rect 349 1144 355 1156
rect 685 1144 691 1436
rect 717 1364 723 1476
rect 765 1464 771 1476
rect 829 1464 835 1476
rect 877 1324 883 1476
rect 1069 1464 1075 1516
rect 925 1364 931 1456
rect 989 1384 995 1436
rect 1069 1384 1075 1456
rect 909 1324 915 1336
rect 781 1304 787 1316
rect 797 1297 812 1303
rect 221 1124 227 1136
rect 717 1124 723 1136
rect 685 1117 700 1123
rect 237 1064 243 1116
rect 317 1103 323 1116
rect 317 1097 348 1103
rect 205 964 211 996
rect 45 924 51 936
rect 61 924 67 936
rect 13 884 19 896
rect 13 664 19 716
rect 61 544 67 916
rect 77 904 83 916
rect 109 904 115 936
rect 157 924 163 936
rect 189 904 195 956
rect 205 944 211 956
rect 221 924 227 936
rect 157 724 163 756
rect 237 743 243 1056
rect 269 1044 275 1076
rect 269 924 275 1036
rect 285 984 291 996
rect 301 944 307 1096
rect 349 1004 355 1096
rect 525 1084 531 1116
rect 557 1084 563 1096
rect 413 944 419 956
rect 349 924 355 936
rect 269 904 275 916
rect 365 904 371 916
rect 445 904 451 956
rect 509 924 515 1036
rect 525 924 531 1076
rect 541 944 547 1036
rect 557 964 563 1076
rect 541 904 547 936
rect 573 924 579 936
rect 349 864 355 896
rect 445 764 451 896
rect 653 884 659 1076
rect 685 1023 691 1117
rect 749 1104 755 1236
rect 797 1064 803 1297
rect 861 1184 867 1296
rect 877 1144 883 1236
rect 829 1104 835 1136
rect 941 1123 947 1356
rect 1213 1344 1219 1643
rect 1245 1463 1251 1643
rect 1309 1637 1331 1643
rect 1325 1584 1331 1637
rect 1229 1457 1251 1463
rect 925 1117 947 1123
rect 877 1104 883 1116
rect 925 1084 931 1117
rect 973 1104 979 1316
rect 1037 1304 1043 1316
rect 1085 1304 1091 1336
rect 1101 1304 1107 1316
rect 989 1284 995 1296
rect 1117 1284 1123 1336
rect 1213 1324 1219 1336
rect 1149 1304 1155 1316
rect 685 1017 707 1023
rect 701 984 707 1017
rect 717 1004 723 1036
rect 749 904 755 956
rect 797 944 803 1056
rect 877 984 883 1036
rect 765 904 771 936
rect 781 924 787 936
rect 813 904 819 976
rect 845 924 851 976
rect 925 963 931 1076
rect 925 957 940 963
rect 957 944 963 1096
rect 989 1084 995 1276
rect 1101 1124 1107 1236
rect 1053 1044 1059 1116
rect 1133 1084 1139 1256
rect 1229 1184 1235 1457
rect 1277 1384 1283 1516
rect 1357 1504 1363 1516
rect 1293 1344 1299 1476
rect 1341 1424 1347 1476
rect 1373 1424 1379 1643
rect 1437 1524 1443 1643
rect 1517 1637 1539 1643
rect 1533 1584 1539 1637
rect 1549 1524 1555 1536
rect 1309 1364 1315 1376
rect 1293 1264 1299 1336
rect 1309 1304 1315 1356
rect 1188 1117 1203 1123
rect 989 944 995 956
rect 957 924 963 936
rect 1133 884 1139 1076
rect 1197 984 1203 1117
rect 1277 1104 1283 1116
rect 1341 1104 1347 1116
rect 1357 1084 1363 1416
rect 1389 1323 1395 1436
rect 1405 1424 1411 1476
rect 1405 1344 1411 1356
rect 1437 1343 1443 1436
rect 1469 1364 1475 1416
rect 1517 1344 1523 1516
rect 1677 1504 1683 1576
rect 1853 1563 1859 1643
rect 1853 1557 1875 1563
rect 1821 1544 1827 1556
rect 1709 1464 1715 1516
rect 1789 1504 1795 1516
rect 1757 1484 1763 1496
rect 1576 1406 1582 1414
rect 1590 1406 1596 1414
rect 1604 1406 1610 1414
rect 1618 1406 1624 1414
rect 1869 1384 1875 1557
rect 1901 1504 1907 1556
rect 1917 1484 1923 1643
rect 1965 1564 1971 1643
rect 1933 1524 1939 1556
rect 2013 1504 2019 1556
rect 2125 1484 2131 1516
rect 1917 1464 1923 1476
rect 1981 1464 1987 1476
rect 2093 1424 2099 1476
rect 1981 1384 1987 1416
rect 2100 1397 2115 1403
rect 1693 1344 1699 1376
rect 2093 1344 2099 1356
rect 1437 1337 1459 1343
rect 1380 1317 1395 1323
rect 1405 1304 1411 1336
rect 1453 1324 1459 1337
rect 1421 1284 1427 1316
rect 1389 1084 1395 1116
rect 1309 1064 1315 1076
rect 1405 1064 1411 1076
rect 1245 923 1251 1036
rect 1293 964 1299 996
rect 1245 917 1260 923
rect 1293 904 1299 956
rect 1325 944 1331 1036
rect 1373 944 1379 1036
rect 1325 924 1331 936
rect 1213 884 1219 896
rect 237 737 259 743
rect 77 684 83 716
rect 109 684 115 716
rect 77 664 83 676
rect 109 644 115 676
rect 173 624 179 716
rect 237 704 243 716
rect 253 704 259 737
rect 228 677 243 683
rect 13 484 19 496
rect 61 304 67 536
rect 77 524 83 556
rect 157 504 163 596
rect 189 564 195 636
rect 205 584 211 616
rect 237 584 243 677
rect 221 504 227 556
rect 269 543 275 696
rect 285 624 291 676
rect 301 644 307 696
rect 381 684 387 716
rect 333 664 339 676
rect 269 537 284 543
rect 333 540 339 636
rect 349 544 355 656
rect 381 644 387 676
rect 365 524 371 636
rect 397 564 403 656
rect 397 544 403 556
rect 429 540 435 636
rect 461 604 467 636
rect 477 544 483 556
rect 493 504 499 676
rect 525 504 531 656
rect 589 544 595 876
rect 616 806 622 814
rect 630 806 636 814
rect 644 806 650 814
rect 658 806 664 814
rect 685 704 691 756
rect 717 724 723 876
rect 701 704 707 716
rect 669 564 675 696
rect 765 664 771 756
rect 829 744 835 756
rect 957 744 963 776
rect 1165 744 1171 756
rect 605 504 611 516
rect 701 504 707 576
rect 717 504 723 636
rect 765 584 771 636
rect 733 524 739 556
rect 781 544 787 716
rect 813 644 819 736
rect 861 724 867 736
rect 1293 724 1299 736
rect 1357 724 1363 916
rect 1373 904 1379 936
rect 1405 924 1411 936
rect 1421 884 1427 956
rect 1437 863 1443 1316
rect 1453 1304 1459 1316
rect 1485 1184 1491 1256
rect 1517 1124 1523 1336
rect 1917 1324 1923 1336
rect 1805 1297 1820 1303
rect 1805 1264 1811 1297
rect 1821 1184 1827 1276
rect 1885 1244 1891 1276
rect 1620 1117 1635 1123
rect 1453 964 1459 1036
rect 1453 924 1459 936
rect 1469 884 1475 1076
rect 1501 983 1507 1116
rect 1629 1104 1635 1117
rect 1636 1097 1651 1103
rect 1492 977 1507 983
rect 1517 964 1523 1076
rect 1533 924 1539 1036
rect 1549 964 1555 1076
rect 1576 1006 1582 1014
rect 1590 1006 1596 1014
rect 1604 1006 1610 1014
rect 1618 1006 1624 1014
rect 1645 924 1651 1097
rect 1677 1064 1683 1156
rect 1709 1084 1715 1096
rect 1661 924 1667 1036
rect 1725 964 1731 1116
rect 1757 1104 1763 1116
rect 1789 1104 1795 1116
rect 1901 1104 1907 1116
rect 1933 1104 1939 1336
rect 1949 1324 1955 1336
rect 1981 1324 1987 1336
rect 1981 1284 1987 1296
rect 2061 1124 2067 1316
rect 2077 1124 2083 1316
rect 2093 1124 2099 1336
rect 2109 1304 2115 1397
rect 2125 1344 2131 1356
rect 2141 1344 2147 1436
rect 2221 1383 2227 1456
rect 2212 1377 2227 1383
rect 2173 1344 2179 1356
rect 2157 1324 2163 1336
rect 2205 1324 2211 1336
rect 2141 1163 2147 1316
rect 2157 1184 2163 1296
rect 2253 1284 2259 1296
rect 2141 1157 2163 1163
rect 2157 1123 2163 1157
rect 2157 1117 2179 1123
rect 2013 1104 2019 1116
rect 2061 1104 2067 1116
rect 1901 1084 1907 1096
rect 1933 1084 1939 1096
rect 2093 1084 2099 1116
rect 2004 1077 2019 1083
rect 1949 1064 1955 1076
rect 2013 1044 2019 1077
rect 2093 1064 2099 1076
rect 2109 1044 2115 1116
rect 2125 1084 2131 1096
rect 1869 964 1875 996
rect 1981 964 1987 996
rect 1997 964 2003 996
rect 2013 984 2019 1036
rect 2045 964 2051 1036
rect 1501 904 1507 916
rect 1645 904 1651 916
rect 1725 904 1731 956
rect 1869 944 1875 956
rect 1853 904 1859 936
rect 1901 904 1907 916
rect 1949 904 1955 916
rect 1476 877 1491 883
rect 1421 857 1443 863
rect 829 584 835 696
rect 909 564 915 676
rect 925 644 931 696
rect 1005 683 1011 716
rect 1197 704 1203 716
rect 1229 684 1235 696
rect 996 677 1011 683
rect 980 657 988 663
rect 973 584 979 636
rect 989 564 995 656
rect 813 544 819 556
rect 877 544 883 556
rect 1005 544 1011 677
rect 1261 677 1331 683
rect 1037 664 1043 676
rect 1117 664 1123 676
rect 829 524 835 536
rect 829 504 835 516
rect 109 324 115 356
rect 157 324 163 336
rect 61 284 67 296
rect 205 284 211 296
rect 61 144 67 276
rect 237 264 243 496
rect 317 284 323 296
rect 285 264 291 276
rect 77 103 83 236
rect 189 144 195 176
rect 285 144 291 256
rect 317 243 323 276
rect 333 264 339 336
rect 397 304 403 496
rect 461 344 467 356
rect 413 304 419 316
rect 317 237 339 243
rect 317 144 323 156
rect 333 144 339 237
rect 381 184 387 256
rect 445 184 451 296
rect 541 284 547 436
rect 557 384 563 496
rect 616 406 622 414
rect 630 406 636 414
rect 644 406 650 414
rect 658 406 664 414
rect 733 344 739 436
rect 909 424 915 516
rect 797 324 803 356
rect 68 97 83 103
rect 13 84 19 96
rect 237 84 243 116
rect 253 104 259 116
rect 333 104 339 136
rect 413 124 419 156
rect 429 124 435 136
rect 509 124 515 156
rect 541 144 547 256
rect 621 244 627 316
rect 717 224 723 296
rect 557 124 563 176
rect 573 144 579 156
rect 589 144 595 156
rect 717 143 723 176
rect 733 164 739 276
rect 749 144 755 276
rect 717 137 739 143
rect 525 104 531 116
rect 445 -23 451 96
rect 557 -23 563 16
rect 589 -23 595 136
rect 733 124 739 137
rect 765 124 771 156
rect 797 124 803 296
rect 877 284 883 416
rect 877 183 883 276
rect 861 177 883 183
rect 861 124 867 177
rect 893 164 899 256
rect 909 244 915 316
rect 909 184 915 216
rect 893 144 899 156
rect 925 144 931 536
rect 1005 524 1011 536
rect 1069 523 1075 636
rect 1213 564 1219 656
rect 1261 644 1267 677
rect 1277 644 1283 656
rect 1325 644 1331 677
rect 1197 544 1203 556
rect 1069 517 1084 523
rect 1085 504 1091 516
rect 1101 504 1107 536
rect 1277 524 1283 556
rect 1133 484 1139 516
rect 1149 504 1155 516
rect 1085 364 1091 436
rect 1133 384 1139 436
rect 1069 344 1075 356
rect 1005 324 1011 336
rect 941 244 947 296
rect 973 284 979 316
rect 1053 284 1059 296
rect 957 264 963 276
rect 621 104 627 116
rect 701 104 707 116
rect 861 104 867 116
rect 941 104 947 116
rect 616 6 622 14
rect 630 6 636 14
rect 644 6 650 14
rect 658 6 664 14
rect 781 -23 787 96
rect 957 -17 963 136
rect 1005 124 1011 236
rect 1021 224 1027 256
rect 1085 244 1091 336
rect 1165 304 1171 316
rect 1140 297 1155 303
rect 1149 264 1155 297
rect 1069 184 1075 236
rect 1149 184 1155 256
rect 1165 164 1171 296
rect 1181 264 1187 476
rect 1213 324 1219 356
rect 1277 324 1283 436
rect 1293 344 1299 636
rect 1325 564 1331 576
rect 1373 544 1379 656
rect 1389 584 1395 616
rect 1309 504 1315 536
rect 1405 524 1411 696
rect 1421 544 1427 857
rect 1485 724 1491 877
rect 1533 744 1539 836
rect 1501 724 1507 736
rect 1677 724 1683 836
rect 1805 724 1811 836
rect 1437 544 1443 656
rect 1453 644 1459 676
rect 1453 544 1459 576
rect 1357 324 1363 456
rect 1437 404 1443 536
rect 1245 284 1251 316
rect 1373 304 1379 316
rect 1437 304 1443 376
rect 1453 304 1459 536
rect 1469 464 1475 636
rect 1485 524 1491 716
rect 1501 564 1507 716
rect 1533 544 1539 716
rect 1725 704 1731 716
rect 1576 606 1582 614
rect 1590 606 1596 614
rect 1604 606 1610 614
rect 1618 606 1624 614
rect 1629 524 1635 536
rect 1645 524 1651 676
rect 1661 664 1667 676
rect 1677 544 1683 696
rect 1773 684 1779 716
rect 1997 704 2003 736
rect 2045 684 2051 836
rect 2061 704 2067 936
rect 2093 904 2099 956
rect 1757 664 1763 676
rect 1725 523 1731 636
rect 1757 524 1763 656
rect 1853 584 1859 676
rect 2061 564 2067 656
rect 2077 564 2083 716
rect 2093 684 2099 876
rect 2109 724 2115 916
rect 2141 724 2147 836
rect 2173 784 2179 1117
rect 2205 1084 2211 1096
rect 2205 924 2211 1076
rect 2221 1064 2227 1116
rect 2221 944 2227 956
rect 2109 604 2115 716
rect 2125 664 2131 676
rect 2157 664 2163 716
rect 2205 704 2211 916
rect 2221 904 2227 936
rect 1805 524 1811 556
rect 1853 524 1859 536
rect 1869 524 1875 536
rect 2029 524 2035 536
rect 2061 524 2067 556
rect 2157 524 2163 636
rect 1716 517 1731 523
rect 1949 517 1996 523
rect 1501 464 1507 496
rect 1469 324 1475 436
rect 1485 304 1491 316
rect 1421 284 1427 296
rect 1229 224 1235 256
rect 1277 184 1283 236
rect 1293 164 1299 216
rect 1133 144 1139 156
rect 1309 144 1315 276
rect 1101 104 1107 116
rect 941 -23 963 -17
rect 973 -17 979 36
rect 973 -23 995 -17
rect 1117 -23 1123 116
rect 1181 104 1187 116
rect 1245 104 1251 136
rect 1325 124 1331 156
rect 1357 124 1363 156
rect 1389 104 1395 236
rect 1437 124 1443 236
rect 1453 164 1459 296
rect 1517 284 1523 296
rect 1476 237 1491 243
rect 1485 124 1491 237
rect 1533 144 1539 516
rect 1661 484 1667 516
rect 1693 504 1699 516
rect 1709 504 1715 516
rect 1949 504 1955 517
rect 2029 504 2035 516
rect 1917 484 1923 496
rect 1613 324 1619 476
rect 1837 384 1843 436
rect 1773 324 1779 356
rect 1821 344 1827 356
rect 1613 264 1619 316
rect 2061 304 2067 516
rect 2141 464 2147 516
rect 2157 504 2163 516
rect 2173 504 2179 536
rect 2077 344 2083 456
rect 2157 384 2163 436
rect 2173 344 2179 476
rect 2189 464 2195 476
rect 2221 324 2227 896
rect 2237 684 2243 1056
rect 2253 964 2259 996
rect 2237 524 2243 656
rect 2237 504 2243 516
rect 1700 297 1715 303
rect 1645 264 1651 276
rect 1661 263 1667 296
rect 1661 257 1683 263
rect 1576 206 1582 214
rect 1590 206 1596 214
rect 1604 206 1610 214
rect 1618 206 1624 214
rect 1677 184 1683 257
rect 1581 144 1587 156
rect 1181 -23 1187 96
rect 1229 -23 1235 16
rect 1421 -17 1427 36
rect 1405 -23 1427 -17
rect 1437 -23 1443 36
rect 1469 -23 1475 36
rect 1517 -17 1523 36
rect 1501 -23 1523 -17
rect 1693 -23 1699 136
rect 1709 124 1715 297
rect 1741 264 1747 276
rect 1725 144 1731 256
rect 1773 184 1779 296
rect 1885 284 1891 296
rect 1789 144 1795 156
rect 1773 124 1779 136
rect 1885 124 1891 276
rect 1917 144 1923 256
rect 1933 244 1939 276
rect 1949 264 1955 276
rect 1933 124 1939 236
rect 2061 144 2067 276
rect 2093 164 2099 296
rect 2237 284 2243 496
rect 2109 184 2115 236
rect 2125 204 2131 276
rect 2253 264 2259 296
rect 1725 -23 1731 116
rect 1773 104 1779 116
rect 1885 104 1891 116
rect 2013 104 2019 136
rect 2141 104 2147 176
rect 2189 144 2195 196
rect 2173 104 2179 116
rect 2029 84 2035 96
rect 2253 84 2259 96
rect 1997 64 2003 76
<< m3contact >>
rect 76 1536 84 1544
rect 156 1536 164 1544
rect 236 1536 244 1544
rect 284 1536 292 1544
rect 60 1496 68 1504
rect 316 1516 324 1524
rect 332 1516 340 1524
rect 124 1496 132 1504
rect 220 1496 228 1504
rect 92 1356 100 1364
rect 12 1296 20 1304
rect 60 1296 68 1304
rect 92 1296 100 1304
rect 156 1336 164 1344
rect 220 1336 228 1344
rect 284 1356 292 1364
rect 300 1336 308 1344
rect 140 1296 148 1304
rect 172 1296 180 1304
rect 622 1606 630 1614
rect 636 1606 644 1614
rect 650 1606 658 1614
rect 412 1536 420 1544
rect 380 1516 388 1524
rect 396 1516 404 1524
rect 428 1516 436 1524
rect 508 1516 516 1524
rect 380 1496 388 1504
rect 428 1496 436 1504
rect 348 1356 356 1364
rect 364 1336 372 1344
rect 332 1316 340 1324
rect 972 1596 980 1604
rect 764 1536 772 1544
rect 940 1536 948 1544
rect 956 1536 964 1544
rect 1180 1536 1188 1544
rect 828 1516 836 1524
rect 940 1516 948 1524
rect 972 1516 980 1524
rect 1052 1516 1060 1524
rect 1068 1516 1076 1524
rect 1132 1516 1140 1524
rect 844 1496 852 1504
rect 604 1476 612 1484
rect 716 1476 724 1484
rect 764 1476 772 1484
rect 780 1476 788 1484
rect 876 1476 884 1484
rect 908 1476 916 1484
rect 956 1496 964 1504
rect 988 1496 996 1504
rect 1004 1496 1012 1504
rect 1020 1476 1028 1484
rect 412 1356 420 1364
rect 428 1356 436 1364
rect 444 1356 452 1364
rect 556 1436 564 1444
rect 588 1436 596 1444
rect 444 1336 452 1344
rect 460 1316 468 1324
rect 572 1356 580 1364
rect 652 1356 660 1364
rect 668 1316 676 1324
rect 284 1296 292 1304
rect 316 1296 324 1304
rect 396 1296 404 1304
rect 412 1296 420 1304
rect 508 1296 516 1304
rect 156 1236 164 1244
rect 188 1236 196 1244
rect 108 1136 116 1144
rect 76 1096 84 1104
rect 124 1096 132 1104
rect 12 1076 20 1084
rect 44 1036 52 1044
rect 140 1076 148 1084
rect 140 1056 148 1064
rect 108 1036 116 1044
rect 76 996 84 1004
rect 622 1206 630 1214
rect 636 1206 644 1214
rect 650 1206 658 1214
rect 764 1456 772 1464
rect 828 1456 836 1464
rect 716 1356 724 1364
rect 1100 1496 1108 1504
rect 1084 1476 1092 1484
rect 908 1456 916 1464
rect 924 1456 932 1464
rect 988 1376 996 1384
rect 940 1356 948 1364
rect 1196 1356 1204 1364
rect 748 1316 756 1324
rect 876 1316 884 1324
rect 908 1316 916 1324
rect 700 1296 708 1304
rect 780 1296 788 1304
rect 220 1136 228 1144
rect 348 1136 356 1144
rect 364 1136 372 1144
rect 396 1136 404 1144
rect 684 1136 692 1144
rect 716 1136 724 1144
rect 172 1116 180 1124
rect 236 1116 244 1124
rect 252 1116 260 1124
rect 332 1116 340 1124
rect 284 1096 292 1104
rect 300 1096 308 1104
rect 460 1096 468 1104
rect 268 1076 276 1084
rect 204 1056 212 1064
rect 204 996 212 1004
rect 188 956 196 964
rect 44 936 52 944
rect 92 936 100 944
rect 108 936 116 944
rect 172 936 180 944
rect 60 916 68 924
rect 12 896 20 904
rect 12 716 20 724
rect 28 676 36 684
rect 156 916 164 924
rect 204 936 212 944
rect 220 916 228 924
rect 76 896 84 904
rect 124 896 132 904
rect 76 736 84 744
rect 140 736 148 744
rect 268 1036 276 1044
rect 284 996 292 1004
rect 316 1056 324 1064
rect 556 1096 564 1104
rect 428 1076 436 1084
rect 476 1080 484 1084
rect 476 1076 484 1080
rect 524 1076 532 1084
rect 348 996 356 1004
rect 396 956 404 964
rect 412 956 420 964
rect 460 956 468 964
rect 300 936 308 944
rect 348 936 356 944
rect 268 916 276 924
rect 364 916 372 924
rect 412 916 420 924
rect 572 1056 580 1064
rect 540 936 548 944
rect 572 916 580 924
rect 348 896 356 904
rect 380 896 388 904
rect 540 896 548 904
rect 620 896 628 904
rect 252 876 260 884
rect 332 876 340 884
rect 844 1276 852 1284
rect 828 1136 836 1144
rect 844 1136 852 1144
rect 876 1136 884 1144
rect 1228 1476 1236 1484
rect 1356 1516 1364 1524
rect 1020 1336 1028 1344
rect 1084 1336 1092 1344
rect 1116 1336 1124 1344
rect 972 1316 980 1324
rect 876 1096 884 1104
rect 988 1296 996 1304
rect 1036 1296 1044 1304
rect 1068 1296 1076 1304
rect 1100 1296 1108 1304
rect 1148 1316 1156 1324
rect 1212 1316 1220 1324
rect 1164 1296 1172 1304
rect 940 1096 948 1104
rect 956 1096 964 1104
rect 972 1096 980 1104
rect 700 1036 708 1044
rect 716 996 724 1004
rect 812 976 820 984
rect 844 976 852 984
rect 876 976 884 984
rect 780 936 788 944
rect 940 956 948 964
rect 1132 1256 1140 1264
rect 1292 1476 1300 1484
rect 1676 1576 1684 1584
rect 1548 1536 1556 1544
rect 1436 1516 1444 1524
rect 1516 1516 1524 1524
rect 1644 1516 1652 1524
rect 1500 1496 1508 1504
rect 1340 1416 1348 1424
rect 1356 1416 1364 1424
rect 1372 1416 1380 1424
rect 1308 1376 1316 1384
rect 1340 1376 1348 1384
rect 1324 1356 1332 1364
rect 1244 1336 1252 1344
rect 1292 1336 1300 1344
rect 1260 1276 1268 1284
rect 1308 1296 1316 1304
rect 1340 1296 1348 1304
rect 1292 1256 1300 1264
rect 988 956 996 964
rect 972 936 980 944
rect 1068 936 1076 944
rect 956 916 964 924
rect 1020 916 1028 924
rect 764 896 772 904
rect 828 896 836 904
rect 876 896 884 904
rect 1276 1116 1284 1124
rect 1340 1116 1348 1124
rect 1404 1416 1412 1424
rect 1404 1356 1412 1364
rect 1468 1416 1476 1424
rect 1468 1356 1476 1364
rect 1500 1356 1508 1364
rect 1868 1576 1876 1584
rect 1820 1536 1828 1544
rect 1836 1536 1844 1544
rect 1708 1516 1716 1524
rect 1724 1516 1732 1524
rect 1804 1516 1812 1524
rect 1564 1496 1572 1504
rect 1692 1476 1700 1484
rect 1788 1496 1796 1504
rect 1820 1496 1828 1504
rect 1756 1476 1764 1484
rect 1788 1436 1796 1444
rect 1582 1406 1590 1414
rect 1596 1406 1604 1414
rect 1610 1406 1618 1414
rect 1900 1556 1908 1564
rect 1932 1556 1940 1564
rect 1964 1556 1972 1564
rect 2012 1556 2020 1564
rect 2076 1536 2084 1544
rect 1932 1496 1940 1504
rect 1996 1476 2004 1484
rect 2124 1476 2132 1484
rect 2188 1476 2196 1484
rect 1916 1456 1924 1464
rect 1980 1456 1988 1464
rect 2012 1456 2020 1464
rect 1980 1416 1988 1424
rect 2092 1416 2100 1424
rect 1692 1376 1700 1384
rect 1772 1336 1780 1344
rect 1916 1336 1924 1344
rect 1980 1336 1988 1344
rect 2044 1336 2052 1344
rect 2092 1336 2100 1344
rect 1452 1316 1460 1324
rect 1404 1296 1412 1304
rect 1420 1276 1428 1284
rect 1388 1116 1396 1124
rect 1308 1076 1316 1084
rect 1356 1076 1364 1084
rect 1404 1076 1412 1084
rect 1228 916 1236 924
rect 1292 996 1300 1004
rect 1276 936 1284 944
rect 1420 956 1428 964
rect 1324 936 1332 944
rect 1372 936 1380 944
rect 1404 936 1412 944
rect 1164 896 1172 904
rect 1228 896 1236 904
rect 1292 896 1300 904
rect 1308 896 1316 904
rect 588 876 596 884
rect 652 876 660 884
rect 716 876 724 884
rect 860 876 868 884
rect 892 876 900 884
rect 1132 876 1140 884
rect 1212 876 1220 884
rect 444 756 452 764
rect 76 716 84 724
rect 156 716 164 724
rect 188 716 196 724
rect 92 696 100 704
rect 156 696 164 704
rect 108 676 116 684
rect 76 656 84 664
rect 108 636 116 644
rect 444 736 452 744
rect 524 736 532 744
rect 460 716 468 724
rect 492 716 500 724
rect 236 696 244 704
rect 268 696 276 704
rect 316 696 324 704
rect 364 696 372 704
rect 172 616 180 624
rect 156 596 164 604
rect 76 556 84 564
rect 60 536 68 544
rect 44 516 52 524
rect 12 496 20 504
rect 124 536 132 544
rect 92 516 100 524
rect 204 616 212 624
rect 172 556 180 564
rect 540 696 548 704
rect 332 656 340 664
rect 348 656 356 664
rect 300 636 308 644
rect 332 636 340 644
rect 284 616 292 624
rect 396 656 404 664
rect 364 636 372 644
rect 380 636 388 644
rect 428 636 436 644
rect 380 556 388 564
rect 460 596 468 604
rect 476 556 484 564
rect 524 656 532 664
rect 572 656 580 664
rect 622 806 630 814
rect 636 806 644 814
rect 650 806 658 814
rect 684 756 692 764
rect 700 696 708 704
rect 748 676 756 684
rect 828 736 836 744
rect 860 736 868 744
rect 1036 736 1044 744
rect 1148 736 1156 744
rect 1164 736 1172 744
rect 1292 736 1300 744
rect 780 716 788 724
rect 764 636 772 644
rect 700 576 708 584
rect 668 556 676 564
rect 588 536 596 544
rect 588 516 596 524
rect 620 516 628 524
rect 732 556 740 564
rect 1388 896 1396 904
rect 1484 1276 1492 1284
rect 1484 1256 1492 1264
rect 1644 1316 1652 1324
rect 1900 1316 1908 1324
rect 1628 1296 1636 1304
rect 1692 1296 1700 1304
rect 1724 1296 1732 1304
rect 1820 1276 1828 1284
rect 1804 1256 1812 1264
rect 1516 1116 1524 1124
rect 1452 956 1460 964
rect 1452 916 1460 924
rect 1452 896 1460 904
rect 1516 956 1524 964
rect 1582 1006 1590 1014
rect 1596 1006 1604 1014
rect 1610 1006 1618 1014
rect 1548 956 1556 964
rect 1612 956 1620 964
rect 1548 936 1556 944
rect 1804 1136 1812 1144
rect 1836 1136 1844 1144
rect 1692 1116 1700 1124
rect 1772 1116 1780 1124
rect 1788 1116 1796 1124
rect 1916 1116 1924 1124
rect 1708 1076 1716 1084
rect 1948 1316 1956 1324
rect 2028 1316 2036 1324
rect 2060 1316 2068 1324
rect 2076 1316 2084 1324
rect 1980 1276 1988 1284
rect 2124 1356 2132 1364
rect 2172 1356 2180 1364
rect 2140 1336 2148 1344
rect 2204 1336 2212 1344
rect 2156 1316 2164 1324
rect 2156 1296 2164 1304
rect 2204 1296 2212 1304
rect 2252 1296 2260 1304
rect 2140 1136 2148 1144
rect 2012 1116 2020 1124
rect 2076 1116 2084 1124
rect 2092 1116 2100 1124
rect 2172 1136 2180 1144
rect 1756 1096 1764 1104
rect 1788 1096 1796 1104
rect 1900 1096 1908 1104
rect 1980 1096 1988 1104
rect 2060 1096 2068 1104
rect 1932 1076 1940 1084
rect 1884 1056 1892 1064
rect 1948 1056 1956 1064
rect 2076 1076 2084 1084
rect 2092 1056 2100 1064
rect 2124 1076 2132 1084
rect 2012 1036 2020 1044
rect 2108 1036 2116 1044
rect 1868 996 1876 1004
rect 1980 996 1988 1004
rect 1868 956 1876 964
rect 2044 956 2052 964
rect 2092 956 2100 964
rect 1500 916 1508 924
rect 1532 916 1540 924
rect 1740 936 1748 944
rect 1996 936 2004 944
rect 2028 936 2036 944
rect 2060 936 2068 944
rect 1772 916 1780 924
rect 1932 916 1940 924
rect 2044 916 2052 924
rect 1484 896 1492 904
rect 1644 896 1652 904
rect 1852 896 1860 904
rect 1900 896 1908 904
rect 1948 896 1956 904
rect 1468 876 1476 884
rect 844 716 852 724
rect 1004 716 1012 724
rect 1068 716 1076 724
rect 1180 716 1188 724
rect 1260 716 1268 724
rect 1340 716 1348 724
rect 1356 716 1364 724
rect 812 636 820 644
rect 876 676 884 684
rect 892 676 900 684
rect 828 576 836 584
rect 940 676 948 684
rect 1116 696 1124 704
rect 1164 696 1172 704
rect 1196 696 1204 704
rect 1372 696 1380 704
rect 988 656 996 664
rect 924 636 932 644
rect 972 636 980 644
rect 908 556 916 564
rect 1228 676 1236 684
rect 1036 656 1044 664
rect 1116 656 1124 664
rect 1212 656 1220 664
rect 1196 636 1204 644
rect 748 536 756 544
rect 780 536 788 544
rect 812 536 820 544
rect 876 536 884 544
rect 924 536 932 544
rect 828 516 836 524
rect 908 516 916 524
rect 396 496 404 504
rect 524 496 532 504
rect 556 496 564 504
rect 604 496 612 504
rect 636 496 644 504
rect 716 496 724 504
rect 108 356 116 364
rect 156 336 164 344
rect 204 296 212 304
rect 332 336 340 344
rect 300 296 308 304
rect 252 280 260 284
rect 252 276 260 280
rect 316 276 324 284
rect 236 256 244 264
rect 60 136 68 144
rect 12 96 20 104
rect 188 176 196 184
rect 348 316 356 324
rect 444 356 452 364
rect 460 356 468 364
rect 492 356 500 364
rect 428 316 436 324
rect 380 296 388 304
rect 412 296 420 304
rect 444 296 452 304
rect 380 256 388 264
rect 622 406 630 414
rect 636 406 644 414
rect 650 406 658 414
rect 876 416 884 424
rect 908 416 916 424
rect 732 336 740 344
rect 812 336 820 344
rect 844 336 852 344
rect 588 316 596 324
rect 796 316 804 324
rect 524 276 532 284
rect 540 276 548 284
rect 524 176 532 184
rect 412 156 420 164
rect 108 136 116 144
rect 284 136 292 144
rect 316 136 324 144
rect 364 136 372 144
rect 252 116 260 124
rect 156 96 164 104
rect 188 96 196 104
rect 476 136 484 144
rect 716 216 724 224
rect 556 176 564 184
rect 716 176 724 184
rect 540 136 548 144
rect 572 156 580 164
rect 588 136 596 144
rect 684 136 692 144
rect 732 156 740 164
rect 764 156 772 164
rect 428 116 436 124
rect 476 116 484 124
rect 508 116 516 124
rect 524 116 532 124
rect 332 96 340 104
rect 444 96 452 104
rect 236 76 244 84
rect 348 76 356 84
rect 556 16 564 24
rect 860 236 868 244
rect 844 136 852 144
rect 908 236 916 244
rect 908 216 916 224
rect 876 156 884 164
rect 940 516 948 524
rect 1004 516 1012 524
rect 1388 676 1396 684
rect 1372 656 1380 664
rect 1260 636 1268 644
rect 1276 636 1284 644
rect 1324 636 1332 644
rect 1276 556 1284 564
rect 1100 536 1108 544
rect 1164 536 1172 544
rect 1196 536 1204 544
rect 1244 516 1252 524
rect 1084 496 1092 504
rect 1116 496 1124 504
rect 1148 496 1156 504
rect 1228 496 1236 504
rect 1036 476 1044 484
rect 1068 476 1076 484
rect 1132 476 1140 484
rect 1180 476 1188 484
rect 1132 436 1140 444
rect 1084 356 1092 364
rect 1004 336 1012 344
rect 1068 336 1076 344
rect 940 316 948 324
rect 972 316 980 324
rect 1068 296 1076 304
rect 1052 276 1060 284
rect 956 256 964 264
rect 940 236 948 244
rect 892 136 900 144
rect 924 136 932 144
rect 956 136 964 144
rect 780 116 788 124
rect 620 96 628 104
rect 700 96 708 104
rect 780 96 788 104
rect 812 96 820 104
rect 860 96 868 104
rect 940 96 948 104
rect 622 6 630 14
rect 636 6 644 14
rect 650 6 658 14
rect 1116 276 1124 284
rect 1164 296 1172 304
rect 1148 256 1156 264
rect 1068 236 1076 244
rect 1084 236 1092 244
rect 1212 356 1220 364
rect 1324 556 1332 564
rect 1388 616 1396 624
rect 1308 536 1316 544
rect 1788 876 1796 884
rect 1820 876 1828 884
rect 1500 736 1508 744
rect 1532 736 1540 744
rect 1676 716 1684 724
rect 1772 716 1780 724
rect 1436 656 1444 664
rect 1452 636 1460 644
rect 1452 576 1460 584
rect 1420 536 1428 544
rect 1356 516 1364 524
rect 1404 516 1412 524
rect 1420 516 1428 524
rect 1356 456 1364 464
rect 1436 396 1444 404
rect 1436 376 1444 384
rect 1244 316 1252 324
rect 1276 316 1284 324
rect 1212 296 1220 304
rect 1500 556 1508 564
rect 1644 696 1652 704
rect 1676 696 1684 704
rect 1724 696 1732 704
rect 1548 676 1556 684
rect 1644 676 1652 684
rect 1582 606 1590 614
rect 1596 606 1604 614
rect 1610 606 1618 614
rect 1548 556 1556 564
rect 1660 656 1668 664
rect 2012 716 2020 724
rect 1884 696 1892 704
rect 1948 696 1956 704
rect 1996 696 2004 704
rect 2108 916 2116 924
rect 2140 916 2148 924
rect 1692 676 1700 684
rect 1852 676 1860 684
rect 1916 676 1924 684
rect 2060 676 2068 684
rect 1708 656 1716 664
rect 1756 656 1764 664
rect 1676 536 1684 544
rect 1484 516 1492 524
rect 1532 516 1540 524
rect 1628 516 1636 524
rect 1692 516 1700 524
rect 1948 656 1956 664
rect 2028 656 2036 664
rect 2060 656 2068 664
rect 1852 576 1860 584
rect 2156 876 2164 884
rect 2220 1116 2228 1124
rect 2204 1096 2212 1104
rect 2220 956 2228 964
rect 2204 916 2212 924
rect 2188 876 2196 884
rect 2140 716 2148 724
rect 2092 676 2100 684
rect 2220 896 2228 904
rect 2124 656 2132 664
rect 2156 656 2164 664
rect 2108 596 2116 604
rect 1820 556 1828 564
rect 1932 556 1940 564
rect 2076 556 2084 564
rect 1788 536 1796 544
rect 1868 536 1876 544
rect 2028 536 2036 544
rect 2108 536 2116 544
rect 2172 536 2180 544
rect 1756 516 1764 524
rect 1804 516 1812 524
rect 1852 516 1860 524
rect 1468 456 1476 464
rect 1500 456 1508 464
rect 1324 296 1332 304
rect 1372 296 1380 304
rect 1420 296 1428 304
rect 1452 296 1460 304
rect 1484 296 1492 304
rect 1260 276 1268 284
rect 1308 276 1316 284
rect 1404 276 1412 284
rect 1276 236 1284 244
rect 1292 236 1300 244
rect 1228 216 1236 224
rect 1292 216 1300 224
rect 1356 236 1364 244
rect 1436 236 1444 244
rect 1324 156 1332 164
rect 1356 156 1364 164
rect 1132 136 1140 144
rect 1212 136 1220 144
rect 1308 136 1316 144
rect 1100 96 1108 104
rect 1372 136 1380 144
rect 1340 116 1348 124
rect 1372 116 1380 124
rect 1484 276 1492 284
rect 1516 276 1524 284
rect 1452 156 1460 164
rect 2060 516 2068 524
rect 2076 516 2084 524
rect 2124 516 2132 524
rect 2156 516 2164 524
rect 1676 496 1684 504
rect 1708 496 1716 504
rect 1900 496 1908 504
rect 1948 496 1956 504
rect 1964 496 1972 504
rect 2028 496 2036 504
rect 1612 476 1620 484
rect 1660 476 1668 484
rect 1724 476 1732 484
rect 1756 476 1764 484
rect 1916 476 1924 484
rect 1708 456 1716 464
rect 1836 376 1844 384
rect 1772 356 1780 364
rect 1804 356 1812 364
rect 1820 356 1828 364
rect 1852 356 1860 364
rect 1756 336 1764 344
rect 1596 316 1604 324
rect 1788 316 1796 324
rect 2188 516 2196 524
rect 2188 476 2196 484
rect 2076 456 2084 464
rect 2140 456 2148 464
rect 2156 436 2164 444
rect 2092 336 2100 344
rect 2252 996 2260 1004
rect 2236 656 2244 664
rect 2236 516 2244 524
rect 2236 496 2244 504
rect 2140 316 2148 324
rect 2220 316 2228 324
rect 1644 256 1652 264
rect 1676 276 1684 284
rect 1582 206 1590 214
rect 1596 206 1604 214
rect 1610 206 1618 214
rect 1580 156 1588 164
rect 1660 156 1668 164
rect 1532 136 1540 144
rect 1692 136 1700 144
rect 1180 96 1188 104
rect 1244 96 1252 104
rect 1324 96 1332 104
rect 1388 96 1396 104
rect 1532 96 1540 104
rect 1436 36 1444 44
rect 1228 16 1236 24
rect 1772 296 1780 304
rect 1804 296 1812 304
rect 1884 296 1892 304
rect 1980 296 1988 304
rect 2060 296 2068 304
rect 1740 256 1748 264
rect 1932 276 1940 284
rect 2028 276 2036 284
rect 1740 136 1748 144
rect 1788 136 1796 144
rect 1852 136 1860 144
rect 1916 256 1924 264
rect 1900 156 1908 164
rect 1948 256 1956 264
rect 1916 136 1924 144
rect 2044 156 2052 164
rect 2252 296 2260 304
rect 2124 276 2132 284
rect 2172 276 2180 284
rect 2124 196 2132 204
rect 2188 196 2196 204
rect 2108 176 2116 184
rect 2140 176 2148 184
rect 2108 156 2116 164
rect 1948 136 1956 144
rect 2012 136 2020 144
rect 1708 116 1716 124
rect 1724 116 1732 124
rect 1772 116 1780 124
rect 1884 116 1892 124
rect 1900 116 1908 124
rect 1996 116 2004 124
rect 2156 116 2164 124
rect 2188 116 2196 124
rect 2012 96 2020 104
rect 2060 96 2068 104
rect 2124 96 2132 104
rect 2172 96 2180 104
rect 2252 96 2260 104
rect 1852 76 1860 84
rect 1980 76 1988 84
rect 1996 76 2004 84
rect 2028 76 2036 84
<< metal3 >>
rect 616 1614 664 1616
rect 616 1606 620 1614
rect 630 1606 636 1614
rect 644 1606 650 1614
rect 660 1606 664 1614
rect 616 1604 664 1606
rect 1684 1577 1868 1583
rect 1908 1557 1932 1563
rect 1940 1557 1964 1563
rect 1972 1557 2012 1563
rect -19 1537 76 1543
rect 84 1537 156 1543
rect 164 1537 236 1543
rect 292 1537 412 1543
rect 772 1537 940 1543
rect 964 1537 1180 1543
rect 1556 1537 1820 1543
rect 1844 1537 2076 1543
rect 324 1517 332 1523
rect 340 1517 380 1523
rect 388 1517 396 1523
rect 436 1517 508 1523
rect 836 1517 940 1523
rect 980 1517 1052 1523
rect 1076 1517 1132 1523
rect 1364 1517 1436 1523
rect 1444 1517 1516 1523
rect 1652 1517 1708 1523
rect 1732 1517 1804 1523
rect -19 1497 60 1503
rect 68 1497 124 1503
rect 132 1497 220 1503
rect 388 1497 428 1503
rect 852 1497 956 1503
rect 964 1497 988 1503
rect 1012 1497 1100 1503
rect 1508 1497 1564 1503
rect 1796 1497 1820 1503
rect 1828 1497 1932 1503
rect 612 1477 716 1483
rect 724 1477 764 1483
rect 788 1477 876 1483
rect 916 1477 1020 1483
rect 1028 1477 1084 1483
rect 1236 1477 1292 1483
rect 1700 1477 1756 1483
rect 1764 1477 1996 1483
rect 2100 1477 2124 1483
rect 2132 1477 2188 1483
rect 772 1457 828 1463
rect 836 1457 908 1463
rect 916 1457 924 1463
rect 1924 1457 1980 1463
rect 1988 1457 2012 1463
rect 564 1437 588 1443
rect 596 1437 1788 1443
rect 1348 1417 1356 1423
rect 1364 1417 1372 1423
rect 1380 1417 1404 1423
rect 1412 1417 1468 1423
rect 1988 1417 2092 1423
rect 1576 1414 1624 1416
rect 1576 1406 1580 1414
rect 1590 1406 1596 1414
rect 1604 1406 1610 1414
rect 1620 1406 1624 1414
rect 1576 1404 1624 1406
rect 996 1377 1308 1383
rect 1348 1377 1692 1383
rect 100 1357 284 1363
rect 356 1357 412 1363
rect 436 1357 444 1363
rect 452 1357 572 1363
rect 660 1357 716 1363
rect 948 1357 972 1363
rect 980 1357 1196 1363
rect 1332 1357 1404 1363
rect 1476 1357 1500 1363
rect 2132 1357 2172 1363
rect 164 1337 220 1343
rect 228 1337 300 1343
rect 372 1337 444 1343
rect 1028 1337 1084 1343
rect 1124 1337 1244 1343
rect 1300 1337 1772 1343
rect 1924 1337 1980 1343
rect 2052 1337 2092 1343
rect 2148 1337 2204 1343
rect 340 1317 460 1323
rect 676 1317 748 1323
rect 756 1317 876 1323
rect 884 1317 908 1323
rect 980 1317 1148 1323
rect 1156 1317 1212 1323
rect 1460 1317 1644 1323
rect 1908 1317 1948 1323
rect 2036 1317 2060 1323
rect 2084 1317 2156 1323
rect -19 1297 12 1303
rect 68 1297 92 1303
rect 148 1297 172 1303
rect 292 1297 316 1303
rect 324 1297 396 1303
rect 420 1297 508 1303
rect 708 1297 780 1303
rect 996 1297 1036 1303
rect 1076 1297 1100 1303
rect 1108 1297 1164 1303
rect 1316 1297 1340 1303
rect 1412 1297 1628 1303
rect 1700 1297 1724 1303
rect 2164 1297 2204 1303
rect 2260 1297 2291 1303
rect 852 1277 1260 1283
rect 1428 1277 1484 1283
rect 1828 1277 1980 1283
rect 1140 1257 1292 1263
rect 1492 1257 1804 1263
rect 164 1237 188 1243
rect 616 1214 664 1216
rect 616 1206 620 1214
rect 630 1206 636 1214
rect 644 1206 650 1214
rect 660 1206 664 1214
rect 616 1204 664 1206
rect -19 1137 108 1143
rect 228 1137 348 1143
rect 372 1137 396 1143
rect 692 1137 716 1143
rect 724 1137 828 1143
rect 852 1137 876 1143
rect 1812 1137 1836 1143
rect 2148 1137 2172 1143
rect 180 1117 236 1123
rect 260 1117 332 1123
rect 1284 1117 1340 1123
rect 1348 1117 1388 1123
rect 1396 1117 1516 1123
rect 1700 1117 1772 1123
rect 1796 1117 1916 1123
rect 2020 1117 2076 1123
rect 2100 1117 2220 1123
rect 2228 1117 2291 1123
rect -19 1097 76 1103
rect 132 1097 284 1103
rect 308 1097 460 1103
rect 468 1097 556 1103
rect 884 1097 940 1103
rect 948 1097 956 1103
rect 964 1097 972 1103
rect 1764 1097 1788 1103
rect 1908 1097 1980 1103
rect 1988 1097 2060 1103
rect 2068 1097 2204 1103
rect 20 1077 140 1083
rect 276 1077 428 1083
rect 436 1077 476 1083
rect 484 1077 524 1083
rect 1316 1077 1356 1083
rect 1364 1077 1404 1083
rect 1716 1077 1932 1083
rect 2084 1077 2124 1083
rect 148 1057 204 1063
rect 324 1057 572 1063
rect 1892 1057 1948 1063
rect 1956 1057 2092 1063
rect 52 1037 108 1043
rect 116 1037 268 1043
rect 708 1037 1292 1043
rect 2020 1037 2108 1043
rect 1576 1014 1624 1016
rect 1576 1006 1580 1014
rect 1590 1006 1596 1014
rect 1604 1006 1610 1014
rect 1620 1006 1624 1014
rect 1576 1004 1624 1006
rect 84 997 204 1003
rect 292 997 348 1003
rect 724 997 1292 1003
rect 1876 997 1980 1003
rect 1988 997 2172 1003
rect 2180 997 2252 1003
rect 2260 997 2291 1003
rect 820 977 844 983
rect 852 977 876 983
rect 196 957 396 963
rect 420 957 460 963
rect 948 957 988 963
rect 1428 957 1452 963
rect 1524 957 1548 963
rect 1556 957 1612 963
rect 1620 957 1868 963
rect 2052 957 2092 963
rect 2228 957 2291 963
rect 52 937 92 943
rect 116 937 172 943
rect 212 937 300 943
rect 356 937 540 943
rect 788 937 972 943
rect 980 937 1068 943
rect 1284 937 1324 943
rect 1380 937 1404 943
rect 1556 937 1740 943
rect 2004 937 2028 943
rect 2036 937 2060 943
rect 68 917 156 923
rect 228 917 268 923
rect 372 917 412 923
rect 420 917 572 923
rect 964 917 1020 923
rect 1236 917 1452 923
rect 1508 917 1532 923
rect 1540 917 1772 923
rect 1940 917 2044 923
rect 2116 917 2140 923
rect 2212 917 2291 923
rect -19 897 12 903
rect 84 897 124 903
rect 356 897 380 903
rect 548 897 620 903
rect 772 897 828 903
rect 884 897 1164 903
rect 1236 897 1292 903
rect 1316 897 1388 903
rect 1460 897 1484 903
rect 1652 897 1852 903
rect 1860 897 1900 903
rect 1908 897 1948 903
rect 1956 897 2220 903
rect 260 877 332 883
rect 596 877 652 883
rect 660 877 716 883
rect 868 877 892 883
rect 1140 877 1212 883
rect 1220 877 1468 883
rect 1796 877 1820 883
rect 2164 877 2188 883
rect 616 814 664 816
rect 616 806 620 814
rect 630 806 636 814
rect 644 806 650 814
rect 660 806 664 814
rect 616 804 664 806
rect 452 757 684 763
rect 84 737 140 743
rect 452 737 524 743
rect 836 737 860 743
rect 1044 737 1148 743
rect 1172 737 1292 743
rect 1508 737 1532 743
rect -19 717 12 723
rect 20 717 76 723
rect 164 717 188 723
rect 468 717 492 723
rect 788 717 844 723
rect 1012 717 1068 723
rect 1188 717 1260 723
rect 1316 717 1340 723
rect 1348 717 1356 723
rect 1684 717 1772 723
rect 2020 717 2140 723
rect 100 697 156 703
rect 164 697 236 703
rect 276 697 316 703
rect 372 697 540 703
rect 548 697 700 703
rect 1124 697 1164 703
rect 1172 697 1196 703
rect 1652 697 1676 703
rect 1684 697 1724 703
rect 1892 697 1948 703
rect 2004 697 2291 703
rect -19 677 28 683
rect 36 677 108 683
rect 756 677 876 683
rect 900 677 940 683
rect 1236 677 1388 683
rect 1556 677 1644 683
rect 1652 677 1692 683
rect 1860 677 1916 683
rect 2068 677 2092 683
rect 84 657 332 663
rect 340 657 348 663
rect 356 657 396 663
rect 532 657 572 663
rect 996 657 1036 663
rect 1044 657 1116 663
rect 1124 657 1212 663
rect 1220 657 1372 663
rect 1380 657 1436 663
rect 1668 657 1708 663
rect 1716 657 1756 663
rect 1956 657 2028 663
rect 2068 657 2124 663
rect 2164 657 2236 663
rect 116 637 300 643
rect 308 637 332 643
rect 340 637 364 643
rect 372 637 380 643
rect 388 637 428 643
rect 772 637 812 643
rect 932 637 972 643
rect 1204 637 1260 643
rect 1284 637 1308 643
rect 1332 637 1452 643
rect 180 617 204 623
rect 212 617 284 623
rect 1380 617 1388 623
rect 1576 614 1624 616
rect 1576 606 1580 614
rect 1590 606 1596 614
rect 1604 606 1610 614
rect 1620 606 1624 614
rect 1576 604 1624 606
rect 164 597 460 603
rect 708 577 828 583
rect 1300 577 1452 583
rect 1460 577 1852 583
rect 1860 577 2092 583
rect 84 557 172 563
rect 388 557 476 563
rect 484 557 668 563
rect 740 557 908 563
rect 1284 557 1324 563
rect 1508 557 1548 563
rect 1828 557 1932 563
rect 1972 557 2076 563
rect 68 537 124 543
rect 132 537 588 543
rect 756 537 780 543
rect 820 537 876 543
rect 884 537 924 543
rect 1108 537 1164 543
rect 1204 537 1308 543
rect 1316 537 1420 543
rect 1684 537 1788 543
rect 1796 537 1868 543
rect 1876 537 2028 543
rect 2116 537 2172 543
rect 52 517 92 523
rect 596 517 620 523
rect 836 517 908 523
rect 916 517 940 523
rect 1012 517 1228 523
rect 1236 517 1244 523
rect 1252 517 1356 523
rect 1364 517 1404 523
rect 1412 517 1420 523
rect 1492 517 1532 523
rect 1636 517 1692 523
rect 1764 517 1804 523
rect 1812 517 1852 523
rect 1860 517 2060 523
rect 2084 517 2124 523
rect 2164 517 2188 523
rect 2244 517 2291 523
rect -19 497 12 503
rect 404 497 524 503
rect 564 497 604 503
rect 644 497 716 503
rect 1092 497 1116 503
rect 1156 497 1228 503
rect 1684 497 1708 503
rect 1908 497 1948 503
rect 2036 497 2236 503
rect 1044 477 1068 483
rect 1140 477 1180 483
rect 1620 477 1660 483
rect 1732 477 1756 483
rect 1924 477 2188 483
rect 1364 457 1468 463
rect 1508 457 1708 463
rect 2084 457 2140 463
rect 1140 437 1644 443
rect 2116 437 2156 443
rect 884 417 908 423
rect 616 414 664 416
rect 616 406 620 414
rect 630 406 636 414
rect 644 406 650 414
rect 660 406 664 414
rect 616 404 664 406
rect 1444 377 1836 383
rect 116 357 444 363
rect 468 357 492 363
rect 1092 357 1212 363
rect 1780 357 1804 363
rect 1828 357 1852 363
rect 164 337 332 343
rect 340 337 732 343
rect 820 337 844 343
rect 1012 337 1068 343
rect 1764 337 2092 343
rect 356 317 428 323
rect 596 317 796 323
rect 948 317 972 323
rect 1252 317 1276 323
rect 1604 317 1788 323
rect 2148 317 2220 323
rect 212 297 300 303
rect 308 297 380 303
rect 420 297 444 303
rect 1076 297 1164 303
rect 1220 297 1324 303
rect 1380 297 1420 303
rect 1428 297 1452 303
rect 1492 297 1772 303
rect 1780 297 1804 303
rect 1892 297 1980 303
rect 2068 297 2252 303
rect 2260 297 2291 303
rect 260 277 316 283
rect 324 277 524 283
rect 548 277 556 283
rect 1060 277 1116 283
rect 1268 277 1308 283
rect 1412 277 1484 283
rect 1524 277 1676 283
rect 1940 277 2028 283
rect 2100 277 2124 283
rect 244 257 380 263
rect 964 257 1148 263
rect 1652 257 1740 263
rect 1924 257 1948 263
rect 868 237 908 243
rect 948 237 1068 243
rect 1092 237 1276 243
rect 1300 237 1324 243
rect 1364 237 1436 243
rect 724 217 908 223
rect 1236 217 1292 223
rect 1576 214 1624 216
rect 1576 206 1580 214
rect 1590 206 1596 214
rect 1604 206 1610 214
rect 1620 206 1624 214
rect 1576 204 1624 206
rect 2132 197 2188 203
rect 196 177 524 183
rect 564 177 716 183
rect 2116 177 2140 183
rect 420 157 572 163
rect 740 157 764 163
rect 772 157 876 163
rect 1332 157 1356 163
rect 1460 157 1580 163
rect 1668 157 1900 163
rect 2052 157 2108 163
rect 68 137 108 143
rect 292 137 316 143
rect 324 137 364 143
rect 372 137 476 143
rect 484 137 540 143
rect 548 137 588 143
rect 596 137 684 143
rect 852 137 892 143
rect 900 137 924 143
rect 932 137 956 143
rect 1140 137 1212 143
rect 1316 137 1372 143
rect 1380 137 1532 143
rect 1700 137 1740 143
rect 1748 137 1788 143
rect 1796 137 1852 143
rect 1860 137 1916 143
rect 1956 137 2012 143
rect 260 117 428 123
rect 436 117 476 123
rect 516 117 524 123
rect 532 117 780 123
rect 1348 117 1372 123
rect 1716 117 1724 123
rect 1732 117 1772 123
rect 1780 117 1884 123
rect 1908 117 1996 123
rect 2164 117 2188 123
rect -19 97 12 103
rect 164 97 188 103
rect 340 97 444 103
rect 452 97 620 103
rect 628 97 700 103
rect 788 97 812 103
rect 820 97 860 103
rect 868 97 940 103
rect 1108 97 1180 103
rect 1188 97 1244 103
rect 1396 97 1532 103
rect 2020 97 2060 103
rect 2132 97 2172 103
rect 2260 97 2291 103
rect 244 77 348 83
rect 1860 77 1980 83
rect 2004 77 2028 83
rect 616 14 664 16
rect 616 6 620 14
rect 630 6 636 14
rect 644 6 650 14
rect 660 6 664 14
rect 616 4 664 6
<< m4contact >>
rect 620 1606 622 1614
rect 622 1606 628 1614
rect 636 1606 644 1614
rect 652 1606 658 1614
rect 658 1606 660 1614
rect 972 1596 980 1604
rect 1644 1516 1652 1524
rect 2092 1476 2100 1484
rect 1580 1406 1582 1414
rect 1582 1406 1588 1414
rect 1596 1406 1604 1414
rect 1612 1406 1618 1414
rect 1618 1406 1620 1414
rect 972 1356 980 1364
rect 620 1206 622 1214
rect 622 1206 628 1214
rect 636 1206 644 1214
rect 652 1206 658 1214
rect 658 1206 660 1214
rect 1292 1036 1300 1044
rect 1580 1006 1582 1014
rect 1582 1006 1588 1014
rect 1596 1006 1604 1014
rect 1612 1006 1618 1014
rect 1618 1006 1620 1014
rect 2172 996 2180 1004
rect 620 806 622 814
rect 622 806 628 814
rect 636 806 644 814
rect 652 806 658 814
rect 658 806 660 814
rect 1308 716 1316 724
rect 1372 696 1380 704
rect 1308 636 1316 644
rect 1372 616 1380 624
rect 1580 606 1582 614
rect 1582 606 1588 614
rect 1596 606 1604 614
rect 1612 606 1618 614
rect 1618 606 1620 614
rect 2108 596 2116 604
rect 1292 576 1300 584
rect 2092 576 2100 584
rect 1964 556 1972 564
rect 1228 516 1236 524
rect 1964 496 1972 504
rect 1644 436 1652 444
rect 2108 436 2116 444
rect 620 406 622 414
rect 622 406 628 414
rect 636 406 644 414
rect 652 406 658 414
rect 658 406 660 414
rect 1436 396 1444 404
rect 556 276 564 284
rect 2092 276 2100 284
rect 2172 276 2180 284
rect 1324 236 1332 244
rect 1580 206 1582 214
rect 1582 206 1588 214
rect 1596 206 1604 214
rect 1612 206 1618 214
rect 1618 206 1620 214
rect 1324 96 1332 104
rect 1436 36 1444 44
rect 556 16 564 24
rect 1228 16 1236 24
rect 620 6 622 14
rect 622 6 628 14
rect 636 6 644 14
rect 652 6 658 14
rect 658 6 660 14
<< metal4 >>
rect 616 1614 664 1640
rect 616 1606 620 1614
rect 628 1606 636 1614
rect 644 1606 652 1614
rect 660 1606 664 1614
rect 616 1214 664 1606
rect 973 1364 979 1596
rect 1576 1414 1624 1640
rect 1576 1406 1580 1414
rect 1588 1406 1596 1414
rect 1604 1406 1612 1414
rect 1620 1406 1624 1414
rect 616 1206 620 1214
rect 628 1206 636 1214
rect 644 1206 652 1214
rect 660 1206 664 1214
rect 616 814 664 1206
rect 616 806 620 814
rect 628 806 636 814
rect 644 806 652 814
rect 660 806 664 814
rect 616 414 664 806
rect 1293 584 1299 1036
rect 1576 1014 1624 1406
rect 1576 1006 1580 1014
rect 1588 1006 1596 1014
rect 1604 1006 1612 1014
rect 1620 1006 1624 1014
rect 1309 644 1315 716
rect 1373 624 1379 696
rect 1576 614 1624 1006
rect 1576 606 1580 614
rect 1588 606 1596 614
rect 1604 606 1612 614
rect 1620 606 1624 614
rect 616 406 620 414
rect 628 406 636 414
rect 644 406 652 414
rect 660 406 664 414
rect 557 24 563 276
rect 616 14 664 406
rect 1229 24 1235 516
rect 1325 104 1331 236
rect 1437 44 1443 396
rect 1576 214 1624 606
rect 1645 444 1651 1516
rect 2093 584 2099 1476
rect 1965 504 1971 556
rect 2093 284 2099 576
rect 2109 444 2115 596
rect 2173 284 2179 996
rect 1576 206 1580 214
rect 1588 206 1596 214
rect 1604 206 1612 214
rect 1620 206 1624 214
rect 616 6 620 14
rect 628 6 636 14
rect 644 6 652 14
rect 660 6 664 14
rect 616 -40 664 6
rect 1576 -40 1624 206
use BUFX2  BUFX2_21
timestamp 1586568500
transform -1 0 56 0 1 1410
box -4 -6 52 206
use OR2X2  OR2X2_26
timestamp 1586568500
transform 1 0 56 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_66
timestamp 1586568500
transform 1 0 120 0 1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_26
timestamp 1586568500
transform -1 0 216 0 1 1410
box -4 -6 52 206
use AND2X2  AND2X2_26
timestamp 1586568500
transform 1 0 216 0 1 1410
box -4 -6 68 206
use OR2X2  OR2X2_28
timestamp 1586568500
transform -1 0 344 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_70
timestamp 1586568500
transform 1 0 344 0 1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_28
timestamp 1586568500
transform -1 0 456 0 1 1410
box -4 -6 68 206
use BUFX2  BUFX2_20
timestamp 1586568500
transform -1 0 504 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_71
timestamp 1586568500
transform -1 0 552 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_4
timestamp 1586568500
transform 1 0 552 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_60
timestamp 1586568500
transform 1 0 600 0 1 1410
box -4 -6 52 206
use FILL  FILL_7_0_0
timestamp 1586568500
transform 1 0 648 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_1
timestamp 1586568500
transform 1 0 664 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_2
timestamp 1586568500
transform 1 0 680 0 1 1410
box -4 -6 20 206
use OR2X2  OR2X2_19
timestamp 1586568500
transform 1 0 696 0 1 1410
box -4 -6 68 206
use AND2X2  AND2X2_19
timestamp 1586568500
transform 1 0 760 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_52
timestamp 1586568500
transform 1 0 824 0 1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_19
timestamp 1586568500
transform -1 0 920 0 1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_19
timestamp 1586568500
transform -1 0 984 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_53
timestamp 1586568500
transform -1 0 1048 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_34
timestamp 1586568500
transform -1 0 1080 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_52
timestamp 1586568500
transform 1 0 1080 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_53
timestamp 1586568500
transform 1 0 1144 0 1 1410
box -4 -6 52 206
use INVX1  INVX1_29
timestamp 1586568500
transform 1 0 1192 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_45
timestamp 1586568500
transform 1 0 1224 0 1 1410
box -4 -6 68 206
use BUFX2  BUFX2_15
timestamp 1586568500
transform 1 0 1288 0 1 1410
box -4 -6 52 206
use AND2X2  AND2X2_20
timestamp 1586568500
transform 1 0 1336 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_54
timestamp 1586568500
transform 1 0 1400 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_19
timestamp 1586568500
transform -1 0 1496 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_3
timestamp 1586568500
transform 1 0 1496 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_69
timestamp 1586568500
transform -1 0 1592 0 1 1410
box -4 -6 52 206
use FILL  FILL_7_1_0
timestamp 1586568500
transform -1 0 1608 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_1
timestamp 1586568500
transform -1 0 1624 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_2
timestamp 1586568500
transform -1 0 1640 0 1 1410
box -4 -6 20 206
use OAI21X1  OAI21X1_68
timestamp 1586568500
transform -1 0 1704 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_42
timestamp 1586568500
transform 1 0 1704 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_69
timestamp 1586568500
transform 1 0 1736 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_27
timestamp 1586568500
transform 1 0 1800 0 1 1410
box -4 -6 68 206
use AND2X2  AND2X2_27
timestamp 1586568500
transform -1 0 1928 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_68
timestamp 1586568500
transform -1 0 1976 0 1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_27
timestamp 1586568500
transform 1 0 1976 0 1 1410
box -4 -6 52 206
use OR2X2  OR2X2_27
timestamp 1586568500
transform 1 0 2024 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_23
timestamp 1586568500
transform 1 0 2088 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_23
timestamp 1586568500
transform -1 0 2200 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_15
timestamp 1586568500
transform -1 0 2232 0 1 1410
box -4 -6 36 206
use FILL  FILL_8_1
timestamp 1586568500
transform 1 0 2232 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_2
timestamp 1586568500
transform 1 0 2248 0 1 1410
box -4 -6 20 206
use BUFX2  BUFX2_5
timestamp 1586568500
transform -1 0 56 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_67
timestamp 1586568500
transform -1 0 104 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_26
timestamp 1586568500
transform -1 0 168 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_67
timestamp 1586568500
transform -1 0 232 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_66
timestamp 1586568500
transform 1 0 232 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_41
timestamp 1586568500
transform -1 0 328 0 -1 1410
box -4 -6 36 206
use NOR2X1  NOR2X1_28
timestamp 1586568500
transform -1 0 376 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_71
timestamp 1586568500
transform -1 0 440 0 -1 1410
box -4 -6 68 206
use AND2X2  AND2X2_28
timestamp 1586568500
transform 1 0 440 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_70
timestamp 1586568500
transform 1 0 504 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_43
timestamp 1586568500
transform -1 0 600 0 -1 1410
box -4 -6 36 206
use FILL  FILL_6_0_0
timestamp 1586568500
transform 1 0 600 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_1
timestamp 1586568500
transform 1 0 616 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_2
timestamp 1586568500
transform 1 0 632 0 -1 1410
box -4 -6 20 206
use AND2X2  AND2X2_23
timestamp 1586568500
transform 1 0 648 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_23
timestamp 1586568500
transform 1 0 712 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_60
timestamp 1586568500
transform 1 0 760 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_61
timestamp 1586568500
transform 1 0 824 0 -1 1410
box -4 -6 52 206
use OR2X2  OR2X2_23
timestamp 1586568500
transform -1 0 936 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_17
timestamp 1586568500
transform 1 0 936 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_32
timestamp 1586568500
transform 1 0 984 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_49
timestamp 1586568500
transform 1 0 1016 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_17
timestamp 1586568500
transform 1 0 1080 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_48
timestamp 1586568500
transform -1 0 1192 0 -1 1410
box -4 -6 52 206
use OR2X2  OR2X2_17
timestamp 1586568500
transform 1 0 1192 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_45
timestamp 1586568500
transform -1 0 1304 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_35
timestamp 1586568500
transform 1 0 1304 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_54
timestamp 1586568500
transform -1 0 1400 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_55
timestamp 1586568500
transform 1 0 1400 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_20
timestamp 1586568500
transform 1 0 1464 0 -1 1410
box -4 -6 52 206
use OR2X2  OR2X2_20
timestamp 1586568500
transform 1 0 1512 0 -1 1410
box -4 -6 68 206
use FILL  FILL_6_1_0
timestamp 1586568500
transform 1 0 1576 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_1
timestamp 1586568500
transform 1 0 1592 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_2
timestamp 1586568500
transform 1 0 1608 0 -1 1410
box -4 -6 20 206
use NAND3X1  NAND3X1_20
timestamp 1586568500
transform 1 0 1624 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_55
timestamp 1586568500
transform 1 0 1688 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_30
timestamp 1586568500
transform 1 0 1736 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_46
timestamp 1586568500
transform 1 0 1768 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_16
timestamp 1586568500
transform 1 0 1832 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_35
timestamp 1586568500
transform -1 0 1944 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_36
timestamp 1586568500
transform 1 0 1944 0 -1 1410
box -4 -6 52 206
use AND2X2  AND2X2_13
timestamp 1586568500
transform -1 0 2056 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_9
timestamp 1586568500
transform -1 0 2104 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_27
timestamp 1586568500
transform -1 0 2168 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_28
timestamp 1586568500
transform 1 0 2168 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_10
timestamp 1586568500
transform 1 0 2216 0 -1 1410
box -4 -6 52 206
use AND2X2  AND2X2_2
timestamp 1586568500
transform -1 0 72 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_2
timestamp 1586568500
transform 1 0 72 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_8
timestamp 1586568500
transform 1 0 120 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_9
timestamp 1586568500
transform 1 0 184 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_7
timestamp 1586568500
transform 1 0 232 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_9
timestamp 1586568500
transform 1 0 264 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_2
timestamp 1586568500
transform 1 0 328 0 1 1010
box -4 -6 68 206
use OR2X2  OR2X2_2
timestamp 1586568500
transform -1 0 456 0 1 1010
box -4 -6 68 206
use AND2X2  AND2X2_6
timestamp 1586568500
transform 1 0 456 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_16
timestamp 1586568500
transform -1 0 568 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_1
timestamp 1586568500
transform 1 0 568 0 1 1010
box -4 -6 36 206
use FILL  FILL_5_0_0
timestamp 1586568500
transform 1 0 600 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_1
timestamp 1586568500
transform 1 0 616 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_2
timestamp 1586568500
transform 1 0 632 0 1 1010
box -4 -6 20 206
use OAI21X1  OAI21X1_1
timestamp 1586568500
transform 1 0 648 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_61
timestamp 1586568500
transform -1 0 776 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_38
timestamp 1586568500
transform -1 0 808 0 1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_23
timestamp 1586568500
transform 1 0 808 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_56
timestamp 1586568500
transform -1 0 920 0 1 1010
box -4 -6 52 206
use AND2X2  AND2X2_17
timestamp 1586568500
transform 1 0 920 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_48
timestamp 1586568500
transform 1 0 984 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_49
timestamp 1586568500
transform 1 0 1048 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_28
timestamp 1586568500
transform 1 0 1096 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_44
timestamp 1586568500
transform 1 0 1128 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_14
timestamp 1586568500
transform 1 0 1192 0 1 1010
box -4 -6 52 206
use AND2X2  AND2X2_24
timestamp 1586568500
transform -1 0 1304 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_24
timestamp 1586568500
transform 1 0 1304 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_62
timestamp 1586568500
transform 1 0 1352 0 1 1010
box -4 -6 52 206
use OR2X2  OR2X2_24
timestamp 1586568500
transform 1 0 1400 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_46
timestamp 1586568500
transform 1 0 1464 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_39
timestamp 1586568500
transform 1 0 1512 0 1 1010
box -4 -6 52 206
use FILL  FILL_5_1_0
timestamp 1586568500
transform 1 0 1560 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_1
timestamp 1586568500
transform 1 0 1576 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_2
timestamp 1586568500
transform 1 0 1592 0 1 1010
box -4 -6 20 206
use AND2X2  AND2X2_15
timestamp 1586568500
transform 1 0 1608 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_23
timestamp 1586568500
transform 1 0 1672 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_36
timestamp 1586568500
transform 1 0 1704 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_13
timestamp 1586568500
transform 1 0 1768 0 1 1010
box -4 -6 68 206
use OR2X2  OR2X2_13
timestamp 1586568500
transform -1 0 1896 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_35
timestamp 1586568500
transform -1 0 1944 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_13
timestamp 1586568500
transform 1 0 1944 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_28
timestamp 1586568500
transform 1 0 1992 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_27
timestamp 1586568500
transform -1 0 2104 0 1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_9
timestamp 1586568500
transform 1 0 2104 0 1 1010
box -4 -6 68 206
use OR2X2  OR2X2_9
timestamp 1586568500
transform -1 0 2232 0 1 1010
box -4 -6 68 206
use FILL  FILL_6_1
timestamp 1586568500
transform 1 0 2232 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_2
timestamp 1586568500
transform 1 0 2248 0 1 1010
box -4 -6 20 206
use BUFX2  BUFX2_9
timestamp 1586568500
transform -1 0 56 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_5
timestamp 1586568500
transform 1 0 56 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_5
timestamp 1586568500
transform -1 0 152 0 -1 1010
box -4 -6 36 206
use NAND2X1  NAND2X1_5
timestamp 1586568500
transform 1 0 152 0 -1 1010
box -4 -6 52 206
use OR2X2  OR2X2_6
timestamp 1586568500
transform 1 0 200 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_8
timestamp 1586568500
transform -1 0 312 0 -1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_6
timestamp 1586568500
transform -1 0 376 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_17
timestamp 1586568500
transform -1 0 424 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_11
timestamp 1586568500
transform -1 0 456 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_16
timestamp 1586568500
transform -1 0 520 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_6
timestamp 1586568500
transform -1 0 568 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_17
timestamp 1586568500
transform 1 0 568 0 -1 1010
box -4 -6 68 206
use FILL  FILL_4_0_0
timestamp 1586568500
transform 1 0 632 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_1
timestamp 1586568500
transform 1 0 648 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_2
timestamp 1586568500
transform 1 0 664 0 -1 1010
box -4 -6 20 206
use NAND2X1  NAND2X1_1
timestamp 1586568500
transform 1 0 680 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_36
timestamp 1586568500
transform -1 0 760 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_57
timestamp 1586568500
transform 1 0 760 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_21
timestamp 1586568500
transform 1 0 824 0 -1 1010
box -4 -6 68 206
use OR2X2  OR2X2_21
timestamp 1586568500
transform -1 0 952 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_21
timestamp 1586568500
transform -1 0 1000 0 -1 1010
box -4 -6 52 206
use AND2X2  AND2X2_21
timestamp 1586568500
transform 1 0 1000 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_56
timestamp 1586568500
transform 1 0 1064 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_57
timestamp 1586568500
transform 1 0 1128 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_44
timestamp 1586568500
transform 1 0 1176 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_62
timestamp 1586568500
transform -1 0 1288 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_39
timestamp 1586568500
transform 1 0 1288 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_63
timestamp 1586568500
transform 1 0 1320 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_24
timestamp 1586568500
transform 1 0 1384 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_63
timestamp 1586568500
transform 1 0 1448 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_40
timestamp 1586568500
transform -1 0 1560 0 -1 1010
box -4 -6 68 206
use FILL  FILL_4_1_0
timestamp 1586568500
transform 1 0 1560 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_1
timestamp 1586568500
transform 1 0 1576 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_2
timestamp 1586568500
transform 1 0 1592 0 -1 1010
box -4 -6 20 206
use NOR2X1  NOR2X1_15
timestamp 1586568500
transform 1 0 1608 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_39
timestamp 1586568500
transform 1 0 1656 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_25
timestamp 1586568500
transform 1 0 1720 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_15
timestamp 1586568500
transform 1 0 1752 0 -1 1010
box -4 -6 68 206
use OR2X2  OR2X2_15
timestamp 1586568500
transform -1 0 1880 0 -1 1010
box -4 -6 68 206
use AND2X2  AND2X2_11
timestamp 1586568500
transform 1 0 1880 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_11
timestamp 1586568500
transform -1 0 1992 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_19
timestamp 1586568500
transform 1 0 1992 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_31
timestamp 1586568500
transform 1 0 2024 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_21
timestamp 1586568500
transform 1 0 2088 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_11
timestamp 1586568500
transform 1 0 2120 0 -1 1010
box -4 -6 68 206
use OR2X2  OR2X2_11
timestamp 1586568500
transform -1 0 2248 0 -1 1010
box -4 -6 68 206
use FILL  FILL_5_1
timestamp 1586568500
transform -1 0 2264 0 -1 1010
box -4 -6 20 206
use OR2X2  OR2X2_4
timestamp 1586568500
transform 1 0 8 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_12
timestamp 1586568500
transform 1 0 72 0 1 610
box -4 -6 52 206
use NAND3X1  NAND3X1_4
timestamp 1586568500
transform -1 0 184 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_13
timestamp 1586568500
transform -1 0 232 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_13
timestamp 1586568500
transform -1 0 296 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_4
timestamp 1586568500
transform -1 0 344 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_20
timestamp 1586568500
transform 1 0 344 0 1 610
box -4 -6 52 206
use OR2X2  OR2X2_8
timestamp 1586568500
transform 1 0 392 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_21
timestamp 1586568500
transform -1 0 504 0 1 610
box -4 -6 52 206
use NAND3X1  NAND3X1_8
timestamp 1586568500
transform -1 0 568 0 1 610
box -4 -6 68 206
use INVX1  INVX1_13
timestamp 1586568500
transform 1 0 568 0 1 610
box -4 -6 36 206
use FILL  FILL_3_0_0
timestamp 1586568500
transform 1 0 600 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_1
timestamp 1586568500
transform 1 0 616 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_2
timestamp 1586568500
transform 1 0 632 0 1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_21
timestamp 1586568500
transform 1 0 648 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_2
timestamp 1586568500
transform -1 0 760 0 1 610
box -4 -6 52 206
use INVX1  INVX1_10
timestamp 1586568500
transform 1 0 760 0 1 610
box -4 -6 36 206
use NAND3X1  NAND3X1_5
timestamp 1586568500
transform -1 0 856 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_15
timestamp 1586568500
transform -1 0 904 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_14
timestamp 1586568500
transform 1 0 904 0 1 610
box -4 -6 68 206
use OR2X2  OR2X2_22
timestamp 1586568500
transform 1 0 968 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_50
timestamp 1586568500
transform 1 0 1032 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_58
timestamp 1586568500
transform -1 0 1128 0 1 610
box -4 -6 52 206
use NAND3X1  NAND3X1_22
timestamp 1586568500
transform -1 0 1192 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_59
timestamp 1586568500
transform -1 0 1256 0 1 610
box -4 -6 68 206
use INVX1  INVX1_37
timestamp 1586568500
transform -1 0 1288 0 1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_59
timestamp 1586568500
transform -1 0 1336 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_58
timestamp 1586568500
transform -1 0 1400 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_22
timestamp 1586568500
transform -1 0 1448 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_43
timestamp 1586568500
transform 1 0 1448 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_41
timestamp 1586568500
transform -1 0 1560 0 1 610
box -4 -6 68 206
use FILL  FILL_3_1_0
timestamp 1586568500
transform -1 0 1576 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_1
timestamp 1586568500
transform -1 0 1592 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_2
timestamp 1586568500
transform -1 0 1608 0 1 610
box -4 -6 20 206
use AND2X2  AND2X2_16
timestamp 1586568500
transform -1 0 1672 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_16
timestamp 1586568500
transform -1 0 1720 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_41
timestamp 1586568500
transform -1 0 1768 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_40
timestamp 1586568500
transform 1 0 1768 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_24
timestamp 1586568500
transform -1 0 1864 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_24
timestamp 1586568500
transform -1 0 1928 0 1 610
box -4 -6 68 206
use INVX1  INVX1_16
timestamp 1586568500
transform -1 0 1960 0 1 610
box -4 -6 36 206
use BUFX2  BUFX2_11
timestamp 1586568500
transform 1 0 1960 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_32
timestamp 1586568500
transform -1 0 2056 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_32
timestamp 1586568500
transform 1 0 2056 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_33
timestamp 1586568500
transform 1 0 2120 0 1 610
box -4 -6 52 206
use AND2X2  AND2X2_9
timestamp 1586568500
transform -1 0 2232 0 1 610
box -4 -6 68 206
use FILL  FILL_4_1
timestamp 1586568500
transform 1 0 2232 0 1 610
box -4 -6 20 206
use FILL  FILL_4_2
timestamp 1586568500
transform 1 0 2248 0 1 610
box -4 -6 20 206
use BUFX2  BUFX2_8
timestamp 1586568500
transform -1 0 56 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_4
timestamp 1586568500
transform 1 0 56 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_4
timestamp 1586568500
transform 1 0 120 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_4
timestamp 1586568500
transform -1 0 200 0 -1 610
box -4 -6 36 206
use INVX1  INVX1_9
timestamp 1586568500
transform -1 0 232 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_12
timestamp 1586568500
transform -1 0 296 0 -1 610
box -4 -6 68 206
use AND2X2  AND2X2_4
timestamp 1586568500
transform -1 0 360 0 -1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_8
timestamp 1586568500
transform -1 0 408 0 -1 610
box -4 -6 52 206
use AND2X2  AND2X2_8
timestamp 1586568500
transform 1 0 408 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_20
timestamp 1586568500
transform 1 0 472 0 -1 610
box -4 -6 68 206
use BUFX2  BUFX2_6
timestamp 1586568500
transform -1 0 584 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_2
timestamp 1586568500
transform 1 0 584 0 -1 610
box -4 -6 68 206
use FILL  FILL_2_0_0
timestamp 1586568500
transform -1 0 664 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1586568500
transform -1 0 680 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_2
timestamp 1586568500
transform -1 0 696 0 -1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_15
timestamp 1586568500
transform -1 0 760 0 -1 610
box -4 -6 68 206
use OR2X2  OR2X2_5
timestamp 1586568500
transform -1 0 824 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_14
timestamp 1586568500
transform -1 0 872 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_5
timestamp 1586568500
transform 1 0 872 0 -1 610
box -4 -6 52 206
use AND2X2  AND2X2_5
timestamp 1586568500
transform 1 0 920 0 -1 610
box -4 -6 68 206
use OR2X2  OR2X2_18
timestamp 1586568500
transform 1 0 984 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_18
timestamp 1586568500
transform -1 0 1112 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_51
timestamp 1586568500
transform -1 0 1176 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_33
timestamp 1586568500
transform -1 0 1208 0 -1 610
box -4 -6 36 206
use NOR2X1  NOR2X1_18
timestamp 1586568500
transform 1 0 1208 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_50
timestamp 1586568500
transform 1 0 1256 0 -1 610
box -4 -6 68 206
use AND2X2  AND2X2_18
timestamp 1586568500
transform -1 0 1384 0 -1 610
box -4 -6 68 206
use AND2X2  AND2X2_22
timestamp 1586568500
transform -1 0 1448 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_25
timestamp 1586568500
transform 1 0 1448 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_42
timestamp 1586568500
transform -1 0 1544 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_26
timestamp 1586568500
transform 1 0 1544 0 -1 610
box -4 -6 36 206
use FILL  FILL_2_1_0
timestamp 1586568500
transform 1 0 1576 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1586568500
transform 1 0 1592 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_2
timestamp 1586568500
transform 1 0 1608 0 -1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_42
timestamp 1586568500
transform 1 0 1624 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_16
timestamp 1586568500
transform 1 0 1688 0 -1 610
box -4 -6 68 206
use OR2X2  OR2X2_16
timestamp 1586568500
transform -1 0 1816 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_17
timestamp 1586568500
transform 1 0 1816 0 -1 610
box -4 -6 36 206
use AND2X2  AND2X2_12
timestamp 1586568500
transform 1 0 1848 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_34
timestamp 1586568500
transform -1 0 1960 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_33
timestamp 1586568500
transform -1 0 2024 0 -1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_12
timestamp 1586568500
transform -1 0 2072 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_22
timestamp 1586568500
transform 1 0 2072 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_34
timestamp 1586568500
transform 1 0 2104 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_12
timestamp 1586568500
transform 1 0 2168 0 -1 610
box -4 -6 68 206
use FILL  FILL_3_1
timestamp 1586568500
transform -1 0 2248 0 -1 610
box -4 -6 20 206
use FILL  FILL_3_2
timestamp 1586568500
transform -1 0 2264 0 -1 610
box -4 -6 20 206
use BUFX2  BUFX2_22
timestamp 1586568500
transform -1 0 56 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_3
timestamp 1586568500
transform 1 0 56 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_19
timestamp 1586568500
transform -1 0 152 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_18
timestamp 1586568500
transform -1 0 216 0 1 210
box -4 -6 68 206
use AND2X2  AND2X2_7
timestamp 1586568500
transform -1 0 280 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_7
timestamp 1586568500
transform 1 0 280 0 1 210
box -4 -6 52 206
use INVX1  INVX1_12
timestamp 1586568500
transform 1 0 328 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_19
timestamp 1586568500
transform 1 0 360 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_7
timestamp 1586568500
transform 1 0 424 0 1 210
box -4 -6 68 206
use OR2X2  OR2X2_7
timestamp 1586568500
transform -1 0 552 0 1 210
box -4 -6 68 206
use INVX1  INVX1_2
timestamp 1586568500
transform -1 0 584 0 1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_7
timestamp 1586568500
transform -1 0 632 0 1 210
box -4 -6 52 206
use FILL  FILL_1_0_0
timestamp 1586568500
transform -1 0 648 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_1
timestamp 1586568500
transform -1 0 664 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_2
timestamp 1586568500
transform -1 0 680 0 1 210
box -4 -6 20 206
use OAI21X1  OAI21X1_6
timestamp 1586568500
transform -1 0 744 0 1 210
box -4 -6 68 206
use INVX1  INVX1_6
timestamp 1586568500
transform 1 0 744 0 1 210
box -4 -6 36 206
use NAND3X1  NAND3X1_1
timestamp 1586568500
transform 1 0 776 0 1 210
box -4 -6 68 206
use OR2X2  OR2X2_1
timestamp 1586568500
transform -1 0 904 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_64
timestamp 1586568500
transform -1 0 968 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_65
timestamp 1586568500
transform 1 0 968 0 1 210
box -4 -6 52 206
use INVX1  INVX1_40
timestamp 1586568500
transform 1 0 1016 0 1 210
box -4 -6 36 206
use NAND3X1  NAND3X1_25
timestamp 1586568500
transform 1 0 1048 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_65
timestamp 1586568500
transform 1 0 1112 0 1 210
box -4 -6 68 206
use INVX1  INVX1_27
timestamp 1586568500
transform 1 0 1176 0 1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_51
timestamp 1586568500
transform -1 0 1256 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_47
timestamp 1586568500
transform 1 0 1256 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_43
timestamp 1586568500
transform 1 0 1304 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_22
timestamp 1586568500
transform -1 0 1416 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_25
timestamp 1586568500
transform 1 0 1416 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_38
timestamp 1586568500
transform -1 0 1544 0 1 210
box -4 -6 68 206
use INVX1  INVX1_24
timestamp 1586568500
transform -1 0 1576 0 1 210
box -4 -6 36 206
use FILL  FILL_1_1_0
timestamp 1586568500
transform -1 0 1592 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_1
timestamp 1586568500
transform -1 0 1608 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_2
timestamp 1586568500
transform -1 0 1624 0 1 210
box -4 -6 20 206
use OAI21X1  OAI21X1_37
timestamp 1586568500
transform -1 0 1688 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_14
timestamp 1586568500
transform -1 0 1736 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_38
timestamp 1586568500
transform 1 0 1736 0 1 210
box -4 -6 52 206
use NAND3X1  NAND3X1_14
timestamp 1586568500
transform 1 0 1784 0 1 210
box -4 -6 68 206
use OR2X2  OR2X2_14
timestamp 1586568500
transform -1 0 1912 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_10
timestamp 1586568500
transform -1 0 1960 0 1 210
box -4 -6 52 206
use AND2X2  AND2X2_10
timestamp 1586568500
transform 1 0 1960 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_29
timestamp 1586568500
transform 1 0 2024 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_26
timestamp 1586568500
transform -1 0 2136 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_31
timestamp 1586568500
transform -1 0 2184 0 1 210
box -4 -6 52 206
use OR2X2  OR2X2_12
timestamp 1586568500
transform -1 0 2248 0 1 210
box -4 -6 68 206
use FILL  FILL_2_1
timestamp 1586568500
transform 1 0 2248 0 1 210
box -4 -6 20 206
use BUFX2  BUFX2_7
timestamp 1586568500
transform -1 0 56 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_3
timestamp 1586568500
transform -1 0 120 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_3
timestamp 1586568500
transform -1 0 152 0 -1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_11
timestamp 1586568500
transform -1 0 200 0 -1 210
box -4 -6 52 206
use NAND3X1  NAND3X1_3
timestamp 1586568500
transform -1 0 264 0 -1 210
box -4 -6 68 206
use OR2X2  OR2X2_3
timestamp 1586568500
transform -1 0 328 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_10
timestamp 1586568500
transform -1 0 376 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_11
timestamp 1586568500
transform -1 0 440 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_18
timestamp 1586568500
transform -1 0 488 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_8
timestamp 1586568500
transform -1 0 520 0 -1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_10
timestamp 1586568500
transform -1 0 584 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_3
timestamp 1586568500
transform 1 0 584 0 -1 210
box -4 -6 52 206
use FILL  FILL_0_0_0
timestamp 1586568500
transform 1 0 632 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1586568500
transform 1 0 648 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_2
timestamp 1586568500
transform 1 0 664 0 -1 210
box -4 -6 20 206
use AND2X2  AND2X2_3
timestamp 1586568500
transform 1 0 680 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_7
timestamp 1586568500
transform 1 0 744 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_6
timestamp 1586568500
transform -1 0 856 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_1
timestamp 1586568500
transform -1 0 904 0 -1 210
box -4 -6 52 206
use AND2X2  AND2X2_1
timestamp 1586568500
transform -1 0 968 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_2
timestamp 1586568500
transform -1 0 1016 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_18
timestamp 1586568500
transform 1 0 1016 0 -1 210
box -4 -6 52 206
use AND2X2  AND2X2_25
timestamp 1586568500
transform -1 0 1128 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_25
timestamp 1586568500
transform 1 0 1128 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_64
timestamp 1586568500
transform -1 0 1224 0 -1 210
box -4 -6 52 206
use OR2X2  OR2X2_25
timestamp 1586568500
transform 1 0 1224 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_31
timestamp 1586568500
transform 1 0 1288 0 -1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_47
timestamp 1586568500
transform -1 0 1384 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_17
timestamp 1586568500
transform 1 0 1384 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_1
timestamp 1586568500
transform 1 0 1432 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_12
timestamp 1586568500
transform 1 0 1480 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_22
timestamp 1586568500
transform -1 0 1592 0 -1 210
box -4 -6 68 206
use FILL  FILL_0_1_0
timestamp 1586568500
transform -1 0 1608 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1586568500
transform -1 0 1624 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_2
timestamp 1586568500
transform -1 0 1640 0 -1 210
box -4 -6 20 206
use INVX1  INVX1_14
timestamp 1586568500
transform -1 0 1672 0 -1 210
box -4 -6 36 206
use AND2X2  AND2X2_14
timestamp 1586568500
transform -1 0 1736 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_37
timestamp 1586568500
transform 1 0 1736 0 -1 210
box -4 -6 52 206
use OR2X2  OR2X2_10
timestamp 1586568500
transform 1 0 1784 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_29
timestamp 1586568500
transform 1 0 1848 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_30
timestamp 1586568500
transform -1 0 1960 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_10
timestamp 1586568500
transform -1 0 2024 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_30
timestamp 1586568500
transform -1 0 2072 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_20
timestamp 1586568500
transform -1 0 2104 0 -1 210
box -4 -6 36 206
use INVX1  INVX1_18
timestamp 1586568500
transform 1 0 2104 0 -1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_26
timestamp 1586568500
transform -1 0 2200 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_13
timestamp 1586568500
transform 1 0 2200 0 -1 210
box -4 -6 52 206
use FILL  FILL_1_1
timestamp 1586568500
transform -1 0 2264 0 -1 210
box -4 -6 20 206
<< labels >>
flabel metal4 s 616 -40 664 -16 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 1576 -40 1624 -16 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 1181 -23 1187 -17 7 FreeSans 24 270 0 0 i_add_term1[0]
port 2 nsew
flabel metal2 s 1965 1637 1971 1643 3 FreeSans 24 90 0 0 i_add_term1[1]
port 3 nsew
flabel metal2 s 397 1637 403 1643 3 FreeSans 24 90 0 0 i_add_term1[2]
port 4 nsew
flabel metal3 s -19 1537 -13 1543 7 FreeSans 24 0 0 0 i_add_term1[3]
port 5 nsew
flabel metal2 s 781 -23 787 -17 7 FreeSans 24 270 0 0 i_add_term1[4]
port 6 nsew
flabel metal2 s 445 -23 451 -17 7 FreeSans 24 270 0 0 i_add_term1[5]
port 7 nsew
flabel metal3 s -19 677 -13 683 7 FreeSans 24 0 0 0 i_add_term1[6]
port 8 nsew
flabel metal3 s -19 1137 -13 1143 7 FreeSans 24 0 0 0 i_add_term1[7]
port 9 nsew
flabel metal3 s 2285 917 2291 923 3 FreeSans 24 0 0 0 i_add_term1[8]
port 10 nsew
flabel metal3 s 2285 957 2291 963 3 FreeSans 24 0 0 0 i_add_term1[9]
port 11 nsew
flabel metal3 s 2285 517 2291 523 3 FreeSans 24 0 0 0 i_add_term1[10]
port 12 nsew
flabel metal2 s 1725 -23 1731 -17 7 FreeSans 24 270 0 0 i_add_term1[11]
port 13 nsew
flabel metal2 s 1213 1637 1219 1643 3 FreeSans 24 90 0 0 i_add_term1[12]
port 14 nsew
flabel metal2 s 669 1637 675 1643 3 FreeSans 24 90 0 0 i_add_term1[13]
port 15 nsew
flabel metal2 s 1437 1637 1443 1643 3 FreeSans 24 90 0 0 i_add_term1[14]
port 16 nsew
flabel metal2 s 1229 -23 1235 -17 7 FreeSans 24 270 0 0 i_add_term1[15]
port 17 nsew
flabel metal2 s 1117 -23 1123 -17 7 FreeSans 24 270 0 0 i_add_term2[0]
port 18 nsew
flabel metal2 s 1917 1637 1923 1643 3 FreeSans 24 90 0 0 i_add_term2[1]
port 19 nsew
flabel metal2 s 349 1637 355 1643 3 FreeSans 24 90 0 0 i_add_term2[2]
port 20 nsew
flabel metal3 s -19 1497 -13 1503 7 FreeSans 24 0 0 0 i_add_term2[3]
port 21 nsew
flabel metal2 s 941 -23 947 -17 7 FreeSans 24 270 0 0 i_add_term2[4]
port 22 nsew
flabel metal2 s 589 -23 595 -17 7 FreeSans 24 270 0 0 i_add_term2[5]
port 23 nsew
flabel metal3 s -19 717 -13 723 7 FreeSans 24 0 0 0 i_add_term2[6]
port 24 nsew
flabel metal3 s -19 1097 -13 1103 7 FreeSans 24 0 0 0 i_add_term2[7]
port 25 nsew
flabel metal3 s 2285 1117 2291 1123 3 FreeSans 24 0 0 0 i_add_term2[8]
port 26 nsew
flabel metal3 s 2285 997 2291 1003 3 FreeSans 24 0 0 0 i_add_term2[9]
port 27 nsew
flabel metal3 s 2285 297 2291 303 3 FreeSans 24 0 0 0 i_add_term2[10]
port 28 nsew
flabel metal2 s 1693 -23 1699 -17 7 FreeSans 24 270 0 0 i_add_term2[11]
port 29 nsew
flabel metal2 s 973 1637 979 1643 3 FreeSans 24 90 0 0 i_add_term2[12]
port 30 nsew
flabel metal2 s 717 1637 723 1643 3 FreeSans 24 90 0 0 i_add_term2[13]
port 31 nsew
flabel metal2 s 1373 1637 1379 1643 3 FreeSans 24 90 0 0 i_add_term2[14]
port 32 nsew
flabel metal2 s 1437 -23 1443 -17 7 FreeSans 24 270 0 0 i_add_term2[15]
port 33 nsew
flabel metal2 s 989 -23 995 -17 7 FreeSans 24 270 0 0 sum[0]
port 34 nsew
flabel metal2 s 1517 1637 1523 1643 3 FreeSans 24 90 0 0 sum[1]
port 35 nsew
flabel metal2 s 573 1637 579 1643 3 FreeSans 24 90 0 0 sum[2]
port 36 nsew
flabel metal3 s -19 1297 -13 1303 7 FreeSans 24 0 0 0 sum[3]
port 37 nsew
flabel metal2 s 557 -23 563 -17 7 FreeSans 24 270 0 0 sum[4]
port 38 nsew
flabel metal3 s -19 97 -13 103 7 FreeSans 24 0 0 0 sum[5]
port 39 nsew
flabel metal3 s -19 497 -13 503 7 FreeSans 24 0 0 0 sum[6]
port 40 nsew
flabel metal3 s -19 897 -13 903 7 FreeSans 24 0 0 0 sum[7]
port 41 nsew
flabel metal3 s 2285 1297 2291 1303 3 FreeSans 24 0 0 0 sum[8]
port 42 nsew
flabel metal3 s 2285 697 2291 703 3 FreeSans 24 0 0 0 sum[9]
port 43 nsew
flabel metal2 s 1501 -23 1507 -17 7 FreeSans 24 270 0 0 sum[10]
port 44 nsew
flabel metal3 s 2285 97 2291 103 3 FreeSans 24 0 0 0 sum[11]
port 45 nsew
flabel metal2 s 1245 1637 1251 1643 3 FreeSans 24 90 0 0 sum[12]
port 46 nsew
flabel metal2 s 1309 1637 1315 1643 3 FreeSans 24 90 0 0 sum[13]
port 47 nsew
flabel metal2 s 1853 1637 1859 1643 3 FreeSans 24 90 0 0 sum[14]
port 48 nsew
flabel metal2 s 1405 -23 1411 -17 7 FreeSans 24 270 0 0 sum[15]
port 49 nsew
flabel metal2 s 1469 -23 1475 -17 7 FreeSans 24 270 0 0 cout
port 50 nsew
<< end >>
