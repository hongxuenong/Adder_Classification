module csa_32bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [31:0] i_add_term1;
input [31:0] i_add_term2;
output [31:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

OAI21X1 OAI21X1_1 ( .A(_369_), .B(_366_), .C(_371_), .Y(_30__3_) );
INVX1 INVX1_1 ( .A(_31_), .Y(_373_) );
NAND2X1 NAND2X1_1 ( .A(_32_), .B(w_cout_5_), .Y(_374_) );
OAI21X1 OAI21X1_2 ( .A(w_cout_5_), .B(_373_), .C(_374_), .Y(w_cout_6_) );
INVX1 INVX1_2 ( .A(_33__0_), .Y(_375_) );
NAND2X1 NAND2X1_2 ( .A(_34__0_), .B(w_cout_5_), .Y(_376_) );
OAI21X1 OAI21X1_3 ( .A(w_cout_5_), .B(_375_), .C(_376_), .Y(_0__24_) );
INVX1 INVX1_3 ( .A(_33__1_), .Y(_377_) );
NAND2X1 NAND2X1_3 ( .A(w_cout_5_), .B(_34__1_), .Y(_378_) );
OAI21X1 OAI21X1_4 ( .A(w_cout_5_), .B(_377_), .C(_378_), .Y(_0__25_) );
INVX1 INVX1_4 ( .A(_33__2_), .Y(_379_) );
NAND2X1 NAND2X1_4 ( .A(w_cout_5_), .B(_34__2_), .Y(_380_) );
OAI21X1 OAI21X1_5 ( .A(w_cout_5_), .B(_379_), .C(_380_), .Y(_0__26_) );
INVX1 INVX1_5 ( .A(_33__3_), .Y(_381_) );
NAND2X1 NAND2X1_5 ( .A(w_cout_5_), .B(_34__3_), .Y(_382_) );
OAI21X1 OAI21X1_6 ( .A(w_cout_5_), .B(_381_), .C(_382_), .Y(_0__27_) );
INVX1 INVX1_6 ( .A(gnd), .Y(_386_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_387_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_388_) );
NAND3X1 NAND3X1_1 ( .A(_386_), .B(_388_), .C(_387_), .Y(_389_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_383_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_384_) );
OAI21X1 OAI21X1_7 ( .A(_383_), .B(_384_), .C(gnd), .Y(_385_) );
NAND2X1 NAND2X1_7 ( .A(_385_), .B(_389_), .Y(_33__0_) );
OAI21X1 OAI21X1_8 ( .A(_386_), .B(_383_), .C(_388_), .Y(_35__1_) );
INVX1 INVX1_7 ( .A(_35__3_), .Y(_393_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_394_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_395_) );
NAND3X1 NAND3X1_2 ( .A(_393_), .B(_395_), .C(_394_), .Y(_396_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_390_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_391_) );
OAI21X1 OAI21X1_9 ( .A(_390_), .B(_391_), .C(_35__3_), .Y(_392_) );
NAND2X1 NAND2X1_9 ( .A(_392_), .B(_396_), .Y(_33__3_) );
OAI21X1 OAI21X1_10 ( .A(_393_), .B(_390_), .C(_395_), .Y(_31_) );
INVX1 INVX1_8 ( .A(_35__1_), .Y(_400_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_401_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_402_) );
NAND3X1 NAND3X1_3 ( .A(_400_), .B(_402_), .C(_401_), .Y(_403_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_397_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_398_) );
OAI21X1 OAI21X1_11 ( .A(_397_), .B(_398_), .C(_35__1_), .Y(_399_) );
NAND2X1 NAND2X1_11 ( .A(_399_), .B(_403_), .Y(_33__1_) );
OAI21X1 OAI21X1_12 ( .A(_400_), .B(_397_), .C(_402_), .Y(_35__2_) );
INVX1 INVX1_9 ( .A(_35__2_), .Y(_407_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_408_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_409_) );
NAND3X1 NAND3X1_4 ( .A(_407_), .B(_409_), .C(_408_), .Y(_410_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_404_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_405_) );
OAI21X1 OAI21X1_13 ( .A(_404_), .B(_405_), .C(_35__2_), .Y(_406_) );
NAND2X1 NAND2X1_13 ( .A(_406_), .B(_410_), .Y(_33__2_) );
OAI21X1 OAI21X1_14 ( .A(_407_), .B(_404_), .C(_409_), .Y(_35__3_) );
INVX1 INVX1_10 ( .A(vdd), .Y(_414_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_415_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_416_) );
NAND3X1 NAND3X1_5 ( .A(_414_), .B(_416_), .C(_415_), .Y(_417_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_411_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_412_) );
OAI21X1 OAI21X1_15 ( .A(_411_), .B(_412_), .C(vdd), .Y(_413_) );
NAND2X1 NAND2X1_15 ( .A(_413_), .B(_417_), .Y(_34__0_) );
OAI21X1 OAI21X1_16 ( .A(_414_), .B(_411_), .C(_416_), .Y(_36__1_) );
INVX1 INVX1_11 ( .A(_36__3_), .Y(_421_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_422_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_423_) );
NAND3X1 NAND3X1_6 ( .A(_421_), .B(_423_), .C(_422_), .Y(_424_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_418_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_419_) );
OAI21X1 OAI21X1_17 ( .A(_418_), .B(_419_), .C(_36__3_), .Y(_420_) );
NAND2X1 NAND2X1_17 ( .A(_420_), .B(_424_), .Y(_34__3_) );
OAI21X1 OAI21X1_18 ( .A(_421_), .B(_418_), .C(_423_), .Y(_32_) );
INVX1 INVX1_12 ( .A(_36__1_), .Y(_428_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_429_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_430_) );
NAND3X1 NAND3X1_7 ( .A(_428_), .B(_430_), .C(_429_), .Y(_431_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_425_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_426_) );
OAI21X1 OAI21X1_19 ( .A(_425_), .B(_426_), .C(_36__1_), .Y(_427_) );
NAND2X1 NAND2X1_19 ( .A(_427_), .B(_431_), .Y(_34__1_) );
OAI21X1 OAI21X1_20 ( .A(_428_), .B(_425_), .C(_430_), .Y(_36__2_) );
INVX1 INVX1_13 ( .A(_36__2_), .Y(_435_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_436_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_437_) );
NAND3X1 NAND3X1_8 ( .A(_435_), .B(_437_), .C(_436_), .Y(_438_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_432_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_433_) );
OAI21X1 OAI21X1_21 ( .A(_432_), .B(_433_), .C(_36__2_), .Y(_434_) );
NAND2X1 NAND2X1_21 ( .A(_434_), .B(_438_), .Y(_34__2_) );
OAI21X1 OAI21X1_22 ( .A(_435_), .B(_432_), .C(_437_), .Y(_36__3_) );
INVX1 INVX1_14 ( .A(_37_), .Y(_439_) );
NAND2X1 NAND2X1_22 ( .A(_38_), .B(w_cout_6_), .Y(_440_) );
OAI21X1 OAI21X1_23 ( .A(w_cout_6_), .B(_439_), .C(_440_), .Y(w_cout_7_) );
INVX1 INVX1_15 ( .A(_39__0_), .Y(_441_) );
NAND2X1 NAND2X1_23 ( .A(_40__0_), .B(w_cout_6_), .Y(_442_) );
OAI21X1 OAI21X1_24 ( .A(w_cout_6_), .B(_441_), .C(_442_), .Y(_0__28_) );
INVX1 INVX1_16 ( .A(_39__1_), .Y(_443_) );
NAND2X1 NAND2X1_24 ( .A(w_cout_6_), .B(_40__1_), .Y(_444_) );
OAI21X1 OAI21X1_25 ( .A(w_cout_6_), .B(_443_), .C(_444_), .Y(_0__29_) );
INVX1 INVX1_17 ( .A(_39__2_), .Y(_445_) );
NAND2X1 NAND2X1_25 ( .A(w_cout_6_), .B(_40__2_), .Y(_446_) );
OAI21X1 OAI21X1_26 ( .A(w_cout_6_), .B(_445_), .C(_446_), .Y(_0__30_) );
INVX1 INVX1_18 ( .A(_39__3_), .Y(_447_) );
NAND2X1 NAND2X1_26 ( .A(w_cout_6_), .B(_40__3_), .Y(_448_) );
OAI21X1 OAI21X1_27 ( .A(w_cout_6_), .B(_447_), .C(_448_), .Y(_0__31_) );
INVX1 INVX1_19 ( .A(gnd), .Y(_452_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_453_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_454_) );
NAND3X1 NAND3X1_9 ( .A(_452_), .B(_454_), .C(_453_), .Y(_455_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_449_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_450_) );
OAI21X1 OAI21X1_28 ( .A(_449_), .B(_450_), .C(gnd), .Y(_451_) );
NAND2X1 NAND2X1_28 ( .A(_451_), .B(_455_), .Y(_39__0_) );
OAI21X1 OAI21X1_29 ( .A(_452_), .B(_449_), .C(_454_), .Y(_41__1_) );
INVX1 INVX1_20 ( .A(_41__3_), .Y(_459_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_460_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_461_) );
NAND3X1 NAND3X1_10 ( .A(_459_), .B(_461_), .C(_460_), .Y(_462_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_456_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_457_) );
OAI21X1 OAI21X1_30 ( .A(_456_), .B(_457_), .C(_41__3_), .Y(_458_) );
NAND2X1 NAND2X1_30 ( .A(_458_), .B(_462_), .Y(_39__3_) );
OAI21X1 OAI21X1_31 ( .A(_459_), .B(_456_), .C(_461_), .Y(_37_) );
INVX1 INVX1_21 ( .A(_41__1_), .Y(_466_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_467_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_468_) );
NAND3X1 NAND3X1_11 ( .A(_466_), .B(_468_), .C(_467_), .Y(_469_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_463_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_464_) );
OAI21X1 OAI21X1_32 ( .A(_463_), .B(_464_), .C(_41__1_), .Y(_465_) );
NAND2X1 NAND2X1_32 ( .A(_465_), .B(_469_), .Y(_39__1_) );
OAI21X1 OAI21X1_33 ( .A(_466_), .B(_463_), .C(_468_), .Y(_41__2_) );
INVX1 INVX1_22 ( .A(_41__2_), .Y(_473_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_474_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_475_) );
NAND3X1 NAND3X1_12 ( .A(_473_), .B(_475_), .C(_474_), .Y(_476_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_470_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_471_) );
OAI21X1 OAI21X1_34 ( .A(_470_), .B(_471_), .C(_41__2_), .Y(_472_) );
NAND2X1 NAND2X1_34 ( .A(_472_), .B(_476_), .Y(_39__2_) );
OAI21X1 OAI21X1_35 ( .A(_473_), .B(_470_), .C(_475_), .Y(_41__3_) );
INVX1 INVX1_23 ( .A(vdd), .Y(_480_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_481_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_482_) );
NAND3X1 NAND3X1_13 ( .A(_480_), .B(_482_), .C(_481_), .Y(_483_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_477_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_478_) );
OAI21X1 OAI21X1_36 ( .A(_477_), .B(_478_), .C(vdd), .Y(_479_) );
NAND2X1 NAND2X1_36 ( .A(_479_), .B(_483_), .Y(_40__0_) );
OAI21X1 OAI21X1_37 ( .A(_480_), .B(_477_), .C(_482_), .Y(_42__1_) );
INVX1 INVX1_24 ( .A(_42__3_), .Y(_487_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_488_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_489_) );
NAND3X1 NAND3X1_14 ( .A(_487_), .B(_489_), .C(_488_), .Y(_490_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_484_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_485_) );
OAI21X1 OAI21X1_38 ( .A(_484_), .B(_485_), .C(_42__3_), .Y(_486_) );
NAND2X1 NAND2X1_38 ( .A(_486_), .B(_490_), .Y(_40__3_) );
OAI21X1 OAI21X1_39 ( .A(_487_), .B(_484_), .C(_489_), .Y(_38_) );
INVX1 INVX1_25 ( .A(_42__1_), .Y(_494_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_495_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_496_) );
NAND3X1 NAND3X1_15 ( .A(_494_), .B(_496_), .C(_495_), .Y(_497_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_491_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_492_) );
OAI21X1 OAI21X1_40 ( .A(_491_), .B(_492_), .C(_42__1_), .Y(_493_) );
NAND2X1 NAND2X1_40 ( .A(_493_), .B(_497_), .Y(_40__1_) );
OAI21X1 OAI21X1_41 ( .A(_494_), .B(_491_), .C(_496_), .Y(_42__2_) );
INVX1 INVX1_26 ( .A(_42__2_), .Y(_501_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_502_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_503_) );
NAND3X1 NAND3X1_16 ( .A(_501_), .B(_503_), .C(_502_), .Y(_504_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_498_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_499_) );
OAI21X1 OAI21X1_42 ( .A(_498_), .B(_499_), .C(_42__2_), .Y(_500_) );
NAND2X1 NAND2X1_42 ( .A(_500_), .B(_504_), .Y(_40__2_) );
OAI21X1 OAI21X1_43 ( .A(_501_), .B(_498_), .C(_503_), .Y(_42__3_) );
INVX1 INVX1_27 ( .A(gnd), .Y(_508_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_509_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_510_) );
NAND3X1 NAND3X1_17 ( .A(_508_), .B(_510_), .C(_509_), .Y(_511_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_505_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_506_) );
OAI21X1 OAI21X1_44 ( .A(_505_), .B(_506_), .C(gnd), .Y(_507_) );
NAND2X1 NAND2X1_44 ( .A(_507_), .B(_511_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_45 ( .A(_508_), .B(_505_), .C(_510_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_28 ( .A(rca_inst_fa31_i_carry), .Y(_515_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_516_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_517_) );
NAND3X1 NAND3X1_18 ( .A(_515_), .B(_517_), .C(_516_), .Y(_518_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_512_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_513_) );
OAI21X1 OAI21X1_46 ( .A(_512_), .B(_513_), .C(rca_inst_fa31_i_carry), .Y(_514_) );
NAND2X1 NAND2X1_46 ( .A(_514_), .B(_518_), .Y(rca_inst_fa31_o_sum) );
OAI21X1 OAI21X1_47 ( .A(_515_), .B(_512_), .C(_517_), .Y(rca_inst_cout) );
INVX1 INVX1_29 ( .A(rca_inst_fa0_o_carry), .Y(_522_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_523_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_524_) );
NAND3X1 NAND3X1_19 ( .A(_522_), .B(_524_), .C(_523_), .Y(_525_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_519_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_520_) );
OAI21X1 OAI21X1_48 ( .A(_519_), .B(_520_), .C(rca_inst_fa0_o_carry), .Y(_521_) );
NAND2X1 NAND2X1_48 ( .A(_521_), .B(_525_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_49 ( .A(_522_), .B(_519_), .C(_524_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_30 ( .A(rca_inst_fa_1__o_carry), .Y(_529_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_530_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_531_) );
NAND3X1 NAND3X1_20 ( .A(_529_), .B(_531_), .C(_530_), .Y(_532_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_526_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_527_) );
OAI21X1 OAI21X1_50 ( .A(_526_), .B(_527_), .C(rca_inst_fa_1__o_carry), .Y(_528_) );
NAND2X1 NAND2X1_50 ( .A(_528_), .B(_532_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_51 ( .A(_529_), .B(_526_), .C(_531_), .Y(rca_inst_fa31_i_carry) );
BUFX2 BUFX2_1 ( .A(w_cout_7_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa31_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
INVX1 INVX1_31 ( .A(_1_), .Y(_43_) );
NAND2X1 NAND2X1_51 ( .A(_2_), .B(rca_inst_cout), .Y(_44_) );
OAI21X1 OAI21X1_52 ( .A(rca_inst_cout), .B(_43_), .C(_44_), .Y(w_cout_1_) );
INVX1 INVX1_32 ( .A(_3__0_), .Y(_45_) );
NAND2X1 NAND2X1_52 ( .A(_4__0_), .B(rca_inst_cout), .Y(_46_) );
OAI21X1 OAI21X1_53 ( .A(rca_inst_cout), .B(_45_), .C(_46_), .Y(_0__4_) );
INVX1 INVX1_33 ( .A(_3__1_), .Y(_47_) );
NAND2X1 NAND2X1_53 ( .A(rca_inst_cout), .B(_4__1_), .Y(_48_) );
OAI21X1 OAI21X1_54 ( .A(rca_inst_cout), .B(_47_), .C(_48_), .Y(_0__5_) );
INVX1 INVX1_34 ( .A(_3__2_), .Y(_49_) );
NAND2X1 NAND2X1_54 ( .A(rca_inst_cout), .B(_4__2_), .Y(_50_) );
OAI21X1 OAI21X1_55 ( .A(rca_inst_cout), .B(_49_), .C(_50_), .Y(_0__6_) );
INVX1 INVX1_35 ( .A(_3__3_), .Y(_51_) );
NAND2X1 NAND2X1_55 ( .A(rca_inst_cout), .B(_4__3_), .Y(_52_) );
OAI21X1 OAI21X1_56 ( .A(rca_inst_cout), .B(_51_), .C(_52_), .Y(_0__7_) );
INVX1 INVX1_36 ( .A(gnd), .Y(_56_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_57_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_58_) );
NAND3X1 NAND3X1_21 ( .A(_56_), .B(_58_), .C(_57_), .Y(_59_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_53_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_54_) );
OAI21X1 OAI21X1_57 ( .A(_53_), .B(_54_), .C(gnd), .Y(_55_) );
NAND2X1 NAND2X1_57 ( .A(_55_), .B(_59_), .Y(_3__0_) );
OAI21X1 OAI21X1_58 ( .A(_56_), .B(_53_), .C(_58_), .Y(_5__1_) );
INVX1 INVX1_37 ( .A(_5__3_), .Y(_63_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_64_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_65_) );
NAND3X1 NAND3X1_22 ( .A(_63_), .B(_65_), .C(_64_), .Y(_66_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_60_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_61_) );
OAI21X1 OAI21X1_59 ( .A(_60_), .B(_61_), .C(_5__3_), .Y(_62_) );
NAND2X1 NAND2X1_59 ( .A(_62_), .B(_66_), .Y(_3__3_) );
OAI21X1 OAI21X1_60 ( .A(_63_), .B(_60_), .C(_65_), .Y(_1_) );
INVX1 INVX1_38 ( .A(_5__1_), .Y(_70_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_71_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_72_) );
NAND3X1 NAND3X1_23 ( .A(_70_), .B(_72_), .C(_71_), .Y(_73_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_67_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_68_) );
OAI21X1 OAI21X1_61 ( .A(_67_), .B(_68_), .C(_5__1_), .Y(_69_) );
NAND2X1 NAND2X1_61 ( .A(_69_), .B(_73_), .Y(_3__1_) );
OAI21X1 OAI21X1_62 ( .A(_70_), .B(_67_), .C(_72_), .Y(_5__2_) );
INVX1 INVX1_39 ( .A(_5__2_), .Y(_77_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_78_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_79_) );
NAND3X1 NAND3X1_24 ( .A(_77_), .B(_79_), .C(_78_), .Y(_80_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_74_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_75_) );
OAI21X1 OAI21X1_63 ( .A(_74_), .B(_75_), .C(_5__2_), .Y(_76_) );
NAND2X1 NAND2X1_63 ( .A(_76_), .B(_80_), .Y(_3__2_) );
OAI21X1 OAI21X1_64 ( .A(_77_), .B(_74_), .C(_79_), .Y(_5__3_) );
INVX1 INVX1_40 ( .A(vdd), .Y(_84_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_85_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_86_) );
NAND3X1 NAND3X1_25 ( .A(_84_), .B(_86_), .C(_85_), .Y(_87_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_81_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_82_) );
OAI21X1 OAI21X1_65 ( .A(_81_), .B(_82_), .C(vdd), .Y(_83_) );
NAND2X1 NAND2X1_65 ( .A(_83_), .B(_87_), .Y(_4__0_) );
OAI21X1 OAI21X1_66 ( .A(_84_), .B(_81_), .C(_86_), .Y(_6__1_) );
INVX1 INVX1_41 ( .A(_6__3_), .Y(_91_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_92_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_93_) );
NAND3X1 NAND3X1_26 ( .A(_91_), .B(_93_), .C(_92_), .Y(_94_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_88_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_89_) );
OAI21X1 OAI21X1_67 ( .A(_88_), .B(_89_), .C(_6__3_), .Y(_90_) );
NAND2X1 NAND2X1_67 ( .A(_90_), .B(_94_), .Y(_4__3_) );
OAI21X1 OAI21X1_68 ( .A(_91_), .B(_88_), .C(_93_), .Y(_2_) );
INVX1 INVX1_42 ( .A(_6__1_), .Y(_98_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_99_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_100_) );
NAND3X1 NAND3X1_27 ( .A(_98_), .B(_100_), .C(_99_), .Y(_101_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_95_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_96_) );
OAI21X1 OAI21X1_69 ( .A(_95_), .B(_96_), .C(_6__1_), .Y(_97_) );
NAND2X1 NAND2X1_69 ( .A(_97_), .B(_101_), .Y(_4__1_) );
OAI21X1 OAI21X1_70 ( .A(_98_), .B(_95_), .C(_100_), .Y(_6__2_) );
INVX1 INVX1_43 ( .A(_6__2_), .Y(_105_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_106_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_107_) );
NAND3X1 NAND3X1_28 ( .A(_105_), .B(_107_), .C(_106_), .Y(_108_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_102_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_103_) );
OAI21X1 OAI21X1_71 ( .A(_102_), .B(_103_), .C(_6__2_), .Y(_104_) );
NAND2X1 NAND2X1_71 ( .A(_104_), .B(_108_), .Y(_4__2_) );
OAI21X1 OAI21X1_72 ( .A(_105_), .B(_102_), .C(_107_), .Y(_6__3_) );
INVX1 INVX1_44 ( .A(_7_), .Y(_109_) );
NAND2X1 NAND2X1_72 ( .A(_8_), .B(w_cout_1_), .Y(_110_) );
OAI21X1 OAI21X1_73 ( .A(w_cout_1_), .B(_109_), .C(_110_), .Y(w_cout_2_) );
INVX1 INVX1_45 ( .A(_9__0_), .Y(_111_) );
NAND2X1 NAND2X1_73 ( .A(_10__0_), .B(w_cout_1_), .Y(_112_) );
OAI21X1 OAI21X1_74 ( .A(w_cout_1_), .B(_111_), .C(_112_), .Y(_0__8_) );
INVX1 INVX1_46 ( .A(_9__1_), .Y(_113_) );
NAND2X1 NAND2X1_74 ( .A(w_cout_1_), .B(_10__1_), .Y(_114_) );
OAI21X1 OAI21X1_75 ( .A(w_cout_1_), .B(_113_), .C(_114_), .Y(_0__9_) );
INVX1 INVX1_47 ( .A(_9__2_), .Y(_115_) );
NAND2X1 NAND2X1_75 ( .A(w_cout_1_), .B(_10__2_), .Y(_116_) );
OAI21X1 OAI21X1_76 ( .A(w_cout_1_), .B(_115_), .C(_116_), .Y(_0__10_) );
INVX1 INVX1_48 ( .A(_9__3_), .Y(_117_) );
NAND2X1 NAND2X1_76 ( .A(w_cout_1_), .B(_10__3_), .Y(_118_) );
OAI21X1 OAI21X1_77 ( .A(w_cout_1_), .B(_117_), .C(_118_), .Y(_0__11_) );
INVX1 INVX1_49 ( .A(gnd), .Y(_122_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_123_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_124_) );
NAND3X1 NAND3X1_29 ( .A(_122_), .B(_124_), .C(_123_), .Y(_125_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_119_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_120_) );
OAI21X1 OAI21X1_78 ( .A(_119_), .B(_120_), .C(gnd), .Y(_121_) );
NAND2X1 NAND2X1_78 ( .A(_121_), .B(_125_), .Y(_9__0_) );
OAI21X1 OAI21X1_79 ( .A(_122_), .B(_119_), .C(_124_), .Y(_11__1_) );
INVX1 INVX1_50 ( .A(_11__3_), .Y(_129_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_130_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_131_) );
NAND3X1 NAND3X1_30 ( .A(_129_), .B(_131_), .C(_130_), .Y(_132_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_126_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_127_) );
OAI21X1 OAI21X1_80 ( .A(_126_), .B(_127_), .C(_11__3_), .Y(_128_) );
NAND2X1 NAND2X1_80 ( .A(_128_), .B(_132_), .Y(_9__3_) );
OAI21X1 OAI21X1_81 ( .A(_129_), .B(_126_), .C(_131_), .Y(_7_) );
INVX1 INVX1_51 ( .A(_11__1_), .Y(_136_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_137_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_138_) );
NAND3X1 NAND3X1_31 ( .A(_136_), .B(_138_), .C(_137_), .Y(_139_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_133_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_134_) );
OAI21X1 OAI21X1_82 ( .A(_133_), .B(_134_), .C(_11__1_), .Y(_135_) );
NAND2X1 NAND2X1_82 ( .A(_135_), .B(_139_), .Y(_9__1_) );
OAI21X1 OAI21X1_83 ( .A(_136_), .B(_133_), .C(_138_), .Y(_11__2_) );
INVX1 INVX1_52 ( .A(_11__2_), .Y(_143_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_144_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_145_) );
NAND3X1 NAND3X1_32 ( .A(_143_), .B(_145_), .C(_144_), .Y(_146_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_140_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_141_) );
OAI21X1 OAI21X1_84 ( .A(_140_), .B(_141_), .C(_11__2_), .Y(_142_) );
NAND2X1 NAND2X1_84 ( .A(_142_), .B(_146_), .Y(_9__2_) );
OAI21X1 OAI21X1_85 ( .A(_143_), .B(_140_), .C(_145_), .Y(_11__3_) );
INVX1 INVX1_53 ( .A(vdd), .Y(_150_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_151_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_152_) );
NAND3X1 NAND3X1_33 ( .A(_150_), .B(_152_), .C(_151_), .Y(_153_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_147_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_148_) );
OAI21X1 OAI21X1_86 ( .A(_147_), .B(_148_), .C(vdd), .Y(_149_) );
NAND2X1 NAND2X1_86 ( .A(_149_), .B(_153_), .Y(_10__0_) );
OAI21X1 OAI21X1_87 ( .A(_150_), .B(_147_), .C(_152_), .Y(_12__1_) );
INVX1 INVX1_54 ( .A(_12__3_), .Y(_157_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_158_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_159_) );
NAND3X1 NAND3X1_34 ( .A(_157_), .B(_159_), .C(_158_), .Y(_160_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_154_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_155_) );
OAI21X1 OAI21X1_88 ( .A(_154_), .B(_155_), .C(_12__3_), .Y(_156_) );
NAND2X1 NAND2X1_88 ( .A(_156_), .B(_160_), .Y(_10__3_) );
OAI21X1 OAI21X1_89 ( .A(_157_), .B(_154_), .C(_159_), .Y(_8_) );
INVX1 INVX1_55 ( .A(_12__1_), .Y(_164_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_165_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_166_) );
NAND3X1 NAND3X1_35 ( .A(_164_), .B(_166_), .C(_165_), .Y(_167_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_161_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_162_) );
OAI21X1 OAI21X1_90 ( .A(_161_), .B(_162_), .C(_12__1_), .Y(_163_) );
NAND2X1 NAND2X1_90 ( .A(_163_), .B(_167_), .Y(_10__1_) );
OAI21X1 OAI21X1_91 ( .A(_164_), .B(_161_), .C(_166_), .Y(_12__2_) );
INVX1 INVX1_56 ( .A(_12__2_), .Y(_171_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_172_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_173_) );
NAND3X1 NAND3X1_36 ( .A(_171_), .B(_173_), .C(_172_), .Y(_174_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_168_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_169_) );
OAI21X1 OAI21X1_92 ( .A(_168_), .B(_169_), .C(_12__2_), .Y(_170_) );
NAND2X1 NAND2X1_92 ( .A(_170_), .B(_174_), .Y(_10__2_) );
OAI21X1 OAI21X1_93 ( .A(_171_), .B(_168_), .C(_173_), .Y(_12__3_) );
INVX1 INVX1_57 ( .A(_13_), .Y(_175_) );
NAND2X1 NAND2X1_93 ( .A(_14_), .B(w_cout_2_), .Y(_176_) );
OAI21X1 OAI21X1_94 ( .A(w_cout_2_), .B(_175_), .C(_176_), .Y(w_cout_3_) );
INVX1 INVX1_58 ( .A(_15__0_), .Y(_177_) );
NAND2X1 NAND2X1_94 ( .A(_16__0_), .B(w_cout_2_), .Y(_178_) );
OAI21X1 OAI21X1_95 ( .A(w_cout_2_), .B(_177_), .C(_178_), .Y(_0__12_) );
INVX1 INVX1_59 ( .A(_15__1_), .Y(_179_) );
NAND2X1 NAND2X1_95 ( .A(w_cout_2_), .B(_16__1_), .Y(_180_) );
OAI21X1 OAI21X1_96 ( .A(w_cout_2_), .B(_179_), .C(_180_), .Y(_0__13_) );
INVX1 INVX1_60 ( .A(_15__2_), .Y(_181_) );
NAND2X1 NAND2X1_96 ( .A(w_cout_2_), .B(_16__2_), .Y(_182_) );
OAI21X1 OAI21X1_97 ( .A(w_cout_2_), .B(_181_), .C(_182_), .Y(_0__14_) );
INVX1 INVX1_61 ( .A(_15__3_), .Y(_183_) );
NAND2X1 NAND2X1_97 ( .A(w_cout_2_), .B(_16__3_), .Y(_184_) );
OAI21X1 OAI21X1_98 ( .A(w_cout_2_), .B(_183_), .C(_184_), .Y(_0__15_) );
INVX1 INVX1_62 ( .A(gnd), .Y(_188_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_189_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_190_) );
NAND3X1 NAND3X1_37 ( .A(_188_), .B(_190_), .C(_189_), .Y(_191_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_185_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_186_) );
OAI21X1 OAI21X1_99 ( .A(_185_), .B(_186_), .C(gnd), .Y(_187_) );
NAND2X1 NAND2X1_99 ( .A(_187_), .B(_191_), .Y(_15__0_) );
OAI21X1 OAI21X1_100 ( .A(_188_), .B(_185_), .C(_190_), .Y(_17__1_) );
INVX1 INVX1_63 ( .A(_17__3_), .Y(_195_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_196_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_197_) );
NAND3X1 NAND3X1_38 ( .A(_195_), .B(_197_), .C(_196_), .Y(_198_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_192_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_193_) );
OAI21X1 OAI21X1_101 ( .A(_192_), .B(_193_), .C(_17__3_), .Y(_194_) );
NAND2X1 NAND2X1_101 ( .A(_194_), .B(_198_), .Y(_15__3_) );
OAI21X1 OAI21X1_102 ( .A(_195_), .B(_192_), .C(_197_), .Y(_13_) );
INVX1 INVX1_64 ( .A(_17__1_), .Y(_202_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_203_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_204_) );
NAND3X1 NAND3X1_39 ( .A(_202_), .B(_204_), .C(_203_), .Y(_205_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_199_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_200_) );
OAI21X1 OAI21X1_103 ( .A(_199_), .B(_200_), .C(_17__1_), .Y(_201_) );
NAND2X1 NAND2X1_103 ( .A(_201_), .B(_205_), .Y(_15__1_) );
OAI21X1 OAI21X1_104 ( .A(_202_), .B(_199_), .C(_204_), .Y(_17__2_) );
INVX1 INVX1_65 ( .A(_17__2_), .Y(_209_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_210_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_211_) );
NAND3X1 NAND3X1_40 ( .A(_209_), .B(_211_), .C(_210_), .Y(_212_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_206_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_207_) );
OAI21X1 OAI21X1_105 ( .A(_206_), .B(_207_), .C(_17__2_), .Y(_208_) );
NAND2X1 NAND2X1_105 ( .A(_208_), .B(_212_), .Y(_15__2_) );
OAI21X1 OAI21X1_106 ( .A(_209_), .B(_206_), .C(_211_), .Y(_17__3_) );
INVX1 INVX1_66 ( .A(vdd), .Y(_216_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_217_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_218_) );
NAND3X1 NAND3X1_41 ( .A(_216_), .B(_218_), .C(_217_), .Y(_219_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_213_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_214_) );
OAI21X1 OAI21X1_107 ( .A(_213_), .B(_214_), .C(vdd), .Y(_215_) );
NAND2X1 NAND2X1_107 ( .A(_215_), .B(_219_), .Y(_16__0_) );
OAI21X1 OAI21X1_108 ( .A(_216_), .B(_213_), .C(_218_), .Y(_18__1_) );
INVX1 INVX1_67 ( .A(_18__3_), .Y(_223_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_224_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_225_) );
NAND3X1 NAND3X1_42 ( .A(_223_), .B(_225_), .C(_224_), .Y(_226_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_220_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_221_) );
OAI21X1 OAI21X1_109 ( .A(_220_), .B(_221_), .C(_18__3_), .Y(_222_) );
NAND2X1 NAND2X1_109 ( .A(_222_), .B(_226_), .Y(_16__3_) );
OAI21X1 OAI21X1_110 ( .A(_223_), .B(_220_), .C(_225_), .Y(_14_) );
INVX1 INVX1_68 ( .A(_18__1_), .Y(_230_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_231_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_232_) );
NAND3X1 NAND3X1_43 ( .A(_230_), .B(_232_), .C(_231_), .Y(_233_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_227_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_228_) );
OAI21X1 OAI21X1_111 ( .A(_227_), .B(_228_), .C(_18__1_), .Y(_229_) );
NAND2X1 NAND2X1_111 ( .A(_229_), .B(_233_), .Y(_16__1_) );
OAI21X1 OAI21X1_112 ( .A(_230_), .B(_227_), .C(_232_), .Y(_18__2_) );
INVX1 INVX1_69 ( .A(_18__2_), .Y(_237_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_238_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_239_) );
NAND3X1 NAND3X1_44 ( .A(_237_), .B(_239_), .C(_238_), .Y(_240_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_234_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_235_) );
OAI21X1 OAI21X1_113 ( .A(_234_), .B(_235_), .C(_18__2_), .Y(_236_) );
NAND2X1 NAND2X1_113 ( .A(_236_), .B(_240_), .Y(_16__2_) );
OAI21X1 OAI21X1_114 ( .A(_237_), .B(_234_), .C(_239_), .Y(_18__3_) );
INVX1 INVX1_70 ( .A(_19_), .Y(_241_) );
NAND2X1 NAND2X1_114 ( .A(_20_), .B(w_cout_3_), .Y(_242_) );
OAI21X1 OAI21X1_115 ( .A(w_cout_3_), .B(_241_), .C(_242_), .Y(w_cout_4_) );
INVX1 INVX1_71 ( .A(_21__0_), .Y(_243_) );
NAND2X1 NAND2X1_115 ( .A(_22__0_), .B(w_cout_3_), .Y(_244_) );
OAI21X1 OAI21X1_116 ( .A(w_cout_3_), .B(_243_), .C(_244_), .Y(_0__16_) );
INVX1 INVX1_72 ( .A(_21__1_), .Y(_245_) );
NAND2X1 NAND2X1_116 ( .A(w_cout_3_), .B(_22__1_), .Y(_246_) );
OAI21X1 OAI21X1_117 ( .A(w_cout_3_), .B(_245_), .C(_246_), .Y(_0__17_) );
INVX1 INVX1_73 ( .A(_21__2_), .Y(_247_) );
NAND2X1 NAND2X1_117 ( .A(w_cout_3_), .B(_22__2_), .Y(_248_) );
OAI21X1 OAI21X1_118 ( .A(w_cout_3_), .B(_247_), .C(_248_), .Y(_0__18_) );
INVX1 INVX1_74 ( .A(_21__3_), .Y(_249_) );
NAND2X1 NAND2X1_118 ( .A(w_cout_3_), .B(_22__3_), .Y(_250_) );
OAI21X1 OAI21X1_119 ( .A(w_cout_3_), .B(_249_), .C(_250_), .Y(_0__19_) );
INVX1 INVX1_75 ( .A(gnd), .Y(_254_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_255_) );
NAND2X1 NAND2X1_119 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_256_) );
NAND3X1 NAND3X1_45 ( .A(_254_), .B(_256_), .C(_255_), .Y(_257_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_251_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_252_) );
OAI21X1 OAI21X1_120 ( .A(_251_), .B(_252_), .C(gnd), .Y(_253_) );
NAND2X1 NAND2X1_120 ( .A(_253_), .B(_257_), .Y(_21__0_) );
OAI21X1 OAI21X1_121 ( .A(_254_), .B(_251_), .C(_256_), .Y(_23__1_) );
INVX1 INVX1_76 ( .A(_23__3_), .Y(_261_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_262_) );
NAND2X1 NAND2X1_121 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_263_) );
NAND3X1 NAND3X1_46 ( .A(_261_), .B(_263_), .C(_262_), .Y(_264_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_258_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_259_) );
OAI21X1 OAI21X1_122 ( .A(_258_), .B(_259_), .C(_23__3_), .Y(_260_) );
NAND2X1 NAND2X1_122 ( .A(_260_), .B(_264_), .Y(_21__3_) );
OAI21X1 OAI21X1_123 ( .A(_261_), .B(_258_), .C(_263_), .Y(_19_) );
INVX1 INVX1_77 ( .A(_23__1_), .Y(_268_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_269_) );
NAND2X1 NAND2X1_123 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_270_) );
NAND3X1 NAND3X1_47 ( .A(_268_), .B(_270_), .C(_269_), .Y(_271_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_265_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_266_) );
OAI21X1 OAI21X1_124 ( .A(_265_), .B(_266_), .C(_23__1_), .Y(_267_) );
NAND2X1 NAND2X1_124 ( .A(_267_), .B(_271_), .Y(_21__1_) );
OAI21X1 OAI21X1_125 ( .A(_268_), .B(_265_), .C(_270_), .Y(_23__2_) );
INVX1 INVX1_78 ( .A(_23__2_), .Y(_275_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_276_) );
NAND2X1 NAND2X1_125 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_277_) );
NAND3X1 NAND3X1_48 ( .A(_275_), .B(_277_), .C(_276_), .Y(_278_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_272_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_273_) );
OAI21X1 OAI21X1_126 ( .A(_272_), .B(_273_), .C(_23__2_), .Y(_274_) );
NAND2X1 NAND2X1_126 ( .A(_274_), .B(_278_), .Y(_21__2_) );
OAI21X1 OAI21X1_127 ( .A(_275_), .B(_272_), .C(_277_), .Y(_23__3_) );
INVX1 INVX1_79 ( .A(vdd), .Y(_282_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_283_) );
NAND2X1 NAND2X1_127 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_284_) );
NAND3X1 NAND3X1_49 ( .A(_282_), .B(_284_), .C(_283_), .Y(_285_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_279_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_280_) );
OAI21X1 OAI21X1_128 ( .A(_279_), .B(_280_), .C(vdd), .Y(_281_) );
NAND2X1 NAND2X1_128 ( .A(_281_), .B(_285_), .Y(_22__0_) );
OAI21X1 OAI21X1_129 ( .A(_282_), .B(_279_), .C(_284_), .Y(_24__1_) );
INVX1 INVX1_80 ( .A(_24__3_), .Y(_289_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_290_) );
NAND2X1 NAND2X1_129 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_291_) );
NAND3X1 NAND3X1_50 ( .A(_289_), .B(_291_), .C(_290_), .Y(_292_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_286_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_287_) );
OAI21X1 OAI21X1_130 ( .A(_286_), .B(_287_), .C(_24__3_), .Y(_288_) );
NAND2X1 NAND2X1_130 ( .A(_288_), .B(_292_), .Y(_22__3_) );
OAI21X1 OAI21X1_131 ( .A(_289_), .B(_286_), .C(_291_), .Y(_20_) );
INVX1 INVX1_81 ( .A(_24__1_), .Y(_296_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_297_) );
NAND2X1 NAND2X1_131 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_298_) );
NAND3X1 NAND3X1_51 ( .A(_296_), .B(_298_), .C(_297_), .Y(_299_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_293_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_294_) );
OAI21X1 OAI21X1_132 ( .A(_293_), .B(_294_), .C(_24__1_), .Y(_295_) );
NAND2X1 NAND2X1_132 ( .A(_295_), .B(_299_), .Y(_22__1_) );
OAI21X1 OAI21X1_133 ( .A(_296_), .B(_293_), .C(_298_), .Y(_24__2_) );
INVX1 INVX1_82 ( .A(_24__2_), .Y(_303_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_304_) );
NAND2X1 NAND2X1_133 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_305_) );
NAND3X1 NAND3X1_52 ( .A(_303_), .B(_305_), .C(_304_), .Y(_306_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_300_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_301_) );
OAI21X1 OAI21X1_134 ( .A(_300_), .B(_301_), .C(_24__2_), .Y(_302_) );
NAND2X1 NAND2X1_134 ( .A(_302_), .B(_306_), .Y(_22__2_) );
OAI21X1 OAI21X1_135 ( .A(_303_), .B(_300_), .C(_305_), .Y(_24__3_) );
INVX1 INVX1_83 ( .A(_25_), .Y(_307_) );
NAND2X1 NAND2X1_135 ( .A(_26_), .B(w_cout_4_), .Y(_308_) );
OAI21X1 OAI21X1_136 ( .A(w_cout_4_), .B(_307_), .C(_308_), .Y(w_cout_5_) );
INVX1 INVX1_84 ( .A(_27__0_), .Y(_309_) );
NAND2X1 NAND2X1_136 ( .A(_28__0_), .B(w_cout_4_), .Y(_310_) );
OAI21X1 OAI21X1_137 ( .A(w_cout_4_), .B(_309_), .C(_310_), .Y(_0__20_) );
INVX1 INVX1_85 ( .A(_27__1_), .Y(_311_) );
NAND2X1 NAND2X1_137 ( .A(w_cout_4_), .B(_28__1_), .Y(_312_) );
OAI21X1 OAI21X1_138 ( .A(w_cout_4_), .B(_311_), .C(_312_), .Y(_0__21_) );
INVX1 INVX1_86 ( .A(_27__2_), .Y(_313_) );
NAND2X1 NAND2X1_138 ( .A(w_cout_4_), .B(_28__2_), .Y(_314_) );
OAI21X1 OAI21X1_139 ( .A(w_cout_4_), .B(_313_), .C(_314_), .Y(_0__22_) );
INVX1 INVX1_87 ( .A(_27__3_), .Y(_315_) );
NAND2X1 NAND2X1_139 ( .A(w_cout_4_), .B(_28__3_), .Y(_316_) );
OAI21X1 OAI21X1_140 ( .A(w_cout_4_), .B(_315_), .C(_316_), .Y(_0__23_) );
INVX1 INVX1_88 ( .A(gnd), .Y(_320_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_321_) );
NAND2X1 NAND2X1_140 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_322_) );
NAND3X1 NAND3X1_53 ( .A(_320_), .B(_322_), .C(_321_), .Y(_323_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_317_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_318_) );
OAI21X1 OAI21X1_141 ( .A(_317_), .B(_318_), .C(gnd), .Y(_319_) );
NAND2X1 NAND2X1_141 ( .A(_319_), .B(_323_), .Y(_27__0_) );
OAI21X1 OAI21X1_142 ( .A(_320_), .B(_317_), .C(_322_), .Y(_29__1_) );
INVX1 INVX1_89 ( .A(_29__3_), .Y(_327_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_328_) );
NAND2X1 NAND2X1_142 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_329_) );
NAND3X1 NAND3X1_54 ( .A(_327_), .B(_329_), .C(_328_), .Y(_330_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_324_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_325_) );
OAI21X1 OAI21X1_143 ( .A(_324_), .B(_325_), .C(_29__3_), .Y(_326_) );
NAND2X1 NAND2X1_143 ( .A(_326_), .B(_330_), .Y(_27__3_) );
OAI21X1 OAI21X1_144 ( .A(_327_), .B(_324_), .C(_329_), .Y(_25_) );
INVX1 INVX1_90 ( .A(_29__1_), .Y(_334_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_335_) );
NAND2X1 NAND2X1_144 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_336_) );
NAND3X1 NAND3X1_55 ( .A(_334_), .B(_336_), .C(_335_), .Y(_337_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_331_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_332_) );
OAI21X1 OAI21X1_145 ( .A(_331_), .B(_332_), .C(_29__1_), .Y(_333_) );
NAND2X1 NAND2X1_145 ( .A(_333_), .B(_337_), .Y(_27__1_) );
OAI21X1 OAI21X1_146 ( .A(_334_), .B(_331_), .C(_336_), .Y(_29__2_) );
INVX1 INVX1_91 ( .A(_29__2_), .Y(_341_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_342_) );
NAND2X1 NAND2X1_146 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_343_) );
NAND3X1 NAND3X1_56 ( .A(_341_), .B(_343_), .C(_342_), .Y(_344_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_338_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_339_) );
OAI21X1 OAI21X1_147 ( .A(_338_), .B(_339_), .C(_29__2_), .Y(_340_) );
NAND2X1 NAND2X1_147 ( .A(_340_), .B(_344_), .Y(_27__2_) );
OAI21X1 OAI21X1_148 ( .A(_341_), .B(_338_), .C(_343_), .Y(_29__3_) );
INVX1 INVX1_92 ( .A(vdd), .Y(_348_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_349_) );
NAND2X1 NAND2X1_148 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_350_) );
NAND3X1 NAND3X1_57 ( .A(_348_), .B(_350_), .C(_349_), .Y(_351_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_345_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_346_) );
OAI21X1 OAI21X1_149 ( .A(_345_), .B(_346_), .C(vdd), .Y(_347_) );
NAND2X1 NAND2X1_149 ( .A(_347_), .B(_351_), .Y(_28__0_) );
OAI21X1 OAI21X1_150 ( .A(_348_), .B(_345_), .C(_350_), .Y(_30__1_) );
INVX1 INVX1_93 ( .A(_30__3_), .Y(_355_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_356_) );
NAND2X1 NAND2X1_150 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_357_) );
NAND3X1 NAND3X1_58 ( .A(_355_), .B(_357_), .C(_356_), .Y(_358_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_352_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_353_) );
OAI21X1 OAI21X1_151 ( .A(_352_), .B(_353_), .C(_30__3_), .Y(_354_) );
NAND2X1 NAND2X1_151 ( .A(_354_), .B(_358_), .Y(_28__3_) );
OAI21X1 OAI21X1_152 ( .A(_355_), .B(_352_), .C(_357_), .Y(_26_) );
INVX1 INVX1_94 ( .A(_30__1_), .Y(_362_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_363_) );
NAND2X1 NAND2X1_152 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_364_) );
NAND3X1 NAND3X1_59 ( .A(_362_), .B(_364_), .C(_363_), .Y(_365_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_359_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_360_) );
OAI21X1 OAI21X1_153 ( .A(_359_), .B(_360_), .C(_30__1_), .Y(_361_) );
NAND2X1 NAND2X1_153 ( .A(_361_), .B(_365_), .Y(_28__1_) );
OAI21X1 OAI21X1_154 ( .A(_362_), .B(_359_), .C(_364_), .Y(_30__2_) );
INVX1 INVX1_95 ( .A(_30__2_), .Y(_369_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_370_) );
NAND2X1 NAND2X1_154 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_371_) );
NAND3X1 NAND3X1_60 ( .A(_369_), .B(_371_), .C(_370_), .Y(_372_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_366_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_367_) );
OAI21X1 OAI21X1_155 ( .A(_366_), .B(_367_), .C(_30__2_), .Y(_368_) );
NAND2X1 NAND2X1_155 ( .A(_368_), .B(_372_), .Y(_28__2_) );
BUFX2 BUFX2_34 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_35 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_36 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_37 ( .A(rca_inst_fa31_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_38 ( .A(rca_inst_cout), .Y(w_cout_0_) );
endmodule
