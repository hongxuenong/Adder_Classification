module cla_50bit (i_add1, i_add2, o_result);

input [49:0] i_add1;
input [49:0] i_add2;
output [50:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX2 BUFX2_1 ( .A(_286__27_), .Y(o_result[27]) );
BUFX2 BUFX2_2 ( .A(_286__28_), .Y(o_result[28]) );
BUFX2 BUFX2_3 ( .A(_286__29_), .Y(o_result[29]) );
BUFX2 BUFX2_4 ( .A(_286__30_), .Y(o_result[30]) );
BUFX2 BUFX2_5 ( .A(_286__31_), .Y(o_result[31]) );
BUFX2 BUFX2_6 ( .A(_286__32_), .Y(o_result[32]) );
BUFX2 BUFX2_7 ( .A(_286__33_), .Y(o_result[33]) );
BUFX2 BUFX2_8 ( .A(_286__34_), .Y(o_result[34]) );
BUFX2 BUFX2_9 ( .A(_286__35_), .Y(o_result[35]) );
BUFX2 BUFX2_10 ( .A(_286__36_), .Y(o_result[36]) );
BUFX2 BUFX2_11 ( .A(_286__37_), .Y(o_result[37]) );
BUFX2 BUFX2_12 ( .A(_286__38_), .Y(o_result[38]) );
BUFX2 BUFX2_13 ( .A(_286__39_), .Y(o_result[39]) );
BUFX2 BUFX2_14 ( .A(_286__40_), .Y(o_result[40]) );
BUFX2 BUFX2_15 ( .A(_286__41_), .Y(o_result[41]) );
BUFX2 BUFX2_16 ( .A(_286__42_), .Y(o_result[42]) );
BUFX2 BUFX2_17 ( .A(_286__43_), .Y(o_result[43]) );
BUFX2 BUFX2_18 ( .A(_286__44_), .Y(o_result[44]) );
BUFX2 BUFX2_19 ( .A(_286__45_), .Y(o_result[45]) );
BUFX2 BUFX2_20 ( .A(_286__46_), .Y(o_result[46]) );
BUFX2 BUFX2_21 ( .A(_286__47_), .Y(o_result[47]) );
BUFX2 BUFX2_22 ( .A(_286__48_), .Y(o_result[48]) );
BUFX2 BUFX2_23 ( .A(_286__49_), .Y(o_result[49]) );
BUFX2 BUFX2_24 ( .A(w_C_50_), .Y(o_result[50]) );
INVX1 INVX1_1 ( .A(w_C_4_), .Y(_290_) );
OR2X2 OR2X2_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_291_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_292_) );
NAND3X1 NAND3X1_1 ( .A(_290_), .B(_292_), .C(_291_), .Y(_293_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_287_) );
AND2X2 AND2X2_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_288_) );
OAI21X1 OAI21X1_1 ( .A(_287_), .B(_288_), .C(w_C_4_), .Y(_289_) );
NAND2X1 NAND2X1_2 ( .A(_289_), .B(_293_), .Y(_286__4_) );
INVX1 INVX1_2 ( .A(w_C_5_), .Y(_297_) );
OR2X2 OR2X2_2 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_298_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_299_) );
NAND3X1 NAND3X1_2 ( .A(_297_), .B(_299_), .C(_298_), .Y(_300_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_294_) );
AND2X2 AND2X2_2 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_295_) );
OAI21X1 OAI21X1_2 ( .A(_294_), .B(_295_), .C(w_C_5_), .Y(_296_) );
NAND2X1 NAND2X1_4 ( .A(_296_), .B(_300_), .Y(_286__5_) );
INVX1 INVX1_3 ( .A(w_C_6_), .Y(_304_) );
OR2X2 OR2X2_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_305_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_306_) );
NAND3X1 NAND3X1_3 ( .A(_304_), .B(_306_), .C(_305_), .Y(_307_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_301_) );
AND2X2 AND2X2_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_302_) );
OAI21X1 OAI21X1_3 ( .A(_301_), .B(_302_), .C(w_C_6_), .Y(_303_) );
NAND2X1 NAND2X1_6 ( .A(_303_), .B(_307_), .Y(_286__6_) );
INVX1 INVX1_4 ( .A(w_C_7_), .Y(_311_) );
OR2X2 OR2X2_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_312_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_313_) );
NAND3X1 NAND3X1_4 ( .A(_311_), .B(_313_), .C(_312_), .Y(_314_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_308_) );
AND2X2 AND2X2_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_309_) );
OAI21X1 OAI21X1_4 ( .A(_308_), .B(_309_), .C(w_C_7_), .Y(_310_) );
NAND2X1 NAND2X1_8 ( .A(_310_), .B(_314_), .Y(_286__7_) );
INVX1 INVX1_5 ( .A(w_C_8_), .Y(_318_) );
OR2X2 OR2X2_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_319_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_320_) );
NAND3X1 NAND3X1_5 ( .A(_318_), .B(_320_), .C(_319_), .Y(_321_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_315_) );
AND2X2 AND2X2_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_316_) );
OAI21X1 OAI21X1_5 ( .A(_315_), .B(_316_), .C(w_C_8_), .Y(_317_) );
NAND2X1 NAND2X1_10 ( .A(_317_), .B(_321_), .Y(_286__8_) );
INVX1 INVX1_6 ( .A(w_C_9_), .Y(_325_) );
OR2X2 OR2X2_6 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_326_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_327_) );
NAND3X1 NAND3X1_6 ( .A(_325_), .B(_327_), .C(_326_), .Y(_328_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_322_) );
AND2X2 AND2X2_6 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_323_) );
OAI21X1 OAI21X1_6 ( .A(_322_), .B(_323_), .C(w_C_9_), .Y(_324_) );
NAND2X1 NAND2X1_12 ( .A(_324_), .B(_328_), .Y(_286__9_) );
INVX1 INVX1_7 ( .A(w_C_10_), .Y(_332_) );
OR2X2 OR2X2_7 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_333_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_334_) );
NAND3X1 NAND3X1_7 ( .A(_332_), .B(_334_), .C(_333_), .Y(_335_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_329_) );
AND2X2 AND2X2_7 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_330_) );
OAI21X1 OAI21X1_7 ( .A(_329_), .B(_330_), .C(w_C_10_), .Y(_331_) );
NAND2X1 NAND2X1_14 ( .A(_331_), .B(_335_), .Y(_286__10_) );
INVX1 INVX1_8 ( .A(w_C_11_), .Y(_339_) );
OR2X2 OR2X2_8 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_340_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_341_) );
NAND3X1 NAND3X1_8 ( .A(_339_), .B(_341_), .C(_340_), .Y(_342_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_336_) );
AND2X2 AND2X2_8 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_337_) );
OAI21X1 OAI21X1_8 ( .A(_336_), .B(_337_), .C(w_C_11_), .Y(_338_) );
NAND2X1 NAND2X1_16 ( .A(_338_), .B(_342_), .Y(_286__11_) );
INVX1 INVX1_9 ( .A(w_C_12_), .Y(_346_) );
OR2X2 OR2X2_9 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_347_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_348_) );
NAND3X1 NAND3X1_9 ( .A(_346_), .B(_348_), .C(_347_), .Y(_349_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_343_) );
AND2X2 AND2X2_9 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_344_) );
OAI21X1 OAI21X1_9 ( .A(_343_), .B(_344_), .C(w_C_12_), .Y(_345_) );
NAND2X1 NAND2X1_18 ( .A(_345_), .B(_349_), .Y(_286__12_) );
INVX1 INVX1_10 ( .A(w_C_13_), .Y(_353_) );
OR2X2 OR2X2_10 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_354_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_355_) );
NAND3X1 NAND3X1_10 ( .A(_353_), .B(_355_), .C(_354_), .Y(_356_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_350_) );
AND2X2 AND2X2_10 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_351_) );
OAI21X1 OAI21X1_10 ( .A(_350_), .B(_351_), .C(w_C_13_), .Y(_352_) );
NAND2X1 NAND2X1_20 ( .A(_352_), .B(_356_), .Y(_286__13_) );
INVX1 INVX1_11 ( .A(w_C_14_), .Y(_360_) );
OR2X2 OR2X2_11 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_361_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_362_) );
NAND3X1 NAND3X1_11 ( .A(_360_), .B(_362_), .C(_361_), .Y(_363_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_357_) );
AND2X2 AND2X2_11 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_358_) );
OAI21X1 OAI21X1_11 ( .A(_357_), .B(_358_), .C(w_C_14_), .Y(_359_) );
NAND2X1 NAND2X1_22 ( .A(_359_), .B(_363_), .Y(_286__14_) );
INVX1 INVX1_12 ( .A(w_C_15_), .Y(_367_) );
OR2X2 OR2X2_12 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_368_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_369_) );
NAND3X1 NAND3X1_12 ( .A(_367_), .B(_369_), .C(_368_), .Y(_370_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_364_) );
AND2X2 AND2X2_12 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_365_) );
OAI21X1 OAI21X1_12 ( .A(_364_), .B(_365_), .C(w_C_15_), .Y(_366_) );
NAND2X1 NAND2X1_24 ( .A(_366_), .B(_370_), .Y(_286__15_) );
INVX1 INVX1_13 ( .A(w_C_16_), .Y(_374_) );
OR2X2 OR2X2_13 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_375_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_376_) );
NAND3X1 NAND3X1_13 ( .A(_374_), .B(_376_), .C(_375_), .Y(_377_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_371_) );
AND2X2 AND2X2_13 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_372_) );
OAI21X1 OAI21X1_13 ( .A(_371_), .B(_372_), .C(w_C_16_), .Y(_373_) );
NAND2X1 NAND2X1_26 ( .A(_373_), .B(_377_), .Y(_286__16_) );
INVX1 INVX1_14 ( .A(w_C_17_), .Y(_381_) );
OR2X2 OR2X2_14 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_382_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_383_) );
NAND3X1 NAND3X1_14 ( .A(_381_), .B(_383_), .C(_382_), .Y(_384_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_378_) );
AND2X2 AND2X2_14 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_379_) );
OAI21X1 OAI21X1_14 ( .A(_378_), .B(_379_), .C(w_C_17_), .Y(_380_) );
NAND2X1 NAND2X1_28 ( .A(_380_), .B(_384_), .Y(_286__17_) );
INVX1 INVX1_15 ( .A(w_C_18_), .Y(_388_) );
OR2X2 OR2X2_15 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_389_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_390_) );
NAND3X1 NAND3X1_15 ( .A(_388_), .B(_390_), .C(_389_), .Y(_391_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_385_) );
AND2X2 AND2X2_15 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_386_) );
OAI21X1 OAI21X1_15 ( .A(_385_), .B(_386_), .C(w_C_18_), .Y(_387_) );
NAND2X1 NAND2X1_30 ( .A(_387_), .B(_391_), .Y(_286__18_) );
INVX1 INVX1_16 ( .A(w_C_19_), .Y(_395_) );
OR2X2 OR2X2_16 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_396_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_397_) );
NAND3X1 NAND3X1_16 ( .A(_395_), .B(_397_), .C(_396_), .Y(_398_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_392_) );
AND2X2 AND2X2_16 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_393_) );
OAI21X1 OAI21X1_16 ( .A(_392_), .B(_393_), .C(w_C_19_), .Y(_394_) );
NAND2X1 NAND2X1_32 ( .A(_394_), .B(_398_), .Y(_286__19_) );
INVX1 INVX1_17 ( .A(w_C_20_), .Y(_402_) );
OR2X2 OR2X2_17 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_403_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_404_) );
NAND3X1 NAND3X1_17 ( .A(_402_), .B(_404_), .C(_403_), .Y(_405_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_399_) );
AND2X2 AND2X2_17 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_400_) );
OAI21X1 OAI21X1_17 ( .A(_399_), .B(_400_), .C(w_C_20_), .Y(_401_) );
NAND2X1 NAND2X1_34 ( .A(_401_), .B(_405_), .Y(_286__20_) );
INVX1 INVX1_18 ( .A(w_C_21_), .Y(_409_) );
OR2X2 OR2X2_18 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_410_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_411_) );
NAND3X1 NAND3X1_18 ( .A(_409_), .B(_411_), .C(_410_), .Y(_412_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_406_) );
AND2X2 AND2X2_18 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_407_) );
OAI21X1 OAI21X1_18 ( .A(_406_), .B(_407_), .C(w_C_21_), .Y(_408_) );
NAND2X1 NAND2X1_36 ( .A(_408_), .B(_412_), .Y(_286__21_) );
INVX1 INVX1_19 ( .A(w_C_22_), .Y(_416_) );
OR2X2 OR2X2_19 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_417_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_418_) );
NAND3X1 NAND3X1_19 ( .A(_416_), .B(_418_), .C(_417_), .Y(_419_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_413_) );
AND2X2 AND2X2_19 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_414_) );
OAI21X1 OAI21X1_19 ( .A(_413_), .B(_414_), .C(w_C_22_), .Y(_415_) );
NAND2X1 NAND2X1_38 ( .A(_415_), .B(_419_), .Y(_286__22_) );
INVX1 INVX1_20 ( .A(w_C_23_), .Y(_423_) );
OR2X2 OR2X2_20 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_424_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_425_) );
NAND3X1 NAND3X1_20 ( .A(_423_), .B(_425_), .C(_424_), .Y(_426_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_420_) );
AND2X2 AND2X2_20 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_421_) );
OAI21X1 OAI21X1_20 ( .A(_420_), .B(_421_), .C(w_C_23_), .Y(_422_) );
NAND2X1 NAND2X1_40 ( .A(_422_), .B(_426_), .Y(_286__23_) );
INVX1 INVX1_21 ( .A(w_C_24_), .Y(_430_) );
OR2X2 OR2X2_21 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_431_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_432_) );
NAND3X1 NAND3X1_21 ( .A(_430_), .B(_432_), .C(_431_), .Y(_433_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_427_) );
AND2X2 AND2X2_21 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_428_) );
OAI21X1 OAI21X1_21 ( .A(_427_), .B(_428_), .C(w_C_24_), .Y(_429_) );
NAND2X1 NAND2X1_42 ( .A(_429_), .B(_433_), .Y(_286__24_) );
INVX1 INVX1_22 ( .A(w_C_25_), .Y(_437_) );
OR2X2 OR2X2_22 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_438_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_439_) );
NAND3X1 NAND3X1_22 ( .A(_437_), .B(_439_), .C(_438_), .Y(_440_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_434_) );
AND2X2 AND2X2_22 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_435_) );
OAI21X1 OAI21X1_22 ( .A(_434_), .B(_435_), .C(w_C_25_), .Y(_436_) );
NAND2X1 NAND2X1_44 ( .A(_436_), .B(_440_), .Y(_286__25_) );
INVX1 INVX1_23 ( .A(w_C_26_), .Y(_444_) );
OR2X2 OR2X2_23 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_445_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_446_) );
NAND3X1 NAND3X1_23 ( .A(_444_), .B(_446_), .C(_445_), .Y(_447_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_441_) );
AND2X2 AND2X2_23 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_442_) );
OAI21X1 OAI21X1_23 ( .A(_441_), .B(_442_), .C(w_C_26_), .Y(_443_) );
NAND2X1 NAND2X1_46 ( .A(_443_), .B(_447_), .Y(_286__26_) );
INVX1 INVX1_24 ( .A(w_C_27_), .Y(_451_) );
OR2X2 OR2X2_24 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_452_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_453_) );
NAND3X1 NAND3X1_24 ( .A(_451_), .B(_453_), .C(_452_), .Y(_454_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_448_) );
AND2X2 AND2X2_24 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_449_) );
OAI21X1 OAI21X1_24 ( .A(_448_), .B(_449_), .C(w_C_27_), .Y(_450_) );
NAND2X1 NAND2X1_48 ( .A(_450_), .B(_454_), .Y(_286__27_) );
INVX1 INVX1_25 ( .A(w_C_28_), .Y(_458_) );
OR2X2 OR2X2_25 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_459_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_460_) );
NAND3X1 NAND3X1_25 ( .A(_458_), .B(_460_), .C(_459_), .Y(_461_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_455_) );
AND2X2 AND2X2_25 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_456_) );
OAI21X1 OAI21X1_25 ( .A(_455_), .B(_456_), .C(w_C_28_), .Y(_457_) );
NAND2X1 NAND2X1_50 ( .A(_457_), .B(_461_), .Y(_286__28_) );
INVX1 INVX1_26 ( .A(w_C_29_), .Y(_465_) );
OR2X2 OR2X2_26 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_466_) );
NAND2X1 NAND2X1_51 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_467_) );
NAND3X1 NAND3X1_26 ( .A(_465_), .B(_467_), .C(_466_), .Y(_468_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_462_) );
AND2X2 AND2X2_26 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_463_) );
OAI21X1 OAI21X1_26 ( .A(_462_), .B(_463_), .C(w_C_29_), .Y(_464_) );
NAND2X1 NAND2X1_52 ( .A(_464_), .B(_468_), .Y(_286__29_) );
INVX1 INVX1_27 ( .A(w_C_30_), .Y(_472_) );
OR2X2 OR2X2_27 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_473_) );
NAND2X1 NAND2X1_53 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_474_) );
NAND3X1 NAND3X1_27 ( .A(_472_), .B(_474_), .C(_473_), .Y(_475_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_469_) );
AND2X2 AND2X2_27 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_470_) );
OAI21X1 OAI21X1_27 ( .A(_469_), .B(_470_), .C(w_C_30_), .Y(_471_) );
NAND2X1 NAND2X1_54 ( .A(_471_), .B(_475_), .Y(_286__30_) );
INVX1 INVX1_28 ( .A(w_C_31_), .Y(_479_) );
OR2X2 OR2X2_28 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_480_) );
NAND2X1 NAND2X1_55 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_481_) );
NAND3X1 NAND3X1_28 ( .A(_479_), .B(_481_), .C(_480_), .Y(_482_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_476_) );
AND2X2 AND2X2_28 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_477_) );
OAI21X1 OAI21X1_28 ( .A(_476_), .B(_477_), .C(w_C_31_), .Y(_478_) );
NAND2X1 NAND2X1_56 ( .A(_478_), .B(_482_), .Y(_286__31_) );
INVX1 INVX1_29 ( .A(w_C_32_), .Y(_486_) );
OR2X2 OR2X2_29 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_487_) );
NAND2X1 NAND2X1_57 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_488_) );
NAND3X1 NAND3X1_29 ( .A(_486_), .B(_488_), .C(_487_), .Y(_489_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_483_) );
AND2X2 AND2X2_29 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_484_) );
OAI21X1 OAI21X1_29 ( .A(_483_), .B(_484_), .C(w_C_32_), .Y(_485_) );
NAND2X1 NAND2X1_58 ( .A(_485_), .B(_489_), .Y(_286__32_) );
INVX1 INVX1_30 ( .A(w_C_33_), .Y(_493_) );
OR2X2 OR2X2_30 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_494_) );
NAND2X1 NAND2X1_59 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_495_) );
NAND3X1 NAND3X1_30 ( .A(_493_), .B(_495_), .C(_494_), .Y(_496_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_490_) );
AND2X2 AND2X2_30 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_491_) );
OAI21X1 OAI21X1_30 ( .A(_490_), .B(_491_), .C(w_C_33_), .Y(_492_) );
NAND2X1 NAND2X1_60 ( .A(_492_), .B(_496_), .Y(_286__33_) );
INVX1 INVX1_31 ( .A(w_C_34_), .Y(_500_) );
OR2X2 OR2X2_31 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_501_) );
NAND2X1 NAND2X1_61 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_502_) );
NAND3X1 NAND3X1_31 ( .A(_500_), .B(_502_), .C(_501_), .Y(_503_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_497_) );
AND2X2 AND2X2_31 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_498_) );
OAI21X1 OAI21X1_31 ( .A(_497_), .B(_498_), .C(w_C_34_), .Y(_499_) );
NAND2X1 NAND2X1_62 ( .A(_499_), .B(_503_), .Y(_286__34_) );
INVX1 INVX1_32 ( .A(w_C_35_), .Y(_507_) );
OR2X2 OR2X2_32 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_508_) );
NAND2X1 NAND2X1_63 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_509_) );
NAND3X1 NAND3X1_32 ( .A(_507_), .B(_509_), .C(_508_), .Y(_510_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_504_) );
AND2X2 AND2X2_32 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_505_) );
OAI21X1 OAI21X1_32 ( .A(_504_), .B(_505_), .C(w_C_35_), .Y(_506_) );
NAND2X1 NAND2X1_64 ( .A(_506_), .B(_510_), .Y(_286__35_) );
INVX1 INVX1_33 ( .A(w_C_36_), .Y(_514_) );
OR2X2 OR2X2_33 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_515_) );
NAND2X1 NAND2X1_65 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_516_) );
NAND3X1 NAND3X1_33 ( .A(_514_), .B(_516_), .C(_515_), .Y(_517_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_511_) );
AND2X2 AND2X2_33 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_512_) );
OAI21X1 OAI21X1_33 ( .A(_511_), .B(_512_), .C(w_C_36_), .Y(_513_) );
NAND2X1 NAND2X1_66 ( .A(_513_), .B(_517_), .Y(_286__36_) );
INVX1 INVX1_34 ( .A(w_C_37_), .Y(_521_) );
OR2X2 OR2X2_34 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_522_) );
NAND2X1 NAND2X1_67 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_523_) );
NAND3X1 NAND3X1_34 ( .A(_521_), .B(_523_), .C(_522_), .Y(_524_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_518_) );
AND2X2 AND2X2_34 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_519_) );
OAI21X1 OAI21X1_34 ( .A(_518_), .B(_519_), .C(w_C_37_), .Y(_520_) );
NAND2X1 NAND2X1_68 ( .A(_520_), .B(_524_), .Y(_286__37_) );
INVX1 INVX1_35 ( .A(w_C_38_), .Y(_528_) );
OR2X2 OR2X2_35 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_529_) );
NAND2X1 NAND2X1_69 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_530_) );
NAND3X1 NAND3X1_35 ( .A(_528_), .B(_530_), .C(_529_), .Y(_531_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_525_) );
AND2X2 AND2X2_35 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_526_) );
OAI21X1 OAI21X1_35 ( .A(_525_), .B(_526_), .C(w_C_38_), .Y(_527_) );
NAND2X1 NAND2X1_70 ( .A(_527_), .B(_531_), .Y(_286__38_) );
INVX1 INVX1_36 ( .A(w_C_39_), .Y(_535_) );
OR2X2 OR2X2_36 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_536_) );
NAND2X1 NAND2X1_71 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_537_) );
NAND3X1 NAND3X1_36 ( .A(_535_), .B(_537_), .C(_536_), .Y(_538_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_532_) );
AND2X2 AND2X2_36 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_533_) );
OAI21X1 OAI21X1_36 ( .A(_532_), .B(_533_), .C(w_C_39_), .Y(_534_) );
NAND2X1 NAND2X1_72 ( .A(_534_), .B(_538_), .Y(_286__39_) );
INVX1 INVX1_37 ( .A(w_C_40_), .Y(_542_) );
OR2X2 OR2X2_37 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_543_) );
NAND2X1 NAND2X1_73 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_544_) );
NAND3X1 NAND3X1_37 ( .A(_542_), .B(_544_), .C(_543_), .Y(_545_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_539_) );
AND2X2 AND2X2_37 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_540_) );
OAI21X1 OAI21X1_37 ( .A(_539_), .B(_540_), .C(w_C_40_), .Y(_541_) );
NAND2X1 NAND2X1_74 ( .A(_541_), .B(_545_), .Y(_286__40_) );
INVX1 INVX1_38 ( .A(w_C_41_), .Y(_549_) );
OR2X2 OR2X2_38 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_550_) );
NAND2X1 NAND2X1_75 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_551_) );
NAND3X1 NAND3X1_38 ( .A(_549_), .B(_551_), .C(_550_), .Y(_552_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_546_) );
AND2X2 AND2X2_38 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_547_) );
OAI21X1 OAI21X1_38 ( .A(_546_), .B(_547_), .C(w_C_41_), .Y(_548_) );
NAND2X1 NAND2X1_76 ( .A(_548_), .B(_552_), .Y(_286__41_) );
INVX1 INVX1_39 ( .A(w_C_42_), .Y(_556_) );
OR2X2 OR2X2_39 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_557_) );
NAND2X1 NAND2X1_77 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_558_) );
NAND3X1 NAND3X1_39 ( .A(_556_), .B(_558_), .C(_557_), .Y(_559_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_553_) );
AND2X2 AND2X2_39 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_554_) );
OAI21X1 OAI21X1_39 ( .A(_553_), .B(_554_), .C(w_C_42_), .Y(_555_) );
NAND2X1 NAND2X1_78 ( .A(_555_), .B(_559_), .Y(_286__42_) );
INVX1 INVX1_40 ( .A(w_C_43_), .Y(_563_) );
OR2X2 OR2X2_40 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_564_) );
NAND2X1 NAND2X1_79 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_565_) );
NAND3X1 NAND3X1_40 ( .A(_563_), .B(_565_), .C(_564_), .Y(_566_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_560_) );
AND2X2 AND2X2_40 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_561_) );
OAI21X1 OAI21X1_40 ( .A(_560_), .B(_561_), .C(w_C_43_), .Y(_562_) );
NAND2X1 NAND2X1_80 ( .A(_562_), .B(_566_), .Y(_286__43_) );
INVX1 INVX1_41 ( .A(w_C_44_), .Y(_570_) );
OR2X2 OR2X2_41 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_571_) );
NAND2X1 NAND2X1_81 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_572_) );
NAND3X1 NAND3X1_41 ( .A(_570_), .B(_572_), .C(_571_), .Y(_573_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_567_) );
AND2X2 AND2X2_41 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_568_) );
OAI21X1 OAI21X1_41 ( .A(_567_), .B(_568_), .C(w_C_44_), .Y(_569_) );
NAND2X1 NAND2X1_82 ( .A(_569_), .B(_573_), .Y(_286__44_) );
INVX1 INVX1_42 ( .A(w_C_45_), .Y(_577_) );
OR2X2 OR2X2_42 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_578_) );
NAND2X1 NAND2X1_83 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_579_) );
NAND3X1 NAND3X1_42 ( .A(_577_), .B(_579_), .C(_578_), .Y(_580_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_574_) );
AND2X2 AND2X2_42 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_575_) );
OAI21X1 OAI21X1_42 ( .A(_574_), .B(_575_), .C(w_C_45_), .Y(_576_) );
NAND2X1 NAND2X1_84 ( .A(_576_), .B(_580_), .Y(_286__45_) );
INVX1 INVX1_43 ( .A(w_C_46_), .Y(_584_) );
OR2X2 OR2X2_43 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_585_) );
NAND2X1 NAND2X1_85 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_586_) );
NAND3X1 NAND3X1_43 ( .A(_584_), .B(_586_), .C(_585_), .Y(_587_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_581_) );
AND2X2 AND2X2_43 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_582_) );
OAI21X1 OAI21X1_43 ( .A(_581_), .B(_582_), .C(w_C_46_), .Y(_583_) );
NAND2X1 NAND2X1_86 ( .A(_583_), .B(_587_), .Y(_286__46_) );
INVX1 INVX1_44 ( .A(w_C_47_), .Y(_591_) );
OR2X2 OR2X2_44 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_592_) );
NAND2X1 NAND2X1_87 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_593_) );
NAND3X1 NAND3X1_44 ( .A(_591_), .B(_593_), .C(_592_), .Y(_594_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_588_) );
AND2X2 AND2X2_44 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_589_) );
OAI21X1 OAI21X1_44 ( .A(_588_), .B(_589_), .C(w_C_47_), .Y(_590_) );
NAND2X1 NAND2X1_88 ( .A(_590_), .B(_594_), .Y(_286__47_) );
INVX1 INVX1_45 ( .A(w_C_48_), .Y(_598_) );
OR2X2 OR2X2_45 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_599_) );
NAND2X1 NAND2X1_89 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_600_) );
NAND3X1 NAND3X1_45 ( .A(_598_), .B(_600_), .C(_599_), .Y(_601_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_595_) );
AND2X2 AND2X2_45 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_596_) );
OAI21X1 OAI21X1_45 ( .A(_595_), .B(_596_), .C(w_C_48_), .Y(_597_) );
NAND2X1 NAND2X1_90 ( .A(_597_), .B(_601_), .Y(_286__48_) );
INVX1 INVX1_46 ( .A(w_C_49_), .Y(_605_) );
OR2X2 OR2X2_46 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_606_) );
NAND2X1 NAND2X1_91 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_607_) );
NAND3X1 NAND3X1_46 ( .A(_605_), .B(_607_), .C(_606_), .Y(_608_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_602_) );
AND2X2 AND2X2_46 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_603_) );
OAI21X1 OAI21X1_46 ( .A(_602_), .B(_603_), .C(w_C_49_), .Y(_604_) );
NAND2X1 NAND2X1_92 ( .A(_604_), .B(_608_), .Y(_286__49_) );
INVX1 INVX1_47 ( .A(gnd), .Y(_612_) );
OR2X2 OR2X2_47 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_613_) );
NAND2X1 NAND2X1_93 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_614_) );
NAND3X1 NAND3X1_47 ( .A(_612_), .B(_614_), .C(_613_), .Y(_615_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_609_) );
AND2X2 AND2X2_47 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_610_) );
OAI21X1 OAI21X1_47 ( .A(_609_), .B(_610_), .C(gnd), .Y(_611_) );
NAND2X1 NAND2X1_94 ( .A(_611_), .B(_615_), .Y(_286__0_) );
INVX1 INVX1_48 ( .A(w_C_1_), .Y(_619_) );
OR2X2 OR2X2_48 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_620_) );
NAND2X1 NAND2X1_95 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_621_) );
NAND3X1 NAND3X1_48 ( .A(_619_), .B(_621_), .C(_620_), .Y(_622_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_616_) );
AND2X2 AND2X2_48 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_617_) );
OAI21X1 OAI21X1_48 ( .A(_616_), .B(_617_), .C(w_C_1_), .Y(_618_) );
NAND2X1 NAND2X1_96 ( .A(_618_), .B(_622_), .Y(_286__1_) );
INVX1 INVX1_49 ( .A(w_C_2_), .Y(_626_) );
OR2X2 OR2X2_49 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_627_) );
NAND2X1 NAND2X1_97 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_628_) );
NAND3X1 NAND3X1_49 ( .A(_626_), .B(_628_), .C(_627_), .Y(_629_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_623_) );
AND2X2 AND2X2_49 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_624_) );
OAI21X1 OAI21X1_49 ( .A(_623_), .B(_624_), .C(w_C_2_), .Y(_625_) );
NAND2X1 NAND2X1_98 ( .A(_625_), .B(_629_), .Y(_286__2_) );
INVX1 INVX1_50 ( .A(w_C_3_), .Y(_633_) );
OR2X2 OR2X2_50 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_634_) );
NAND2X1 NAND2X1_99 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_635_) );
NAND3X1 NAND3X1_50 ( .A(_633_), .B(_635_), .C(_634_), .Y(_636_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_630_) );
AND2X2 AND2X2_50 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_631_) );
OAI21X1 OAI21X1_50 ( .A(_630_), .B(_631_), .C(w_C_3_), .Y(_632_) );
NAND2X1 NAND2X1_100 ( .A(_632_), .B(_636_), .Y(_286__3_) );
INVX1 INVX1_51 ( .A(i_add1[33]), .Y(_190_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_191_) );
INVX1 INVX1_52 ( .A(_191_), .Y(_192_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_193_) );
INVX1 INVX1_53 ( .A(_193_), .Y(_194_) );
NAND3X1 NAND3X1_51 ( .A(_192_), .B(_194_), .C(_187_), .Y(_195_) );
OAI21X1 OAI21X1_51 ( .A(_189_), .B(_190_), .C(_195_), .Y(w_C_34_) );
NOR2X1 NOR2X1_53 ( .A(_189_), .B(_190_), .Y(_196_) );
INVX1 INVX1_54 ( .A(_196_), .Y(_197_) );
AND2X2 AND2X2_51 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_198_) );
INVX1 INVX1_55 ( .A(_198_), .Y(_199_) );
NAND3X1 NAND3X1_52 ( .A(_197_), .B(_199_), .C(_195_), .Y(_200_) );
OAI21X1 OAI21X1_52 ( .A(i_add2[34]), .B(i_add1[34]), .C(_200_), .Y(_201_) );
INVX1 INVX1_56 ( .A(_201_), .Y(w_C_35_) );
INVX1 INVX1_57 ( .A(i_add2[35]), .Y(_202_) );
INVX1 INVX1_58 ( .A(i_add1[35]), .Y(_203_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_204_) );
INVX1 INVX1_59 ( .A(_204_), .Y(_205_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_206_) );
INVX1 INVX1_60 ( .A(_206_), .Y(_207_) );
NAND3X1 NAND3X1_53 ( .A(_205_), .B(_207_), .C(_200_), .Y(_208_) );
OAI21X1 OAI21X1_53 ( .A(_202_), .B(_203_), .C(_208_), .Y(w_C_36_) );
NOR2X1 NOR2X1_56 ( .A(_202_), .B(_203_), .Y(_209_) );
INVX1 INVX1_61 ( .A(_209_), .Y(_210_) );
AND2X2 AND2X2_52 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_211_) );
INVX1 INVX1_62 ( .A(_211_), .Y(_212_) );
NAND3X1 NAND3X1_54 ( .A(_210_), .B(_212_), .C(_208_), .Y(_213_) );
OAI21X1 OAI21X1_54 ( .A(i_add2[36]), .B(i_add1[36]), .C(_213_), .Y(_214_) );
INVX1 INVX1_63 ( .A(_214_), .Y(w_C_37_) );
INVX1 INVX1_64 ( .A(i_add2[37]), .Y(_215_) );
INVX1 INVX1_65 ( .A(i_add1[37]), .Y(_216_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_217_) );
INVX1 INVX1_66 ( .A(_217_), .Y(_218_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_219_) );
INVX1 INVX1_67 ( .A(_219_), .Y(_220_) );
NAND3X1 NAND3X1_55 ( .A(_218_), .B(_220_), .C(_213_), .Y(_221_) );
OAI21X1 OAI21X1_55 ( .A(_215_), .B(_216_), .C(_221_), .Y(w_C_38_) );
NOR2X1 NOR2X1_59 ( .A(_215_), .B(_216_), .Y(_222_) );
INVX1 INVX1_68 ( .A(_222_), .Y(_223_) );
AND2X2 AND2X2_53 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_224_) );
INVX1 INVX1_69 ( .A(_224_), .Y(_225_) );
NAND3X1 NAND3X1_56 ( .A(_223_), .B(_225_), .C(_221_), .Y(_226_) );
OAI21X1 OAI21X1_56 ( .A(i_add2[38]), .B(i_add1[38]), .C(_226_), .Y(_227_) );
INVX1 INVX1_70 ( .A(_227_), .Y(w_C_39_) );
INVX1 INVX1_71 ( .A(i_add2[39]), .Y(_228_) );
INVX1 INVX1_72 ( .A(i_add1[39]), .Y(_229_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_230_) );
INVX1 INVX1_73 ( .A(_230_), .Y(_231_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_232_) );
INVX1 INVX1_74 ( .A(_232_), .Y(_233_) );
NAND3X1 NAND3X1_57 ( .A(_231_), .B(_233_), .C(_226_), .Y(_234_) );
OAI21X1 OAI21X1_57 ( .A(_228_), .B(_229_), .C(_234_), .Y(w_C_40_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_235_) );
INVX1 INVX1_75 ( .A(_235_), .Y(_236_) );
NOR2X1 NOR2X1_63 ( .A(_228_), .B(_229_), .Y(_237_) );
INVX1 INVX1_76 ( .A(_237_), .Y(_238_) );
NAND2X1 NAND2X1_101 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_239_) );
NAND3X1 NAND3X1_58 ( .A(_238_), .B(_239_), .C(_234_), .Y(_240_) );
AND2X2 AND2X2_54 ( .A(_240_), .B(_236_), .Y(w_C_41_) );
INVX1 INVX1_77 ( .A(i_add2[41]), .Y(_241_) );
INVX1 INVX1_78 ( .A(i_add1[41]), .Y(_242_) );
NAND2X1 NAND2X1_102 ( .A(_241_), .B(_242_), .Y(_243_) );
NAND3X1 NAND3X1_59 ( .A(_236_), .B(_243_), .C(_240_), .Y(_244_) );
OAI21X1 OAI21X1_58 ( .A(_241_), .B(_242_), .C(_244_), .Y(w_C_42_) );
INVX1 INVX1_79 ( .A(i_add2[42]), .Y(_245_) );
INVX1 INVX1_80 ( .A(i_add1[42]), .Y(_246_) );
OAI21X1 OAI21X1_59 ( .A(i_add2[42]), .B(i_add1[42]), .C(w_C_42_), .Y(_247_) );
OAI21X1 OAI21X1_60 ( .A(_245_), .B(_246_), .C(_247_), .Y(w_C_43_) );
INVX1 INVX1_81 ( .A(i_add2[43]), .Y(_248_) );
INVX1 INVX1_82 ( .A(i_add1[43]), .Y(_249_) );
NOR2X1 NOR2X1_64 ( .A(_248_), .B(_249_), .Y(_250_) );
OR2X2 OR2X2_51 ( .A(w_C_43_), .B(_250_), .Y(_251_) );
OAI21X1 OAI21X1_61 ( .A(i_add2[43]), .B(i_add1[43]), .C(_251_), .Y(_252_) );
INVX1 INVX1_83 ( .A(_252_), .Y(w_C_44_) );
INVX1 INVX1_84 ( .A(_250_), .Y(_253_) );
NAND2X1 NAND2X1_103 ( .A(_245_), .B(_246_), .Y(_254_) );
NAND2X1 NAND2X1_104 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_255_) );
NAND2X1 NAND2X1_105 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_256_) );
NAND3X1 NAND3X1_60 ( .A(_255_), .B(_256_), .C(_244_), .Y(_257_) );
NAND2X1 NAND2X1_106 ( .A(_248_), .B(_249_), .Y(_258_) );
NAND3X1 NAND3X1_61 ( .A(_254_), .B(_258_), .C(_257_), .Y(_259_) );
NAND2X1 NAND2X1_107 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_260_) );
NAND3X1 NAND3X1_62 ( .A(_253_), .B(_260_), .C(_259_), .Y(_261_) );
OAI21X1 OAI21X1_62 ( .A(i_add2[44]), .B(i_add1[44]), .C(_261_), .Y(_262_) );
INVX1 INVX1_85 ( .A(_262_), .Y(w_C_45_) );
INVX1 INVX1_86 ( .A(i_add2[45]), .Y(_263_) );
INVX1 INVX1_87 ( .A(i_add1[45]), .Y(_264_) );
OAI21X1 OAI21X1_63 ( .A(_263_), .B(_264_), .C(_262_), .Y(_265_) );
OAI21X1 OAI21X1_64 ( .A(i_add2[45]), .B(i_add1[45]), .C(_265_), .Y(_266_) );
INVX1 INVX1_88 ( .A(_266_), .Y(w_C_46_) );
NAND2X1 NAND2X1_108 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_267_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_268_) );
OAI21X1 OAI21X1_65 ( .A(_268_), .B(_266_), .C(_267_), .Y(w_C_47_) );
NAND2X1 NAND2X1_109 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_269_) );
INVX1 INVX1_89 ( .A(_268_), .Y(_270_) );
NOR2X1 NOR2X1_66 ( .A(_263_), .B(_264_), .Y(_271_) );
INVX1 INVX1_90 ( .A(_271_), .Y(_272_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_273_) );
INVX1 INVX1_91 ( .A(_273_), .Y(_274_) );
NAND2X1 NAND2X1_110 ( .A(_263_), .B(_264_), .Y(_275_) );
NAND3X1 NAND3X1_63 ( .A(_274_), .B(_275_), .C(_261_), .Y(_276_) );
NAND3X1 NAND3X1_64 ( .A(_272_), .B(_267_), .C(_276_), .Y(_277_) );
OR2X2 OR2X2_52 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_278_) );
NAND3X1 NAND3X1_65 ( .A(_270_), .B(_278_), .C(_277_), .Y(_279_) );
NAND2X1 NAND2X1_111 ( .A(_269_), .B(_279_), .Y(w_C_48_) );
OR2X2 OR2X2_53 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_280_) );
NAND2X1 NAND2X1_112 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_281_) );
NAND3X1 NAND3X1_66 ( .A(_269_), .B(_281_), .C(_279_), .Y(_282_) );
AND2X2 AND2X2_55 ( .A(_282_), .B(_280_), .Y(w_C_49_) );
NAND2X1 NAND2X1_113 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_283_) );
OR2X2 OR2X2_54 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_284_) );
NAND3X1 NAND3X1_67 ( .A(_280_), .B(_284_), .C(_282_), .Y(_285_) );
NAND2X1 NAND2X1_114 ( .A(_283_), .B(_285_), .Y(w_C_50_) );
NAND2X1 NAND2X1_115 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_92 ( .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_68 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_69 ( .A(_1_), .B(_2_), .Y(w_C_2_) );
INVX1 INVX1_93 ( .A(i_add2[2]), .Y(_3_) );
INVX1 INVX1_94 ( .A(i_add1[2]), .Y(_4_) );
NAND2X1 NAND2X1_116 ( .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_117 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
OAI21X1 OAI21X1_66 ( .A(_1_), .B(_2_), .C(_6_), .Y(_7_) );
AND2X2 AND2X2_56 ( .A(_7_), .B(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_118 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
OR2X2 OR2X2_55 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_68 ( .A(_5_), .B(_9_), .C(_7_), .Y(_10_) );
NAND2X1 NAND2X1_119 ( .A(_8_), .B(_10_), .Y(w_C_4_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
INVX1 INVX1_95 ( .A(_11_), .Y(_12_) );
NAND2X1 NAND2X1_120 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
NAND3X1 NAND3X1_69 ( .A(_8_), .B(_13_), .C(_10_), .Y(_14_) );
AND2X2 AND2X2_57 ( .A(_14_), .B(_12_), .Y(w_C_5_) );
INVX1 INVX1_96 ( .A(i_add2[5]), .Y(_15_) );
INVX1 INVX1_97 ( .A(i_add1[5]), .Y(_16_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_17_) );
INVX1 INVX1_98 ( .A(_17_), .Y(_18_) );
NAND3X1 NAND3X1_70 ( .A(_12_), .B(_18_), .C(_14_), .Y(_19_) );
OAI21X1 OAI21X1_67 ( .A(_15_), .B(_16_), .C(_19_), .Y(w_C_6_) );
NOR2X1 NOR2X1_72 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_20_) );
INVX1 INVX1_99 ( .A(_20_), .Y(_21_) );
NOR2X1 NOR2X1_73 ( .A(_15_), .B(_16_), .Y(_22_) );
INVX1 INVX1_100 ( .A(_22_), .Y(_23_) );
AND2X2 AND2X2_58 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_24_) );
INVX1 INVX1_101 ( .A(_24_), .Y(_25_) );
NAND3X1 NAND3X1_71 ( .A(_23_), .B(_25_), .C(_19_), .Y(_26_) );
AND2X2 AND2X2_59 ( .A(_26_), .B(_21_), .Y(w_C_7_) );
AND2X2 AND2X2_60 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_27_) );
INVX1 INVX1_102 ( .A(_27_), .Y(_28_) );
NOR2X1 NOR2X1_74 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_29_) );
INVX1 INVX1_103 ( .A(_29_), .Y(_30_) );
NAND3X1 NAND3X1_72 ( .A(_21_), .B(_30_), .C(_26_), .Y(_31_) );
AND2X2 AND2X2_61 ( .A(_31_), .B(_28_), .Y(_32_) );
INVX1 INVX1_104 ( .A(_32_), .Y(w_C_8_) );
AND2X2 AND2X2_62 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_33_) );
INVX1 INVX1_105 ( .A(_33_), .Y(_34_) );
NOR2X1 NOR2X1_75 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_35_) );
OAI21X1 OAI21X1_68 ( .A(_35_), .B(_32_), .C(_34_), .Y(w_C_9_) );
AND2X2 AND2X2_63 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_36_) );
INVX1 INVX1_106 ( .A(_36_), .Y(_37_) );
INVX1 INVX1_107 ( .A(_35_), .Y(_38_) );
NAND3X1 NAND3X1_73 ( .A(_28_), .B(_34_), .C(_31_), .Y(_39_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_40_) );
INVX1 INVX1_108 ( .A(_40_), .Y(_41_) );
NAND3X1 NAND3X1_74 ( .A(_38_), .B(_41_), .C(_39_), .Y(_42_) );
AND2X2 AND2X2_64 ( .A(_42_), .B(_37_), .Y(_43_) );
INVX1 INVX1_109 ( .A(_43_), .Y(w_C_10_) );
AND2X2 AND2X2_65 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_44_) );
INVX1 INVX1_110 ( .A(_44_), .Y(_45_) );
NOR2X1 NOR2X1_77 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_46_) );
OAI21X1 OAI21X1_69 ( .A(_46_), .B(_43_), .C(_45_), .Y(w_C_11_) );
AND2X2 AND2X2_66 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_47_) );
INVX1 INVX1_111 ( .A(_47_), .Y(_48_) );
INVX1 INVX1_112 ( .A(_46_), .Y(_49_) );
NAND3X1 NAND3X1_75 ( .A(_37_), .B(_45_), .C(_42_), .Y(_50_) );
NOR2X1 NOR2X1_78 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_51_) );
INVX1 INVX1_113 ( .A(_51_), .Y(_52_) );
NAND3X1 NAND3X1_76 ( .A(_49_), .B(_52_), .C(_50_), .Y(_53_) );
AND2X2 AND2X2_67 ( .A(_53_), .B(_48_), .Y(_54_) );
INVX1 INVX1_114 ( .A(_54_), .Y(w_C_12_) );
AND2X2 AND2X2_68 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_55_) );
INVX1 INVX1_115 ( .A(_55_), .Y(_56_) );
NAND3X1 NAND3X1_77 ( .A(_48_), .B(_56_), .C(_53_), .Y(_57_) );
OAI21X1 OAI21X1_70 ( .A(i_add2[12]), .B(i_add1[12]), .C(_57_), .Y(_58_) );
INVX1 INVX1_116 ( .A(_58_), .Y(w_C_13_) );
INVX1 INVX1_117 ( .A(i_add2[13]), .Y(_59_) );
INVX1 INVX1_118 ( .A(i_add1[13]), .Y(_60_) );
NOR2X1 NOR2X1_79 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_61_) );
INVX1 INVX1_119 ( .A(_61_), .Y(_62_) );
NOR2X1 NOR2X1_80 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_63_) );
INVX1 INVX1_120 ( .A(_63_), .Y(_64_) );
NAND3X1 NAND3X1_78 ( .A(_62_), .B(_64_), .C(_57_), .Y(_65_) );
OAI21X1 OAI21X1_71 ( .A(_59_), .B(_60_), .C(_65_), .Y(w_C_14_) );
NOR2X1 NOR2X1_81 ( .A(_59_), .B(_60_), .Y(_66_) );
INVX1 INVX1_121 ( .A(_66_), .Y(_67_) );
AND2X2 AND2X2_69 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_68_) );
INVX1 INVX1_122 ( .A(_68_), .Y(_69_) );
NAND3X1 NAND3X1_79 ( .A(_67_), .B(_69_), .C(_65_), .Y(_70_) );
OAI21X1 OAI21X1_72 ( .A(i_add2[14]), .B(i_add1[14]), .C(_70_), .Y(_71_) );
INVX1 INVX1_123 ( .A(_71_), .Y(w_C_15_) );
INVX1 INVX1_124 ( .A(i_add2[15]), .Y(_72_) );
INVX1 INVX1_125 ( .A(i_add1[15]), .Y(_73_) );
NOR2X1 NOR2X1_82 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_74_) );
INVX1 INVX1_126 ( .A(_74_), .Y(_75_) );
NOR2X1 NOR2X1_83 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_76_) );
INVX1 INVX1_127 ( .A(_76_), .Y(_77_) );
NAND3X1 NAND3X1_80 ( .A(_75_), .B(_77_), .C(_70_), .Y(_78_) );
OAI21X1 OAI21X1_73 ( .A(_72_), .B(_73_), .C(_78_), .Y(w_C_16_) );
NOR2X1 NOR2X1_84 ( .A(_72_), .B(_73_), .Y(_79_) );
INVX1 INVX1_128 ( .A(_79_), .Y(_80_) );
AND2X2 AND2X2_70 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_81_) );
INVX1 INVX1_129 ( .A(_81_), .Y(_82_) );
NAND3X1 NAND3X1_81 ( .A(_80_), .B(_82_), .C(_78_), .Y(_83_) );
OAI21X1 OAI21X1_74 ( .A(i_add2[16]), .B(i_add1[16]), .C(_83_), .Y(_84_) );
INVX1 INVX1_130 ( .A(_84_), .Y(w_C_17_) );
INVX1 INVX1_131 ( .A(i_add2[17]), .Y(_85_) );
INVX1 INVX1_132 ( .A(i_add1[17]), .Y(_86_) );
NOR2X1 NOR2X1_85 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_87_) );
INVX1 INVX1_133 ( .A(_87_), .Y(_88_) );
NOR2X1 NOR2X1_86 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_89_) );
INVX1 INVX1_134 ( .A(_89_), .Y(_90_) );
NAND3X1 NAND3X1_82 ( .A(_88_), .B(_90_), .C(_83_), .Y(_91_) );
OAI21X1 OAI21X1_75 ( .A(_85_), .B(_86_), .C(_91_), .Y(w_C_18_) );
NOR2X1 NOR2X1_87 ( .A(_85_), .B(_86_), .Y(_92_) );
INVX1 INVX1_135 ( .A(_92_), .Y(_93_) );
AND2X2 AND2X2_71 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_94_) );
INVX1 INVX1_136 ( .A(_94_), .Y(_95_) );
NAND3X1 NAND3X1_83 ( .A(_93_), .B(_95_), .C(_91_), .Y(_96_) );
OAI21X1 OAI21X1_76 ( .A(i_add2[18]), .B(i_add1[18]), .C(_96_), .Y(_97_) );
INVX1 INVX1_137 ( .A(_97_), .Y(w_C_19_) );
INVX1 INVX1_138 ( .A(i_add2[19]), .Y(_98_) );
INVX1 INVX1_139 ( .A(i_add1[19]), .Y(_99_) );
NOR2X1 NOR2X1_88 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_100_) );
INVX1 INVX1_140 ( .A(_100_), .Y(_101_) );
NOR2X1 NOR2X1_89 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_102_) );
INVX1 INVX1_141 ( .A(_102_), .Y(_103_) );
NAND3X1 NAND3X1_84 ( .A(_101_), .B(_103_), .C(_96_), .Y(_104_) );
OAI21X1 OAI21X1_77 ( .A(_98_), .B(_99_), .C(_104_), .Y(w_C_20_) );
NOR2X1 NOR2X1_90 ( .A(_98_), .B(_99_), .Y(_105_) );
INVX1 INVX1_142 ( .A(_105_), .Y(_106_) );
AND2X2 AND2X2_72 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_107_) );
INVX1 INVX1_143 ( .A(_107_), .Y(_108_) );
NAND3X1 NAND3X1_85 ( .A(_106_), .B(_108_), .C(_104_), .Y(_109_) );
OAI21X1 OAI21X1_78 ( .A(i_add2[20]), .B(i_add1[20]), .C(_109_), .Y(_110_) );
INVX1 INVX1_144 ( .A(_110_), .Y(w_C_21_) );
INVX1 INVX1_145 ( .A(i_add2[21]), .Y(_111_) );
INVX1 INVX1_146 ( .A(i_add1[21]), .Y(_112_) );
NOR2X1 NOR2X1_91 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_113_) );
INVX1 INVX1_147 ( .A(_113_), .Y(_114_) );
NOR2X1 NOR2X1_92 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_115_) );
INVX1 INVX1_148 ( .A(_115_), .Y(_116_) );
NAND3X1 NAND3X1_86 ( .A(_114_), .B(_116_), .C(_109_), .Y(_117_) );
OAI21X1 OAI21X1_79 ( .A(_111_), .B(_112_), .C(_117_), .Y(w_C_22_) );
NOR2X1 NOR2X1_93 ( .A(_111_), .B(_112_), .Y(_118_) );
INVX1 INVX1_149 ( .A(_118_), .Y(_119_) );
AND2X2 AND2X2_73 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_120_) );
INVX1 INVX1_150 ( .A(_120_), .Y(_121_) );
NAND3X1 NAND3X1_87 ( .A(_119_), .B(_121_), .C(_117_), .Y(_122_) );
OAI21X1 OAI21X1_80 ( .A(i_add2[22]), .B(i_add1[22]), .C(_122_), .Y(_123_) );
INVX1 INVX1_151 ( .A(_123_), .Y(w_C_23_) );
INVX1 INVX1_152 ( .A(i_add2[23]), .Y(_124_) );
INVX1 INVX1_153 ( .A(i_add1[23]), .Y(_125_) );
NOR2X1 NOR2X1_94 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_126_) );
INVX1 INVX1_154 ( .A(_126_), .Y(_127_) );
NOR2X1 NOR2X1_95 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_128_) );
INVX1 INVX1_155 ( .A(_128_), .Y(_129_) );
NAND3X1 NAND3X1_88 ( .A(_127_), .B(_129_), .C(_122_), .Y(_130_) );
OAI21X1 OAI21X1_81 ( .A(_124_), .B(_125_), .C(_130_), .Y(w_C_24_) );
NOR2X1 NOR2X1_96 ( .A(_124_), .B(_125_), .Y(_131_) );
INVX1 INVX1_156 ( .A(_131_), .Y(_132_) );
AND2X2 AND2X2_74 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_133_) );
INVX1 INVX1_157 ( .A(_133_), .Y(_134_) );
NAND3X1 NAND3X1_89 ( .A(_132_), .B(_134_), .C(_130_), .Y(_135_) );
OAI21X1 OAI21X1_82 ( .A(i_add2[24]), .B(i_add1[24]), .C(_135_), .Y(_136_) );
INVX1 INVX1_158 ( .A(_136_), .Y(w_C_25_) );
INVX1 INVX1_159 ( .A(i_add2[25]), .Y(_137_) );
INVX1 INVX1_160 ( .A(i_add1[25]), .Y(_138_) );
NOR2X1 NOR2X1_97 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_139_) );
INVX1 INVX1_161 ( .A(_139_), .Y(_140_) );
NOR2X1 NOR2X1_98 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_141_) );
INVX1 INVX1_162 ( .A(_141_), .Y(_142_) );
NAND3X1 NAND3X1_90 ( .A(_140_), .B(_142_), .C(_135_), .Y(_143_) );
OAI21X1 OAI21X1_83 ( .A(_137_), .B(_138_), .C(_143_), .Y(w_C_26_) );
NOR2X1 NOR2X1_99 ( .A(_137_), .B(_138_), .Y(_144_) );
INVX1 INVX1_163 ( .A(_144_), .Y(_145_) );
AND2X2 AND2X2_75 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_146_) );
INVX1 INVX1_164 ( .A(_146_), .Y(_147_) );
NAND3X1 NAND3X1_91 ( .A(_145_), .B(_147_), .C(_143_), .Y(_148_) );
OAI21X1 OAI21X1_84 ( .A(i_add2[26]), .B(i_add1[26]), .C(_148_), .Y(_149_) );
INVX1 INVX1_165 ( .A(_149_), .Y(w_C_27_) );
INVX1 INVX1_166 ( .A(i_add2[27]), .Y(_150_) );
INVX1 INVX1_167 ( .A(i_add1[27]), .Y(_151_) );
NOR2X1 NOR2X1_100 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_152_) );
INVX1 INVX1_168 ( .A(_152_), .Y(_153_) );
NOR2X1 NOR2X1_101 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_154_) );
INVX1 INVX1_169 ( .A(_154_), .Y(_155_) );
NAND3X1 NAND3X1_92 ( .A(_153_), .B(_155_), .C(_148_), .Y(_156_) );
OAI21X1 OAI21X1_85 ( .A(_150_), .B(_151_), .C(_156_), .Y(w_C_28_) );
NOR2X1 NOR2X1_102 ( .A(_150_), .B(_151_), .Y(_157_) );
INVX1 INVX1_170 ( .A(_157_), .Y(_158_) );
AND2X2 AND2X2_76 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_159_) );
INVX1 INVX1_171 ( .A(_159_), .Y(_160_) );
NAND3X1 NAND3X1_93 ( .A(_158_), .B(_160_), .C(_156_), .Y(_161_) );
OAI21X1 OAI21X1_86 ( .A(i_add2[28]), .B(i_add1[28]), .C(_161_), .Y(_162_) );
INVX1 INVX1_172 ( .A(_162_), .Y(w_C_29_) );
INVX1 INVX1_173 ( .A(i_add2[29]), .Y(_163_) );
INVX1 INVX1_174 ( .A(i_add1[29]), .Y(_164_) );
NOR2X1 NOR2X1_103 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_165_) );
INVX1 INVX1_175 ( .A(_165_), .Y(_166_) );
NOR2X1 NOR2X1_104 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_167_) );
INVX1 INVX1_176 ( .A(_167_), .Y(_168_) );
NAND3X1 NAND3X1_94 ( .A(_166_), .B(_168_), .C(_161_), .Y(_169_) );
OAI21X1 OAI21X1_87 ( .A(_163_), .B(_164_), .C(_169_), .Y(w_C_30_) );
NOR2X1 NOR2X1_105 ( .A(_163_), .B(_164_), .Y(_170_) );
INVX1 INVX1_177 ( .A(_170_), .Y(_171_) );
AND2X2 AND2X2_77 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_172_) );
INVX1 INVX1_178 ( .A(_172_), .Y(_173_) );
NAND3X1 NAND3X1_95 ( .A(_171_), .B(_173_), .C(_169_), .Y(_174_) );
OAI21X1 OAI21X1_88 ( .A(i_add2[30]), .B(i_add1[30]), .C(_174_), .Y(_175_) );
INVX1 INVX1_179 ( .A(_175_), .Y(w_C_31_) );
INVX1 INVX1_180 ( .A(i_add2[31]), .Y(_176_) );
INVX1 INVX1_181 ( .A(i_add1[31]), .Y(_177_) );
NOR2X1 NOR2X1_106 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_178_) );
INVX1 INVX1_182 ( .A(_178_), .Y(_179_) );
NOR2X1 NOR2X1_107 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_180_) );
INVX1 INVX1_183 ( .A(_180_), .Y(_181_) );
NAND3X1 NAND3X1_96 ( .A(_179_), .B(_181_), .C(_174_), .Y(_182_) );
OAI21X1 OAI21X1_89 ( .A(_176_), .B(_177_), .C(_182_), .Y(w_C_32_) );
NOR2X1 NOR2X1_108 ( .A(_176_), .B(_177_), .Y(_183_) );
INVX1 INVX1_184 ( .A(_183_), .Y(_184_) );
AND2X2 AND2X2_78 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_185_) );
INVX1 INVX1_185 ( .A(_185_), .Y(_186_) );
NAND3X1 NAND3X1_97 ( .A(_184_), .B(_186_), .C(_182_), .Y(_187_) );
OAI21X1 OAI21X1_90 ( .A(i_add2[32]), .B(i_add1[32]), .C(_187_), .Y(_188_) );
INVX1 INVX1_186 ( .A(_188_), .Y(w_C_33_) );
INVX1 INVX1_187 ( .A(i_add2[33]), .Y(_189_) );
BUFX2 BUFX2_25 ( .A(_286__0_), .Y(o_result[0]) );
BUFX2 BUFX2_26 ( .A(_286__1_), .Y(o_result[1]) );
BUFX2 BUFX2_27 ( .A(_286__2_), .Y(o_result[2]) );
BUFX2 BUFX2_28 ( .A(_286__3_), .Y(o_result[3]) );
BUFX2 BUFX2_29 ( .A(_286__4_), .Y(o_result[4]) );
BUFX2 BUFX2_30 ( .A(_286__5_), .Y(o_result[5]) );
BUFX2 BUFX2_31 ( .A(_286__6_), .Y(o_result[6]) );
BUFX2 BUFX2_32 ( .A(_286__7_), .Y(o_result[7]) );
BUFX2 BUFX2_33 ( .A(_286__8_), .Y(o_result[8]) );
BUFX2 BUFX2_34 ( .A(_286__9_), .Y(o_result[9]) );
BUFX2 BUFX2_35 ( .A(_286__10_), .Y(o_result[10]) );
BUFX2 BUFX2_36 ( .A(_286__11_), .Y(o_result[11]) );
BUFX2 BUFX2_37 ( .A(_286__12_), .Y(o_result[12]) );
BUFX2 BUFX2_38 ( .A(_286__13_), .Y(o_result[13]) );
BUFX2 BUFX2_39 ( .A(_286__14_), .Y(o_result[14]) );
BUFX2 BUFX2_40 ( .A(_286__15_), .Y(o_result[15]) );
BUFX2 BUFX2_41 ( .A(_286__16_), .Y(o_result[16]) );
BUFX2 BUFX2_42 ( .A(_286__17_), .Y(o_result[17]) );
BUFX2 BUFX2_43 ( .A(_286__18_), .Y(o_result[18]) );
BUFX2 BUFX2_44 ( .A(_286__19_), .Y(o_result[19]) );
BUFX2 BUFX2_45 ( .A(_286__20_), .Y(o_result[20]) );
BUFX2 BUFX2_46 ( .A(_286__21_), .Y(o_result[21]) );
BUFX2 BUFX2_47 ( .A(_286__22_), .Y(o_result[22]) );
BUFX2 BUFX2_48 ( .A(_286__23_), .Y(o_result[23]) );
BUFX2 BUFX2_49 ( .A(_286__24_), .Y(o_result[24]) );
BUFX2 BUFX2_50 ( .A(_286__25_), .Y(o_result[25]) );
BUFX2 BUFX2_51 ( .A(_286__26_), .Y(o_result[26]) );
BUFX2 BUFX2_52 ( .A(w_C_50_), .Y(_286__50_) );
BUFX2 BUFX2_53 ( .A(gnd), .Y(w_C_0_) );
endmodule
