module cla_30bit (i_add1, i_add2, o_result);

input [29:0] i_add1;
input [29:0] i_add2;
output [30:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_159_) );
INVX1 INVX1_1 ( .A(_159_), .Y(w_C_1_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_160_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_161_) );
NOR2X1 NOR2X1_2 ( .A(_160_), .B(_161_), .Y(w_C_2_) );
INVX1 INVX1_2 ( .A(i_add2[2]), .Y(_162_) );
INVX1 INVX1_3 ( .A(i_add1[2]), .Y(_163_) );
NAND2X1 NAND2X1_2 ( .A(_162_), .B(_163_), .Y(_164_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_165_) );
OAI21X1 OAI21X1_1 ( .A(_160_), .B(_161_), .C(_165_), .Y(_0_) );
AND2X2 AND2X2_1 ( .A(_0_), .B(_164_), .Y(w_C_3_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_1_) );
OR2X2 OR2X2_1 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_2_) );
NAND3X1 NAND3X1_1 ( .A(_164_), .B(_2_), .C(_0_), .Y(_3_) );
NAND2X1 NAND2X1_5 ( .A(_1_), .B(_3_), .Y(w_C_4_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_4_) );
NAND3X1 NAND3X1_2 ( .A(_1_), .B(_4_), .C(_3_), .Y(_5_) );
OAI21X1 OAI21X1_2 ( .A(i_add2[4]), .B(i_add1[4]), .C(_5_), .Y(_6_) );
INVX1 INVX1_4 ( .A(_6_), .Y(w_C_5_) );
INVX1 INVX1_5 ( .A(i_add2[5]), .Y(_7_) );
INVX1 INVX1_6 ( .A(i_add1[5]), .Y(_8_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_9_) );
INVX1 INVX1_7 ( .A(_9_), .Y(_10_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_11_) );
INVX1 INVX1_8 ( .A(_11_), .Y(_12_) );
NAND3X1 NAND3X1_3 ( .A(_10_), .B(_12_), .C(_5_), .Y(_13_) );
OAI21X1 OAI21X1_3 ( .A(_7_), .B(_8_), .C(_13_), .Y(w_C_6_) );
NOR2X1 NOR2X1_5 ( .A(_7_), .B(_8_), .Y(_14_) );
INVX1 INVX1_9 ( .A(_14_), .Y(_15_) );
AND2X2 AND2X2_2 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_16_) );
INVX1 INVX1_10 ( .A(_16_), .Y(_17_) );
NAND3X1 NAND3X1_4 ( .A(_15_), .B(_17_), .C(_13_), .Y(_18_) );
OAI21X1 OAI21X1_4 ( .A(i_add2[6]), .B(i_add1[6]), .C(_18_), .Y(_19_) );
INVX1 INVX1_11 ( .A(_19_), .Y(w_C_7_) );
INVX1 INVX1_12 ( .A(i_add2[7]), .Y(_20_) );
INVX1 INVX1_13 ( .A(i_add1[7]), .Y(_21_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_14 ( .A(_22_), .Y(_23_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_24_) );
INVX1 INVX1_15 ( .A(_24_), .Y(_25_) );
NAND3X1 NAND3X1_5 ( .A(_23_), .B(_25_), .C(_18_), .Y(_26_) );
OAI21X1 OAI21X1_5 ( .A(_20_), .B(_21_), .C(_26_), .Y(w_C_8_) );
NOR2X1 NOR2X1_8 ( .A(_20_), .B(_21_), .Y(_27_) );
INVX1 INVX1_16 ( .A(_27_), .Y(_28_) );
AND2X2 AND2X2_3 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_29_) );
INVX1 INVX1_17 ( .A(_29_), .Y(_30_) );
NAND3X1 NAND3X1_6 ( .A(_28_), .B(_30_), .C(_26_), .Y(_31_) );
OAI21X1 OAI21X1_6 ( .A(i_add2[8]), .B(i_add1[8]), .C(_31_), .Y(_32_) );
INVX1 INVX1_18 ( .A(_32_), .Y(w_C_9_) );
INVX1 INVX1_19 ( .A(i_add2[9]), .Y(_33_) );
INVX1 INVX1_20 ( .A(i_add1[9]), .Y(_34_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_35_) );
INVX1 INVX1_21 ( .A(_35_), .Y(_36_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_37_) );
INVX1 INVX1_22 ( .A(_37_), .Y(_38_) );
NAND3X1 NAND3X1_7 ( .A(_36_), .B(_38_), .C(_31_), .Y(_39_) );
OAI21X1 OAI21X1_7 ( .A(_33_), .B(_34_), .C(_39_), .Y(w_C_10_) );
NOR2X1 NOR2X1_11 ( .A(_33_), .B(_34_), .Y(_40_) );
INVX1 INVX1_23 ( .A(_40_), .Y(_41_) );
AND2X2 AND2X2_4 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_42_) );
INVX1 INVX1_24 ( .A(_42_), .Y(_43_) );
NAND3X1 NAND3X1_8 ( .A(_41_), .B(_43_), .C(_39_), .Y(_44_) );
OAI21X1 OAI21X1_8 ( .A(i_add2[10]), .B(i_add1[10]), .C(_44_), .Y(_45_) );
INVX1 INVX1_25 ( .A(_45_), .Y(w_C_11_) );
INVX1 INVX1_26 ( .A(i_add2[11]), .Y(_46_) );
INVX1 INVX1_27 ( .A(i_add1[11]), .Y(_47_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_48_) );
INVX1 INVX1_28 ( .A(_48_), .Y(_49_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_50_) );
INVX1 INVX1_29 ( .A(_50_), .Y(_51_) );
NAND3X1 NAND3X1_9 ( .A(_49_), .B(_51_), .C(_44_), .Y(_52_) );
OAI21X1 OAI21X1_9 ( .A(_46_), .B(_47_), .C(_52_), .Y(w_C_12_) );
NOR2X1 NOR2X1_14 ( .A(_46_), .B(_47_), .Y(_53_) );
INVX1 INVX1_30 ( .A(_53_), .Y(_54_) );
AND2X2 AND2X2_5 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_55_) );
INVX1 INVX1_31 ( .A(_55_), .Y(_56_) );
NAND3X1 NAND3X1_10 ( .A(_54_), .B(_56_), .C(_52_), .Y(_57_) );
OAI21X1 OAI21X1_10 ( .A(i_add2[12]), .B(i_add1[12]), .C(_57_), .Y(_58_) );
INVX1 INVX1_32 ( .A(_58_), .Y(w_C_13_) );
INVX1 INVX1_33 ( .A(i_add2[13]), .Y(_59_) );
INVX1 INVX1_34 ( .A(i_add1[13]), .Y(_60_) );
NOR2X1 NOR2X1_15 ( .A(_59_), .B(_60_), .Y(_61_) );
INVX1 INVX1_35 ( .A(_61_), .Y(_62_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_63_) );
INVX1 INVX1_36 ( .A(_63_), .Y(_64_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_65_) );
INVX1 INVX1_37 ( .A(_65_), .Y(_66_) );
NAND3X1 NAND3X1_11 ( .A(_64_), .B(_66_), .C(_57_), .Y(_67_) );
AND2X2 AND2X2_6 ( .A(_67_), .B(_62_), .Y(_68_) );
INVX1 INVX1_38 ( .A(_68_), .Y(w_C_14_) );
AND2X2 AND2X2_7 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_69_) );
INVX1 INVX1_39 ( .A(_69_), .Y(_70_) );
NAND3X1 NAND3X1_12 ( .A(_62_), .B(_70_), .C(_67_), .Y(_71_) );
OAI21X1 OAI21X1_11 ( .A(i_add2[14]), .B(i_add1[14]), .C(_71_), .Y(_72_) );
INVX1 INVX1_40 ( .A(_72_), .Y(w_C_15_) );
INVX1 INVX1_41 ( .A(i_add2[15]), .Y(_73_) );
INVX1 INVX1_42 ( .A(i_add1[15]), .Y(_74_) );
NOR2X1 NOR2X1_18 ( .A(_73_), .B(_74_), .Y(_75_) );
INVX1 INVX1_43 ( .A(_75_), .Y(_76_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_77_) );
INVX1 INVX1_44 ( .A(_77_), .Y(_78_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_79_) );
INVX1 INVX1_45 ( .A(_79_), .Y(_80_) );
NAND3X1 NAND3X1_13 ( .A(_78_), .B(_80_), .C(_71_), .Y(_81_) );
AND2X2 AND2X2_8 ( .A(_81_), .B(_76_), .Y(_82_) );
INVX1 INVX1_46 ( .A(_82_), .Y(w_C_16_) );
AND2X2 AND2X2_9 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_83_) );
INVX1 INVX1_47 ( .A(_83_), .Y(_84_) );
NAND3X1 NAND3X1_14 ( .A(_76_), .B(_84_), .C(_81_), .Y(_85_) );
OAI21X1 OAI21X1_12 ( .A(i_add2[16]), .B(i_add1[16]), .C(_85_), .Y(_86_) );
INVX1 INVX1_48 ( .A(_86_), .Y(w_C_17_) );
INVX1 INVX1_49 ( .A(i_add2[17]), .Y(_87_) );
INVX1 INVX1_50 ( .A(i_add1[17]), .Y(_88_) );
NOR2X1 NOR2X1_21 ( .A(_87_), .B(_88_), .Y(_89_) );
INVX1 INVX1_51 ( .A(_89_), .Y(_90_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_91_) );
INVX1 INVX1_52 ( .A(_91_), .Y(_92_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_93_) );
INVX1 INVX1_53 ( .A(_93_), .Y(_94_) );
NAND3X1 NAND3X1_15 ( .A(_92_), .B(_94_), .C(_85_), .Y(_95_) );
AND2X2 AND2X2_10 ( .A(_95_), .B(_90_), .Y(_96_) );
INVX1 INVX1_54 ( .A(_96_), .Y(w_C_18_) );
AND2X2 AND2X2_11 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_97_) );
INVX1 INVX1_55 ( .A(_97_), .Y(_98_) );
NAND3X1 NAND3X1_16 ( .A(_90_), .B(_98_), .C(_95_), .Y(_99_) );
OAI21X1 OAI21X1_13 ( .A(i_add2[18]), .B(i_add1[18]), .C(_99_), .Y(_100_) );
INVX1 INVX1_56 ( .A(_100_), .Y(w_C_19_) );
INVX1 INVX1_57 ( .A(i_add2[19]), .Y(_101_) );
INVX1 INVX1_58 ( .A(i_add1[19]), .Y(_102_) );
NOR2X1 NOR2X1_24 ( .A(_101_), .B(_102_), .Y(_103_) );
INVX1 INVX1_59 ( .A(_103_), .Y(_104_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_105_) );
INVX1 INVX1_60 ( .A(_105_), .Y(_106_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_107_) );
INVX1 INVX1_61 ( .A(_107_), .Y(_108_) );
NAND3X1 NAND3X1_17 ( .A(_106_), .B(_108_), .C(_99_), .Y(_109_) );
AND2X2 AND2X2_12 ( .A(_109_), .B(_104_), .Y(_110_) );
INVX1 INVX1_62 ( .A(_110_), .Y(w_C_20_) );
AND2X2 AND2X2_13 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_111_) );
INVX1 INVX1_63 ( .A(_111_), .Y(_112_) );
NAND3X1 NAND3X1_18 ( .A(_104_), .B(_112_), .C(_109_), .Y(_113_) );
OAI21X1 OAI21X1_14 ( .A(i_add2[20]), .B(i_add1[20]), .C(_113_), .Y(_114_) );
INVX1 INVX1_64 ( .A(_114_), .Y(w_C_21_) );
INVX1 INVX1_65 ( .A(i_add2[21]), .Y(_115_) );
INVX1 INVX1_66 ( .A(i_add1[21]), .Y(_116_) );
NOR2X1 NOR2X1_27 ( .A(_115_), .B(_116_), .Y(_117_) );
INVX1 INVX1_67 ( .A(_117_), .Y(_118_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_119_) );
INVX1 INVX1_68 ( .A(_119_), .Y(_120_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_121_) );
INVX1 INVX1_69 ( .A(_121_), .Y(_122_) );
NAND3X1 NAND3X1_19 ( .A(_120_), .B(_122_), .C(_113_), .Y(_123_) );
AND2X2 AND2X2_14 ( .A(_123_), .B(_118_), .Y(_124_) );
INVX1 INVX1_70 ( .A(_124_), .Y(w_C_22_) );
AND2X2 AND2X2_15 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_125_) );
INVX1 INVX1_71 ( .A(_125_), .Y(_126_) );
NAND3X1 NAND3X1_20 ( .A(_118_), .B(_126_), .C(_123_), .Y(_127_) );
OAI21X1 OAI21X1_15 ( .A(i_add2[22]), .B(i_add1[22]), .C(_127_), .Y(_128_) );
INVX1 INVX1_72 ( .A(_128_), .Y(w_C_23_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_129_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_130_) );
OAI21X1 OAI21X1_16 ( .A(_130_), .B(_128_), .C(_129_), .Y(w_C_24_) );
OR2X2 OR2X2_2 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_131_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_132_) );
INVX1 INVX1_73 ( .A(_132_), .Y(_133_) );
INVX1 INVX1_74 ( .A(_130_), .Y(_134_) );
NAND3X1 NAND3X1_21 ( .A(_133_), .B(_134_), .C(_127_), .Y(_135_) );
NAND2X1 NAND2X1_8 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_136_) );
NAND3X1 NAND3X1_22 ( .A(_129_), .B(_136_), .C(_135_), .Y(_137_) );
AND2X2 AND2X2_16 ( .A(_137_), .B(_131_), .Y(w_C_25_) );
INVX1 INVX1_75 ( .A(i_add2[25]), .Y(_138_) );
INVX1 INVX1_76 ( .A(i_add1[25]), .Y(_139_) );
NAND2X1 NAND2X1_9 ( .A(_138_), .B(_139_), .Y(_140_) );
NAND3X1 NAND3X1_23 ( .A(_131_), .B(_140_), .C(_137_), .Y(_141_) );
OAI21X1 OAI21X1_17 ( .A(_138_), .B(_139_), .C(_141_), .Y(w_C_26_) );
INVX1 INVX1_77 ( .A(i_add2[26]), .Y(_142_) );
INVX1 INVX1_78 ( .A(i_add1[26]), .Y(_143_) );
NAND2X1 NAND2X1_10 ( .A(_142_), .B(_143_), .Y(_144_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_145_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_146_) );
NAND3X1 NAND3X1_24 ( .A(_145_), .B(_146_), .C(_141_), .Y(_147_) );
AND2X2 AND2X2_17 ( .A(_147_), .B(_144_), .Y(w_C_27_) );
INVX1 INVX1_79 ( .A(i_add2[27]), .Y(_148_) );
INVX1 INVX1_80 ( .A(i_add1[27]), .Y(_149_) );
NAND2X1 NAND2X1_13 ( .A(_148_), .B(_149_), .Y(_150_) );
NAND3X1 NAND3X1_25 ( .A(_144_), .B(_150_), .C(_147_), .Y(_151_) );
OAI21X1 OAI21X1_18 ( .A(_148_), .B(_149_), .C(_151_), .Y(w_C_28_) );
OR2X2 OR2X2_3 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_152_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_153_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_154_) );
NAND3X1 NAND3X1_26 ( .A(_153_), .B(_154_), .C(_151_), .Y(_155_) );
AND2X2 AND2X2_18 ( .A(_155_), .B(_152_), .Y(w_C_29_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_156_) );
OR2X2 OR2X2_4 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_157_) );
NAND3X1 NAND3X1_27 ( .A(_152_), .B(_157_), .C(_155_), .Y(_158_) );
NAND2X1 NAND2X1_17 ( .A(_156_), .B(_158_), .Y(w_C_30_) );
BUFX2 BUFX2_1 ( .A(_166__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_166__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_166__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_166__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_166__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_166__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_166__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_166__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_166__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_166__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_166__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_166__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_166__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_166__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_166__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_166__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_166__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_166__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_166__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_166__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_166__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_166__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_166__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_166__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_166__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_166__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_166__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_166__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_166__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_166__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(w_C_30_), .Y(o_result[30]) );
INVX1 INVX1_81 ( .A(w_C_4_), .Y(_170_) );
OR2X2 OR2X2_5 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_171_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_172_) );
NAND3X1 NAND3X1_28 ( .A(_170_), .B(_172_), .C(_171_), .Y(_173_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_167_) );
AND2X2 AND2X2_19 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_168_) );
OAI21X1 OAI21X1_19 ( .A(_167_), .B(_168_), .C(w_C_4_), .Y(_169_) );
NAND2X1 NAND2X1_19 ( .A(_169_), .B(_173_), .Y(_166__4_) );
INVX1 INVX1_82 ( .A(w_C_5_), .Y(_177_) );
OR2X2 OR2X2_6 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_178_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_179_) );
NAND3X1 NAND3X1_29 ( .A(_177_), .B(_179_), .C(_178_), .Y(_180_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_174_) );
AND2X2 AND2X2_20 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_175_) );
OAI21X1 OAI21X1_20 ( .A(_174_), .B(_175_), .C(w_C_5_), .Y(_176_) );
NAND2X1 NAND2X1_21 ( .A(_176_), .B(_180_), .Y(_166__5_) );
INVX1 INVX1_83 ( .A(w_C_6_), .Y(_184_) );
OR2X2 OR2X2_7 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_185_) );
NAND2X1 NAND2X1_22 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_186_) );
NAND3X1 NAND3X1_30 ( .A(_184_), .B(_186_), .C(_185_), .Y(_187_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_181_) );
AND2X2 AND2X2_21 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_182_) );
OAI21X1 OAI21X1_21 ( .A(_181_), .B(_182_), .C(w_C_6_), .Y(_183_) );
NAND2X1 NAND2X1_23 ( .A(_183_), .B(_187_), .Y(_166__6_) );
INVX1 INVX1_84 ( .A(w_C_7_), .Y(_191_) );
OR2X2 OR2X2_8 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_192_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_193_) );
NAND3X1 NAND3X1_31 ( .A(_191_), .B(_193_), .C(_192_), .Y(_194_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_188_) );
AND2X2 AND2X2_22 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_189_) );
OAI21X1 OAI21X1_22 ( .A(_188_), .B(_189_), .C(w_C_7_), .Y(_190_) );
NAND2X1 NAND2X1_25 ( .A(_190_), .B(_194_), .Y(_166__7_) );
INVX1 INVX1_85 ( .A(w_C_8_), .Y(_198_) );
OR2X2 OR2X2_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_199_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_200_) );
NAND3X1 NAND3X1_32 ( .A(_198_), .B(_200_), .C(_199_), .Y(_201_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_195_) );
AND2X2 AND2X2_23 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_196_) );
OAI21X1 OAI21X1_23 ( .A(_195_), .B(_196_), .C(w_C_8_), .Y(_197_) );
NAND2X1 NAND2X1_27 ( .A(_197_), .B(_201_), .Y(_166__8_) );
INVX1 INVX1_86 ( .A(w_C_9_), .Y(_205_) );
OR2X2 OR2X2_10 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_206_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_207_) );
NAND3X1 NAND3X1_33 ( .A(_205_), .B(_207_), .C(_206_), .Y(_208_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_202_) );
AND2X2 AND2X2_24 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_203_) );
OAI21X1 OAI21X1_24 ( .A(_202_), .B(_203_), .C(w_C_9_), .Y(_204_) );
NAND2X1 NAND2X1_29 ( .A(_204_), .B(_208_), .Y(_166__9_) );
INVX1 INVX1_87 ( .A(w_C_10_), .Y(_212_) );
OR2X2 OR2X2_11 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_213_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_214_) );
NAND3X1 NAND3X1_34 ( .A(_212_), .B(_214_), .C(_213_), .Y(_215_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_209_) );
AND2X2 AND2X2_25 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_210_) );
OAI21X1 OAI21X1_25 ( .A(_209_), .B(_210_), .C(w_C_10_), .Y(_211_) );
NAND2X1 NAND2X1_31 ( .A(_211_), .B(_215_), .Y(_166__10_) );
INVX1 INVX1_88 ( .A(w_C_11_), .Y(_219_) );
OR2X2 OR2X2_12 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_220_) );
NAND2X1 NAND2X1_32 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_221_) );
NAND3X1 NAND3X1_35 ( .A(_219_), .B(_221_), .C(_220_), .Y(_222_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_216_) );
AND2X2 AND2X2_26 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_217_) );
OAI21X1 OAI21X1_26 ( .A(_216_), .B(_217_), .C(w_C_11_), .Y(_218_) );
NAND2X1 NAND2X1_33 ( .A(_218_), .B(_222_), .Y(_166__11_) );
INVX1 INVX1_89 ( .A(w_C_12_), .Y(_226_) );
OR2X2 OR2X2_13 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_227_) );
NAND2X1 NAND2X1_34 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_228_) );
NAND3X1 NAND3X1_36 ( .A(_226_), .B(_228_), .C(_227_), .Y(_229_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_223_) );
AND2X2 AND2X2_27 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_224_) );
OAI21X1 OAI21X1_27 ( .A(_223_), .B(_224_), .C(w_C_12_), .Y(_225_) );
NAND2X1 NAND2X1_35 ( .A(_225_), .B(_229_), .Y(_166__12_) );
INVX1 INVX1_90 ( .A(w_C_13_), .Y(_233_) );
OR2X2 OR2X2_14 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_234_) );
NAND2X1 NAND2X1_36 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_235_) );
NAND3X1 NAND3X1_37 ( .A(_233_), .B(_235_), .C(_234_), .Y(_236_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_230_) );
AND2X2 AND2X2_28 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_231_) );
OAI21X1 OAI21X1_28 ( .A(_230_), .B(_231_), .C(w_C_13_), .Y(_232_) );
NAND2X1 NAND2X1_37 ( .A(_232_), .B(_236_), .Y(_166__13_) );
INVX1 INVX1_91 ( .A(w_C_14_), .Y(_240_) );
OR2X2 OR2X2_15 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_241_) );
NAND2X1 NAND2X1_38 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_242_) );
NAND3X1 NAND3X1_38 ( .A(_240_), .B(_242_), .C(_241_), .Y(_243_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_237_) );
AND2X2 AND2X2_29 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_238_) );
OAI21X1 OAI21X1_29 ( .A(_237_), .B(_238_), .C(w_C_14_), .Y(_239_) );
NAND2X1 NAND2X1_39 ( .A(_239_), .B(_243_), .Y(_166__14_) );
INVX1 INVX1_92 ( .A(w_C_15_), .Y(_247_) );
OR2X2 OR2X2_16 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_248_) );
NAND2X1 NAND2X1_40 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_249_) );
NAND3X1 NAND3X1_39 ( .A(_247_), .B(_249_), .C(_248_), .Y(_250_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_244_) );
AND2X2 AND2X2_30 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_245_) );
OAI21X1 OAI21X1_30 ( .A(_244_), .B(_245_), .C(w_C_15_), .Y(_246_) );
NAND2X1 NAND2X1_41 ( .A(_246_), .B(_250_), .Y(_166__15_) );
INVX1 INVX1_93 ( .A(w_C_16_), .Y(_254_) );
OR2X2 OR2X2_17 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_255_) );
NAND2X1 NAND2X1_42 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_256_) );
NAND3X1 NAND3X1_40 ( .A(_254_), .B(_256_), .C(_255_), .Y(_257_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_251_) );
AND2X2 AND2X2_31 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_252_) );
OAI21X1 OAI21X1_31 ( .A(_251_), .B(_252_), .C(w_C_16_), .Y(_253_) );
NAND2X1 NAND2X1_43 ( .A(_253_), .B(_257_), .Y(_166__16_) );
INVX1 INVX1_94 ( .A(w_C_17_), .Y(_261_) );
OR2X2 OR2X2_18 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_262_) );
NAND2X1 NAND2X1_44 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_263_) );
NAND3X1 NAND3X1_41 ( .A(_261_), .B(_263_), .C(_262_), .Y(_264_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_258_) );
AND2X2 AND2X2_32 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_259_) );
OAI21X1 OAI21X1_32 ( .A(_258_), .B(_259_), .C(w_C_17_), .Y(_260_) );
NAND2X1 NAND2X1_45 ( .A(_260_), .B(_264_), .Y(_166__17_) );
INVX1 INVX1_95 ( .A(w_C_18_), .Y(_268_) );
OR2X2 OR2X2_19 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_269_) );
NAND2X1 NAND2X1_46 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_270_) );
NAND3X1 NAND3X1_42 ( .A(_268_), .B(_270_), .C(_269_), .Y(_271_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_265_) );
AND2X2 AND2X2_33 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_266_) );
OAI21X1 OAI21X1_33 ( .A(_265_), .B(_266_), .C(w_C_18_), .Y(_267_) );
NAND2X1 NAND2X1_47 ( .A(_267_), .B(_271_), .Y(_166__18_) );
INVX1 INVX1_96 ( .A(w_C_19_), .Y(_275_) );
OR2X2 OR2X2_20 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_276_) );
NAND2X1 NAND2X1_48 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_277_) );
NAND3X1 NAND3X1_43 ( .A(_275_), .B(_277_), .C(_276_), .Y(_278_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_272_) );
AND2X2 AND2X2_34 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_273_) );
OAI21X1 OAI21X1_34 ( .A(_272_), .B(_273_), .C(w_C_19_), .Y(_274_) );
NAND2X1 NAND2X1_49 ( .A(_274_), .B(_278_), .Y(_166__19_) );
INVX1 INVX1_97 ( .A(w_C_20_), .Y(_282_) );
OR2X2 OR2X2_21 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_283_) );
NAND2X1 NAND2X1_50 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_284_) );
NAND3X1 NAND3X1_44 ( .A(_282_), .B(_284_), .C(_283_), .Y(_285_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_279_) );
AND2X2 AND2X2_35 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_280_) );
OAI21X1 OAI21X1_35 ( .A(_279_), .B(_280_), .C(w_C_20_), .Y(_281_) );
NAND2X1 NAND2X1_51 ( .A(_281_), .B(_285_), .Y(_166__20_) );
INVX1 INVX1_98 ( .A(w_C_21_), .Y(_289_) );
OR2X2 OR2X2_22 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_290_) );
NAND2X1 NAND2X1_52 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_291_) );
NAND3X1 NAND3X1_45 ( .A(_289_), .B(_291_), .C(_290_), .Y(_292_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_286_) );
AND2X2 AND2X2_36 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_287_) );
OAI21X1 OAI21X1_36 ( .A(_286_), .B(_287_), .C(w_C_21_), .Y(_288_) );
NAND2X1 NAND2X1_53 ( .A(_288_), .B(_292_), .Y(_166__21_) );
INVX1 INVX1_99 ( .A(w_C_22_), .Y(_296_) );
OR2X2 OR2X2_23 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_297_) );
NAND2X1 NAND2X1_54 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_298_) );
NAND3X1 NAND3X1_46 ( .A(_296_), .B(_298_), .C(_297_), .Y(_299_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_293_) );
AND2X2 AND2X2_37 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_294_) );
OAI21X1 OAI21X1_37 ( .A(_293_), .B(_294_), .C(w_C_22_), .Y(_295_) );
NAND2X1 NAND2X1_55 ( .A(_295_), .B(_299_), .Y(_166__22_) );
INVX1 INVX1_100 ( .A(w_C_23_), .Y(_303_) );
OR2X2 OR2X2_24 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_304_) );
NAND2X1 NAND2X1_56 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_305_) );
NAND3X1 NAND3X1_47 ( .A(_303_), .B(_305_), .C(_304_), .Y(_306_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_300_) );
AND2X2 AND2X2_38 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_301_) );
OAI21X1 OAI21X1_38 ( .A(_300_), .B(_301_), .C(w_C_23_), .Y(_302_) );
NAND2X1 NAND2X1_57 ( .A(_302_), .B(_306_), .Y(_166__23_) );
INVX1 INVX1_101 ( .A(w_C_24_), .Y(_310_) );
OR2X2 OR2X2_25 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_311_) );
NAND2X1 NAND2X1_58 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_312_) );
NAND3X1 NAND3X1_48 ( .A(_310_), .B(_312_), .C(_311_), .Y(_313_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_307_) );
AND2X2 AND2X2_39 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_308_) );
OAI21X1 OAI21X1_39 ( .A(_307_), .B(_308_), .C(w_C_24_), .Y(_309_) );
NAND2X1 NAND2X1_59 ( .A(_309_), .B(_313_), .Y(_166__24_) );
INVX1 INVX1_102 ( .A(w_C_25_), .Y(_317_) );
OR2X2 OR2X2_26 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_318_) );
NAND2X1 NAND2X1_60 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_319_) );
NAND3X1 NAND3X1_49 ( .A(_317_), .B(_319_), .C(_318_), .Y(_320_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_314_) );
AND2X2 AND2X2_40 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_315_) );
OAI21X1 OAI21X1_40 ( .A(_314_), .B(_315_), .C(w_C_25_), .Y(_316_) );
NAND2X1 NAND2X1_61 ( .A(_316_), .B(_320_), .Y(_166__25_) );
INVX1 INVX1_103 ( .A(w_C_26_), .Y(_324_) );
OR2X2 OR2X2_27 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_325_) );
NAND2X1 NAND2X1_62 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_326_) );
NAND3X1 NAND3X1_50 ( .A(_324_), .B(_326_), .C(_325_), .Y(_327_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_321_) );
AND2X2 AND2X2_41 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_322_) );
OAI21X1 OAI21X1_41 ( .A(_321_), .B(_322_), .C(w_C_26_), .Y(_323_) );
NAND2X1 NAND2X1_63 ( .A(_323_), .B(_327_), .Y(_166__26_) );
INVX1 INVX1_104 ( .A(w_C_27_), .Y(_331_) );
OR2X2 OR2X2_28 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_332_) );
NAND2X1 NAND2X1_64 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_333_) );
NAND3X1 NAND3X1_51 ( .A(_331_), .B(_333_), .C(_332_), .Y(_334_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_328_) );
AND2X2 AND2X2_42 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_329_) );
OAI21X1 OAI21X1_42 ( .A(_328_), .B(_329_), .C(w_C_27_), .Y(_330_) );
NAND2X1 NAND2X1_65 ( .A(_330_), .B(_334_), .Y(_166__27_) );
INVX1 INVX1_105 ( .A(w_C_28_), .Y(_338_) );
OR2X2 OR2X2_29 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_339_) );
NAND2X1 NAND2X1_66 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_340_) );
NAND3X1 NAND3X1_52 ( .A(_338_), .B(_340_), .C(_339_), .Y(_341_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_335_) );
AND2X2 AND2X2_43 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_336_) );
OAI21X1 OAI21X1_43 ( .A(_335_), .B(_336_), .C(w_C_28_), .Y(_337_) );
NAND2X1 NAND2X1_67 ( .A(_337_), .B(_341_), .Y(_166__28_) );
INVX1 INVX1_106 ( .A(w_C_29_), .Y(_345_) );
OR2X2 OR2X2_30 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_346_) );
NAND2X1 NAND2X1_68 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_347_) );
NAND3X1 NAND3X1_53 ( .A(_345_), .B(_347_), .C(_346_), .Y(_348_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_342_) );
AND2X2 AND2X2_44 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_343_) );
OAI21X1 OAI21X1_44 ( .A(_342_), .B(_343_), .C(w_C_29_), .Y(_344_) );
NAND2X1 NAND2X1_69 ( .A(_344_), .B(_348_), .Y(_166__29_) );
INVX1 INVX1_107 ( .A(gnd), .Y(_352_) );
OR2X2 OR2X2_31 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_353_) );
NAND2X1 NAND2X1_70 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_354_) );
NAND3X1 NAND3X1_54 ( .A(_352_), .B(_354_), .C(_353_), .Y(_355_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_349_) );
AND2X2 AND2X2_45 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_350_) );
OAI21X1 OAI21X1_45 ( .A(_349_), .B(_350_), .C(gnd), .Y(_351_) );
NAND2X1 NAND2X1_71 ( .A(_351_), .B(_355_), .Y(_166__0_) );
INVX1 INVX1_108 ( .A(w_C_1_), .Y(_359_) );
OR2X2 OR2X2_32 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_360_) );
NAND2X1 NAND2X1_72 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_361_) );
NAND3X1 NAND3X1_55 ( .A(_359_), .B(_361_), .C(_360_), .Y(_362_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_356_) );
AND2X2 AND2X2_46 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_357_) );
OAI21X1 OAI21X1_46 ( .A(_356_), .B(_357_), .C(w_C_1_), .Y(_358_) );
NAND2X1 NAND2X1_73 ( .A(_358_), .B(_362_), .Y(_166__1_) );
INVX1 INVX1_109 ( .A(w_C_2_), .Y(_366_) );
OR2X2 OR2X2_33 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_367_) );
NAND2X1 NAND2X1_74 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_368_) );
NAND3X1 NAND3X1_56 ( .A(_366_), .B(_368_), .C(_367_), .Y(_369_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_363_) );
AND2X2 AND2X2_47 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_364_) );
OAI21X1 OAI21X1_47 ( .A(_363_), .B(_364_), .C(w_C_2_), .Y(_365_) );
NAND2X1 NAND2X1_75 ( .A(_365_), .B(_369_), .Y(_166__2_) );
INVX1 INVX1_110 ( .A(w_C_3_), .Y(_373_) );
OR2X2 OR2X2_34 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_374_) );
NAND2X1 NAND2X1_76 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_375_) );
NAND3X1 NAND3X1_57 ( .A(_373_), .B(_375_), .C(_374_), .Y(_376_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_370_) );
AND2X2 AND2X2_48 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_371_) );
OAI21X1 OAI21X1_48 ( .A(_370_), .B(_371_), .C(w_C_3_), .Y(_372_) );
NAND2X1 NAND2X1_77 ( .A(_372_), .B(_376_), .Y(_166__3_) );
BUFX2 BUFX2_32 ( .A(w_C_30_), .Y(_166__30_) );
BUFX2 BUFX2_33 ( .A(gnd), .Y(w_C_0_) );
endmodule
