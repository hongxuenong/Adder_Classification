module cla_13bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];

NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_4_) );
INVX1 INVX1_1 ( .A(_4_), .Y(w_C_1_) );
NAND2X1 NAND2X1_2 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
NAND2X1 NAND2X1_3 ( .A(_4_), .B(_5_), .Y(_6_) );
OAI21X1 OAI21X1_1 ( .A(i_add2[1]), .B(i_add1[1]), .C(_6_), .Y(_7_) );
INVX1 INVX1_2 ( .A(_7_), .Y(w_C_2_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_8_) );
OR2X2 OR2X2_1 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_9_) );
OR2X2 OR2X2_2 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_10_) );
NAND3X1 NAND3X1_1 ( .A(_9_), .B(_10_), .C(_6_), .Y(_11_) );
NAND2X1 NAND2X1_5 ( .A(_8_), .B(_11_), .Y(w_C_3_) );
OR2X2 OR2X2_3 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_12_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_13_) );
NAND3X1 NAND3X1_2 ( .A(_8_), .B(_13_), .C(_11_), .Y(_14_) );
AND2X2 AND2X2_1 ( .A(_14_), .B(_12_), .Y(w_C_4_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_15_) );
OR2X2 OR2X2_4 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_16_) );
NAND3X1 NAND3X1_3 ( .A(_12_), .B(_16_), .C(_14_), .Y(_17_) );
NAND2X1 NAND2X1_8 ( .A(_15_), .B(_17_), .Y(w_C_5_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_18_) );
INVX1 INVX1_3 ( .A(_18_), .Y(_19_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_20_) );
NAND3X1 NAND3X1_4 ( .A(_15_), .B(_20_), .C(_17_), .Y(_21_) );
AND2X2 AND2X2_2 ( .A(_21_), .B(_19_), .Y(w_C_6_) );
INVX1 INVX1_4 ( .A(i_add2[6]), .Y(_22_) );
INVX1 INVX1_5 ( .A(i_add1[6]), .Y(_23_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_24_) );
INVX1 INVX1_6 ( .A(_24_), .Y(_25_) );
NAND3X1 NAND3X1_5 ( .A(_19_), .B(_25_), .C(_21_), .Y(_26_) );
OAI21X1 OAI21X1_2 ( .A(_22_), .B(_23_), .C(_26_), .Y(w_C_7_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_27_) );
INVX1 INVX1_7 ( .A(_27_), .Y(_28_) );
NOR2X1 NOR2X1_4 ( .A(_22_), .B(_23_), .Y(_29_) );
INVX1 INVX1_8 ( .A(_29_), .Y(_30_) );
AND2X2 AND2X2_3 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_31_) );
INVX1 INVX1_9 ( .A(_31_), .Y(_32_) );
NAND3X1 NAND3X1_6 ( .A(_30_), .B(_32_), .C(_26_), .Y(_33_) );
AND2X2 AND2X2_4 ( .A(_33_), .B(_28_), .Y(w_C_8_) );
INVX1 INVX1_10 ( .A(i_add2[8]), .Y(_34_) );
INVX1 INVX1_11 ( .A(i_add1[8]), .Y(_35_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_36_) );
INVX1 INVX1_12 ( .A(_36_), .Y(_37_) );
NAND3X1 NAND3X1_7 ( .A(_28_), .B(_37_), .C(_33_), .Y(_38_) );
OAI21X1 OAI21X1_3 ( .A(_34_), .B(_35_), .C(_38_), .Y(w_C_9_) );
NOR2X1 NOR2X1_6 ( .A(_34_), .B(_35_), .Y(_39_) );
INVX1 INVX1_13 ( .A(_39_), .Y(_40_) );
AND2X2 AND2X2_5 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_41_) );
INVX1 INVX1_14 ( .A(_41_), .Y(_42_) );
NAND3X1 NAND3X1_8 ( .A(_40_), .B(_42_), .C(_38_), .Y(_43_) );
OAI21X1 OAI21X1_4 ( .A(i_add2[9]), .B(i_add1[9]), .C(_43_), .Y(_44_) );
INVX1 INVX1_15 ( .A(_44_), .Y(w_C_10_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_45_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_46_) );
OAI21X1 OAI21X1_5 ( .A(_46_), .B(_44_), .C(_45_), .Y(w_C_11_) );
OR2X2 OR2X2_5 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_47_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_48_) );
INVX1 INVX1_16 ( .A(_48_), .Y(_49_) );
INVX1 INVX1_17 ( .A(_46_), .Y(_50_) );
NAND3X1 NAND3X1_9 ( .A(_49_), .B(_50_), .C(_43_), .Y(_51_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_52_) );
NAND3X1 NAND3X1_10 ( .A(_45_), .B(_52_), .C(_51_), .Y(_0_) );
AND2X2 AND2X2_6 ( .A(_0_), .B(_47_), .Y(w_C_12_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_1_) );
OR2X2 OR2X2_6 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_2_) );
NAND3X1 NAND3X1_11 ( .A(_47_), .B(_2_), .C(_0_), .Y(_3_) );
NAND2X1 NAND2X1_13 ( .A(_1_), .B(_3_), .Y(w_C_13_) );
BUFX2 BUFX2_1 ( .A(_53__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_53__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_53__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_53__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_53__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_53__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_53__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_53__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_53__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_53__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_53__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_53__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_53__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(w_C_13_), .Y(o_result[13]) );
INVX1 INVX1_18 ( .A(w_C_4_), .Y(_57_) );
OR2X2 OR2X2_7 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_58_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_59_) );
NAND3X1 NAND3X1_12 ( .A(_57_), .B(_59_), .C(_58_), .Y(_60_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_54_) );
AND2X2 AND2X2_7 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_55_) );
OAI21X1 OAI21X1_6 ( .A(_54_), .B(_55_), .C(w_C_4_), .Y(_56_) );
NAND2X1 NAND2X1_15 ( .A(_56_), .B(_60_), .Y(_53__4_) );
INVX1 INVX1_19 ( .A(w_C_5_), .Y(_64_) );
OR2X2 OR2X2_8 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_65_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_66_) );
NAND3X1 NAND3X1_13 ( .A(_64_), .B(_66_), .C(_65_), .Y(_67_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_61_) );
AND2X2 AND2X2_8 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_62_) );
OAI21X1 OAI21X1_7 ( .A(_61_), .B(_62_), .C(w_C_5_), .Y(_63_) );
NAND2X1 NAND2X1_17 ( .A(_63_), .B(_67_), .Y(_53__5_) );
INVX1 INVX1_20 ( .A(w_C_6_), .Y(_71_) );
OR2X2 OR2X2_9 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_72_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_73_) );
NAND3X1 NAND3X1_14 ( .A(_71_), .B(_73_), .C(_72_), .Y(_74_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_68_) );
AND2X2 AND2X2_9 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_69_) );
OAI21X1 OAI21X1_8 ( .A(_68_), .B(_69_), .C(w_C_6_), .Y(_70_) );
NAND2X1 NAND2X1_19 ( .A(_70_), .B(_74_), .Y(_53__6_) );
INVX1 INVX1_21 ( .A(w_C_7_), .Y(_78_) );
OR2X2 OR2X2_10 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_79_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_80_) );
NAND3X1 NAND3X1_15 ( .A(_78_), .B(_80_), .C(_79_), .Y(_81_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_75_) );
AND2X2 AND2X2_10 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_76_) );
OAI21X1 OAI21X1_9 ( .A(_75_), .B(_76_), .C(w_C_7_), .Y(_77_) );
NAND2X1 NAND2X1_21 ( .A(_77_), .B(_81_), .Y(_53__7_) );
INVX1 INVX1_22 ( .A(w_C_8_), .Y(_85_) );
OR2X2 OR2X2_11 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_86_) );
NAND2X1 NAND2X1_22 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_87_) );
NAND3X1 NAND3X1_16 ( .A(_85_), .B(_87_), .C(_86_), .Y(_88_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_82_) );
AND2X2 AND2X2_11 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_83_) );
OAI21X1 OAI21X1_10 ( .A(_82_), .B(_83_), .C(w_C_8_), .Y(_84_) );
NAND2X1 NAND2X1_23 ( .A(_84_), .B(_88_), .Y(_53__8_) );
INVX1 INVX1_23 ( .A(w_C_9_), .Y(_92_) );
OR2X2 OR2X2_12 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_93_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_94_) );
NAND3X1 NAND3X1_17 ( .A(_92_), .B(_94_), .C(_93_), .Y(_95_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_89_) );
AND2X2 AND2X2_12 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_90_) );
OAI21X1 OAI21X1_11 ( .A(_89_), .B(_90_), .C(w_C_9_), .Y(_91_) );
NAND2X1 NAND2X1_25 ( .A(_91_), .B(_95_), .Y(_53__9_) );
INVX1 INVX1_24 ( .A(w_C_10_), .Y(_99_) );
OR2X2 OR2X2_13 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_100_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_101_) );
NAND3X1 NAND3X1_18 ( .A(_99_), .B(_101_), .C(_100_), .Y(_102_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_96_) );
AND2X2 AND2X2_13 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_97_) );
OAI21X1 OAI21X1_12 ( .A(_96_), .B(_97_), .C(w_C_10_), .Y(_98_) );
NAND2X1 NAND2X1_27 ( .A(_98_), .B(_102_), .Y(_53__10_) );
INVX1 INVX1_25 ( .A(w_C_11_), .Y(_106_) );
OR2X2 OR2X2_14 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_107_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_108_) );
NAND3X1 NAND3X1_19 ( .A(_106_), .B(_108_), .C(_107_), .Y(_109_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_103_) );
AND2X2 AND2X2_14 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_104_) );
OAI21X1 OAI21X1_13 ( .A(_103_), .B(_104_), .C(w_C_11_), .Y(_105_) );
NAND2X1 NAND2X1_29 ( .A(_105_), .B(_109_), .Y(_53__11_) );
INVX1 INVX1_26 ( .A(w_C_12_), .Y(_113_) );
OR2X2 OR2X2_15 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_114_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_115_) );
NAND3X1 NAND3X1_20 ( .A(_113_), .B(_115_), .C(_114_), .Y(_116_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_110_) );
AND2X2 AND2X2_15 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_111_) );
OAI21X1 OAI21X1_14 ( .A(_110_), .B(_111_), .C(w_C_12_), .Y(_112_) );
NAND2X1 NAND2X1_31 ( .A(_112_), .B(_116_), .Y(_53__12_) );
INVX1 INVX1_27 ( .A(1'b0), .Y(_120_) );
OR2X2 OR2X2_16 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_121_) );
NAND2X1 NAND2X1_32 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_122_) );
NAND3X1 NAND3X1_21 ( .A(_120_), .B(_122_), .C(_121_), .Y(_123_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_117_) );
AND2X2 AND2X2_16 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_118_) );
OAI21X1 OAI21X1_15 ( .A(_117_), .B(_118_), .C(1'b0), .Y(_119_) );
NAND2X1 NAND2X1_33 ( .A(_119_), .B(_123_), .Y(_53__0_) );
INVX1 INVX1_28 ( .A(w_C_1_), .Y(_127_) );
OR2X2 OR2X2_17 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_128_) );
NAND2X1 NAND2X1_34 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_129_) );
NAND3X1 NAND3X1_22 ( .A(_127_), .B(_129_), .C(_128_), .Y(_130_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_124_) );
AND2X2 AND2X2_17 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_125_) );
OAI21X1 OAI21X1_16 ( .A(_124_), .B(_125_), .C(w_C_1_), .Y(_126_) );
NAND2X1 NAND2X1_35 ( .A(_126_), .B(_130_), .Y(_53__1_) );
INVX1 INVX1_29 ( .A(w_C_2_), .Y(_134_) );
OR2X2 OR2X2_18 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_135_) );
NAND2X1 NAND2X1_36 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_136_) );
NAND3X1 NAND3X1_23 ( .A(_134_), .B(_136_), .C(_135_), .Y(_137_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_131_) );
AND2X2 AND2X2_18 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_132_) );
OAI21X1 OAI21X1_17 ( .A(_131_), .B(_132_), .C(w_C_2_), .Y(_133_) );
NAND2X1 NAND2X1_37 ( .A(_133_), .B(_137_), .Y(_53__2_) );
INVX1 INVX1_30 ( .A(w_C_3_), .Y(_141_) );
OR2X2 OR2X2_19 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_142_) );
NAND2X1 NAND2X1_38 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_143_) );
NAND3X1 NAND3X1_24 ( .A(_141_), .B(_143_), .C(_142_), .Y(_144_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_138_) );
AND2X2 AND2X2_19 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_139_) );
OAI21X1 OAI21X1_18 ( .A(_138_), .B(_139_), .C(w_C_3_), .Y(_140_) );
NAND2X1 NAND2X1_39 ( .A(_140_), .B(_144_), .Y(_53__3_) );
BUFX2 BUFX2_15 ( .A(w_C_13_), .Y(_53__13_) );
BUFX2 BUFX2_16 ( .A(1'b0), .Y(w_C_0_) );
endmodule
