module cla_10bit (i_add1, i_add2, o_result);

input [9:0] i_add1;
input [9:0] i_add2;
output [10:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_1 ( .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_2 ( .A(_1_), .B(_2_), .Y(w_C_2_) );
INVX1 INVX1_2 ( .A(i_add2[2]), .Y(_3_) );
INVX1 INVX1_3 ( .A(i_add1[2]), .Y(_4_) );
NAND2X1 NAND2X1_2 ( .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
OAI21X1 OAI21X1_1 ( .A(_1_), .B(_2_), .C(_6_), .Y(_7_) );
AND2X2 AND2X2_1 ( .A(_7_), .B(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
OR2X2 OR2X2_1 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_1 ( .A(_5_), .B(_9_), .C(_7_), .Y(_10_) );
AND2X2 AND2X2_2 ( .A(_10_), .B(_8_), .Y(_11_) );
INVX1 INVX1_4 ( .A(_11_), .Y(w_C_4_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_12_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
OAI21X1 OAI21X1_2 ( .A(_13_), .B(_11_), .C(_12_), .Y(w_C_5_) );
AND2X2 AND2X2_3 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_14_) );
INVX1 INVX1_5 ( .A(_14_), .Y(_15_) );
INVX1 INVX1_6 ( .A(_13_), .Y(_16_) );
NAND3X1 NAND3X1_2 ( .A(_8_), .B(_12_), .C(_10_), .Y(_17_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_18_) );
INVX1 INVX1_7 ( .A(_18_), .Y(_19_) );
NAND3X1 NAND3X1_3 ( .A(_16_), .B(_19_), .C(_17_), .Y(_20_) );
AND2X2 AND2X2_4 ( .A(_20_), .B(_15_), .Y(_21_) );
INVX1 INVX1_8 ( .A(_21_), .Y(w_C_6_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_23_) );
OAI21X1 OAI21X1_3 ( .A(_23_), .B(_21_), .C(_22_), .Y(w_C_7_) );
INVX1 INVX1_9 ( .A(i_add2[7]), .Y(_24_) );
INVX1 INVX1_10 ( .A(i_add1[7]), .Y(_25_) );
INVX1 INVX1_11 ( .A(_23_), .Y(_26_) );
NAND3X1 NAND3X1_4 ( .A(_15_), .B(_22_), .C(_20_), .Y(_27_) );
NAND2X1 NAND2X1_7 ( .A(_24_), .B(_25_), .Y(_28_) );
NAND3X1 NAND3X1_5 ( .A(_26_), .B(_28_), .C(_27_), .Y(_29_) );
OAI21X1 OAI21X1_4 ( .A(_24_), .B(_25_), .C(_29_), .Y(w_C_8_) );
OR2X2 OR2X2_2 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_30_) );
NAND2X1 NAND2X1_8 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_31_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_32_) );
NAND3X1 NAND3X1_6 ( .A(_31_), .B(_32_), .C(_29_), .Y(_33_) );
AND2X2 AND2X2_5 ( .A(_33_), .B(_30_), .Y(w_C_9_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_34_) );
OR2X2 OR2X2_3 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_35_) );
NAND3X1 NAND3X1_7 ( .A(_30_), .B(_35_), .C(_33_), .Y(_36_) );
NAND2X1 NAND2X1_11 ( .A(_34_), .B(_36_), .Y(w_C_10_) );
BUFX2 BUFX2_1 ( .A(_37__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_37__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_37__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_37__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_37__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_37__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_37__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_37__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_37__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_37__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(w_C_10_), .Y(o_result[10]) );
INVX1 INVX1_12 ( .A(w_C_4_), .Y(_41_) );
OR2X2 OR2X2_4 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_42_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_43_) );
NAND3X1 NAND3X1_8 ( .A(_41_), .B(_43_), .C(_42_), .Y(_44_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_38_) );
AND2X2 AND2X2_6 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_39_) );
OAI21X1 OAI21X1_5 ( .A(_38_), .B(_39_), .C(w_C_4_), .Y(_40_) );
NAND2X1 NAND2X1_13 ( .A(_40_), .B(_44_), .Y(_37__4_) );
INVX1 INVX1_13 ( .A(w_C_5_), .Y(_48_) );
OR2X2 OR2X2_5 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_49_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_50_) );
NAND3X1 NAND3X1_9 ( .A(_48_), .B(_50_), .C(_49_), .Y(_51_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_45_) );
AND2X2 AND2X2_7 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_46_) );
OAI21X1 OAI21X1_6 ( .A(_45_), .B(_46_), .C(w_C_5_), .Y(_47_) );
NAND2X1 NAND2X1_15 ( .A(_47_), .B(_51_), .Y(_37__5_) );
INVX1 INVX1_14 ( .A(w_C_6_), .Y(_55_) );
OR2X2 OR2X2_6 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_56_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_57_) );
NAND3X1 NAND3X1_10 ( .A(_55_), .B(_57_), .C(_56_), .Y(_58_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_52_) );
AND2X2 AND2X2_8 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_53_) );
OAI21X1 OAI21X1_7 ( .A(_52_), .B(_53_), .C(w_C_6_), .Y(_54_) );
NAND2X1 NAND2X1_17 ( .A(_54_), .B(_58_), .Y(_37__6_) );
INVX1 INVX1_15 ( .A(w_C_7_), .Y(_62_) );
OR2X2 OR2X2_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_63_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_64_) );
NAND3X1 NAND3X1_11 ( .A(_62_), .B(_64_), .C(_63_), .Y(_65_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_59_) );
AND2X2 AND2X2_9 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_60_) );
OAI21X1 OAI21X1_8 ( .A(_59_), .B(_60_), .C(w_C_7_), .Y(_61_) );
NAND2X1 NAND2X1_19 ( .A(_61_), .B(_65_), .Y(_37__7_) );
INVX1 INVX1_16 ( .A(w_C_8_), .Y(_69_) );
OR2X2 OR2X2_8 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_70_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_71_) );
NAND3X1 NAND3X1_12 ( .A(_69_), .B(_71_), .C(_70_), .Y(_72_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_66_) );
AND2X2 AND2X2_10 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_67_) );
OAI21X1 OAI21X1_9 ( .A(_66_), .B(_67_), .C(w_C_8_), .Y(_68_) );
NAND2X1 NAND2X1_21 ( .A(_68_), .B(_72_), .Y(_37__8_) );
INVX1 INVX1_17 ( .A(w_C_9_), .Y(_76_) );
OR2X2 OR2X2_9 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_77_) );
NAND2X1 NAND2X1_22 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_78_) );
NAND3X1 NAND3X1_13 ( .A(_76_), .B(_78_), .C(_77_), .Y(_79_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_73_) );
AND2X2 AND2X2_11 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_74_) );
OAI21X1 OAI21X1_10 ( .A(_73_), .B(_74_), .C(w_C_9_), .Y(_75_) );
NAND2X1 NAND2X1_23 ( .A(_75_), .B(_79_), .Y(_37__9_) );
INVX1 INVX1_18 ( .A(gnd), .Y(_83_) );
OR2X2 OR2X2_10 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_84_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_85_) );
NAND3X1 NAND3X1_14 ( .A(_83_), .B(_85_), .C(_84_), .Y(_86_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_80_) );
AND2X2 AND2X2_12 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_81_) );
OAI21X1 OAI21X1_11 ( .A(_80_), .B(_81_), .C(gnd), .Y(_82_) );
NAND2X1 NAND2X1_25 ( .A(_82_), .B(_86_), .Y(_37__0_) );
INVX1 INVX1_19 ( .A(w_C_1_), .Y(_90_) );
OR2X2 OR2X2_11 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_91_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_92_) );
NAND3X1 NAND3X1_15 ( .A(_90_), .B(_92_), .C(_91_), .Y(_93_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_87_) );
AND2X2 AND2X2_13 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_88_) );
OAI21X1 OAI21X1_12 ( .A(_87_), .B(_88_), .C(w_C_1_), .Y(_89_) );
NAND2X1 NAND2X1_27 ( .A(_89_), .B(_93_), .Y(_37__1_) );
INVX1 INVX1_20 ( .A(w_C_2_), .Y(_97_) );
OR2X2 OR2X2_12 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_98_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_99_) );
NAND3X1 NAND3X1_16 ( .A(_97_), .B(_99_), .C(_98_), .Y(_100_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_94_) );
AND2X2 AND2X2_14 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_95_) );
OAI21X1 OAI21X1_13 ( .A(_94_), .B(_95_), .C(w_C_2_), .Y(_96_) );
NAND2X1 NAND2X1_29 ( .A(_96_), .B(_100_), .Y(_37__2_) );
INVX1 INVX1_21 ( .A(w_C_3_), .Y(_104_) );
OR2X2 OR2X2_13 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_105_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_106_) );
NAND3X1 NAND3X1_17 ( .A(_104_), .B(_106_), .C(_105_), .Y(_107_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_101_) );
AND2X2 AND2X2_15 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_102_) );
OAI21X1 OAI21X1_14 ( .A(_101_), .B(_102_), .C(w_C_3_), .Y(_103_) );
NAND2X1 NAND2X1_31 ( .A(_103_), .B(_107_), .Y(_37__3_) );
BUFX2 BUFX2_12 ( .A(w_C_10_), .Y(_37__10_) );
BUFX2 BUFX2_13 ( .A(gnd), .Y(w_C_0_) );
endmodule
