module cla_53bit (i_add1, i_add2, o_result);

input [52:0] i_add1;
input [52:0] i_add2;
output [53:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

INVX1 INVX1_1 ( .A(i_add1[18]), .Y(_99_) );
NOR2X1 NOR2X1_1 ( .A(_98_), .B(_99_), .Y(_100_) );
INVX1 INVX1_2 ( .A(_100_), .Y(_101_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_102_) );
INVX1 INVX1_3 ( .A(_102_), .Y(_103_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_104_) );
INVX1 INVX1_4 ( .A(_104_), .Y(_105_) );
NAND3X1 NAND3X1_1 ( .A(_103_), .B(_105_), .C(_96_), .Y(_106_) );
AND2X2 AND2X2_1 ( .A(_106_), .B(_101_), .Y(_107_) );
INVX1 INVX1_5 ( .A(_107_), .Y(w_C_19_) );
AND2X2 AND2X2_2 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_108_) );
INVX1 INVX1_6 ( .A(_108_), .Y(_109_) );
NAND3X1 NAND3X1_2 ( .A(_101_), .B(_109_), .C(_106_), .Y(_110_) );
OAI21X1 OAI21X1_1 ( .A(i_add2[19]), .B(i_add1[19]), .C(_110_), .Y(_111_) );
INVX1 INVX1_7 ( .A(_111_), .Y(w_C_20_) );
INVX1 INVX1_8 ( .A(i_add2[20]), .Y(_112_) );
INVX1 INVX1_9 ( .A(i_add1[20]), .Y(_113_) );
NOR2X1 NOR2X1_4 ( .A(_112_), .B(_113_), .Y(_114_) );
INVX1 INVX1_10 ( .A(_114_), .Y(_115_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_116_) );
INVX1 INVX1_11 ( .A(_116_), .Y(_117_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_118_) );
INVX1 INVX1_12 ( .A(_118_), .Y(_119_) );
NAND3X1 NAND3X1_3 ( .A(_117_), .B(_119_), .C(_110_), .Y(_120_) );
AND2X2 AND2X2_3 ( .A(_120_), .B(_115_), .Y(_121_) );
INVX1 INVX1_13 ( .A(_121_), .Y(w_C_21_) );
AND2X2 AND2X2_4 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_122_) );
INVX1 INVX1_14 ( .A(_122_), .Y(_123_) );
NAND3X1 NAND3X1_4 ( .A(_115_), .B(_123_), .C(_120_), .Y(_124_) );
OAI21X1 OAI21X1_2 ( .A(i_add2[21]), .B(i_add1[21]), .C(_124_), .Y(_125_) );
INVX1 INVX1_15 ( .A(_125_), .Y(w_C_22_) );
INVX1 INVX1_16 ( .A(i_add2[22]), .Y(_126_) );
INVX1 INVX1_17 ( .A(i_add1[22]), .Y(_127_) );
NOR2X1 NOR2X1_7 ( .A(_126_), .B(_127_), .Y(_128_) );
INVX1 INVX1_18 ( .A(_128_), .Y(_129_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_130_) );
INVX1 INVX1_19 ( .A(_130_), .Y(_131_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_132_) );
INVX1 INVX1_20 ( .A(_132_), .Y(_133_) );
NAND3X1 NAND3X1_5 ( .A(_131_), .B(_133_), .C(_124_), .Y(_134_) );
AND2X2 AND2X2_5 ( .A(_134_), .B(_129_), .Y(_135_) );
INVX1 INVX1_21 ( .A(_135_), .Y(w_C_23_) );
AND2X2 AND2X2_6 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_136_) );
INVX1 INVX1_22 ( .A(_136_), .Y(_137_) );
NAND3X1 NAND3X1_6 ( .A(_129_), .B(_137_), .C(_134_), .Y(_138_) );
OAI21X1 OAI21X1_3 ( .A(i_add2[23]), .B(i_add1[23]), .C(_138_), .Y(_139_) );
INVX1 INVX1_23 ( .A(_139_), .Y(w_C_24_) );
INVX1 INVX1_24 ( .A(i_add2[24]), .Y(_140_) );
INVX1 INVX1_25 ( .A(i_add1[24]), .Y(_141_) );
NOR2X1 NOR2X1_10 ( .A(_140_), .B(_141_), .Y(_142_) );
INVX1 INVX1_26 ( .A(_142_), .Y(_143_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_144_) );
INVX1 INVX1_27 ( .A(_144_), .Y(_145_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_146_) );
INVX1 INVX1_28 ( .A(_146_), .Y(_147_) );
NAND3X1 NAND3X1_7 ( .A(_145_), .B(_147_), .C(_138_), .Y(_148_) );
AND2X2 AND2X2_7 ( .A(_148_), .B(_143_), .Y(_149_) );
INVX1 INVX1_29 ( .A(_149_), .Y(w_C_25_) );
AND2X2 AND2X2_8 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_150_) );
INVX1 INVX1_30 ( .A(_150_), .Y(_151_) );
NAND3X1 NAND3X1_8 ( .A(_143_), .B(_151_), .C(_148_), .Y(_152_) );
OAI21X1 OAI21X1_4 ( .A(i_add2[25]), .B(i_add1[25]), .C(_152_), .Y(_153_) );
INVX1 INVX1_31 ( .A(_153_), .Y(w_C_26_) );
BUFX2 BUFX2_1 ( .A(_319__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_319__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_319__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_319__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_319__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_319__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_319__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_319__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_319__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_319__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_319__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_319__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_319__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_319__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_319__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_319__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_319__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_319__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_319__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_319__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_319__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_319__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_319__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_319__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_319__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_319__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_319__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_319__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_319__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_319__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_319__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_319__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_319__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_319__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_319__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_319__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_319__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(_319__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .A(_319__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .A(_319__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .A(_319__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .A(_319__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .A(_319__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .A(_319__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .A(_319__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .A(_319__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .A(_319__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .A(_319__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .A(_319__48_), .Y(o_result[48]) );
BUFX2 BUFX2_50 ( .A(_319__49_), .Y(o_result[49]) );
BUFX2 BUFX2_51 ( .A(_319__50_), .Y(o_result[50]) );
BUFX2 BUFX2_52 ( .A(_319__51_), .Y(o_result[51]) );
BUFX2 BUFX2_53 ( .A(_319__52_), .Y(o_result[52]) );
BUFX2 BUFX2_54 ( .A(w_C_53_), .Y(o_result[53]) );
INVX1 INVX1_32 ( .A(w_C_4_), .Y(_323_) );
OR2X2 OR2X2_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_324_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_325_) );
NAND3X1 NAND3X1_9 ( .A(_323_), .B(_325_), .C(_324_), .Y(_326_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_320_) );
AND2X2 AND2X2_9 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_321_) );
OAI21X1 OAI21X1_5 ( .A(_320_), .B(_321_), .C(w_C_4_), .Y(_322_) );
NAND2X1 NAND2X1_2 ( .A(_322_), .B(_326_), .Y(_319__4_) );
INVX1 INVX1_33 ( .A(w_C_5_), .Y(_330_) );
OR2X2 OR2X2_2 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_331_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_332_) );
NAND3X1 NAND3X1_10 ( .A(_330_), .B(_332_), .C(_331_), .Y(_333_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_327_) );
AND2X2 AND2X2_10 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_328_) );
OAI21X1 OAI21X1_6 ( .A(_327_), .B(_328_), .C(w_C_5_), .Y(_329_) );
NAND2X1 NAND2X1_4 ( .A(_329_), .B(_333_), .Y(_319__5_) );
INVX1 INVX1_34 ( .A(w_C_6_), .Y(_337_) );
OR2X2 OR2X2_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_338_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_339_) );
NAND3X1 NAND3X1_11 ( .A(_337_), .B(_339_), .C(_338_), .Y(_340_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_334_) );
AND2X2 AND2X2_11 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_335_) );
OAI21X1 OAI21X1_7 ( .A(_334_), .B(_335_), .C(w_C_6_), .Y(_336_) );
NAND2X1 NAND2X1_6 ( .A(_336_), .B(_340_), .Y(_319__6_) );
INVX1 INVX1_35 ( .A(w_C_7_), .Y(_344_) );
OR2X2 OR2X2_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_345_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_346_) );
NAND3X1 NAND3X1_12 ( .A(_344_), .B(_346_), .C(_345_), .Y(_347_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_341_) );
AND2X2 AND2X2_12 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_342_) );
OAI21X1 OAI21X1_8 ( .A(_341_), .B(_342_), .C(w_C_7_), .Y(_343_) );
NAND2X1 NAND2X1_8 ( .A(_343_), .B(_347_), .Y(_319__7_) );
INVX1 INVX1_36 ( .A(w_C_8_), .Y(_351_) );
OR2X2 OR2X2_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_352_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_353_) );
NAND3X1 NAND3X1_13 ( .A(_351_), .B(_353_), .C(_352_), .Y(_354_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_348_) );
AND2X2 AND2X2_13 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_349_) );
OAI21X1 OAI21X1_9 ( .A(_348_), .B(_349_), .C(w_C_8_), .Y(_350_) );
NAND2X1 NAND2X1_10 ( .A(_350_), .B(_354_), .Y(_319__8_) );
INVX1 INVX1_37 ( .A(w_C_9_), .Y(_358_) );
OR2X2 OR2X2_6 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_359_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_360_) );
NAND3X1 NAND3X1_14 ( .A(_358_), .B(_360_), .C(_359_), .Y(_361_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_355_) );
AND2X2 AND2X2_14 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_356_) );
OAI21X1 OAI21X1_10 ( .A(_355_), .B(_356_), .C(w_C_9_), .Y(_357_) );
NAND2X1 NAND2X1_12 ( .A(_357_), .B(_361_), .Y(_319__9_) );
INVX1 INVX1_38 ( .A(w_C_10_), .Y(_365_) );
OR2X2 OR2X2_7 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_366_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_367_) );
NAND3X1 NAND3X1_15 ( .A(_365_), .B(_367_), .C(_366_), .Y(_368_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_362_) );
AND2X2 AND2X2_15 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_363_) );
OAI21X1 OAI21X1_11 ( .A(_362_), .B(_363_), .C(w_C_10_), .Y(_364_) );
NAND2X1 NAND2X1_14 ( .A(_364_), .B(_368_), .Y(_319__10_) );
INVX1 INVX1_39 ( .A(w_C_11_), .Y(_372_) );
OR2X2 OR2X2_8 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_373_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_374_) );
NAND3X1 NAND3X1_16 ( .A(_372_), .B(_374_), .C(_373_), .Y(_375_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_369_) );
AND2X2 AND2X2_16 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_370_) );
OAI21X1 OAI21X1_12 ( .A(_369_), .B(_370_), .C(w_C_11_), .Y(_371_) );
NAND2X1 NAND2X1_16 ( .A(_371_), .B(_375_), .Y(_319__11_) );
INVX1 INVX1_40 ( .A(w_C_12_), .Y(_379_) );
OR2X2 OR2X2_9 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_380_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_381_) );
NAND3X1 NAND3X1_17 ( .A(_379_), .B(_381_), .C(_380_), .Y(_382_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_376_) );
AND2X2 AND2X2_17 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_377_) );
OAI21X1 OAI21X1_13 ( .A(_376_), .B(_377_), .C(w_C_12_), .Y(_378_) );
NAND2X1 NAND2X1_18 ( .A(_378_), .B(_382_), .Y(_319__12_) );
INVX1 INVX1_41 ( .A(w_C_13_), .Y(_386_) );
OR2X2 OR2X2_10 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_387_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_388_) );
NAND3X1 NAND3X1_18 ( .A(_386_), .B(_388_), .C(_387_), .Y(_389_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_383_) );
AND2X2 AND2X2_18 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_384_) );
OAI21X1 OAI21X1_14 ( .A(_383_), .B(_384_), .C(w_C_13_), .Y(_385_) );
NAND2X1 NAND2X1_20 ( .A(_385_), .B(_389_), .Y(_319__13_) );
INVX1 INVX1_42 ( .A(w_C_14_), .Y(_393_) );
OR2X2 OR2X2_11 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_394_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_395_) );
NAND3X1 NAND3X1_19 ( .A(_393_), .B(_395_), .C(_394_), .Y(_396_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_390_) );
AND2X2 AND2X2_19 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_391_) );
OAI21X1 OAI21X1_15 ( .A(_390_), .B(_391_), .C(w_C_14_), .Y(_392_) );
NAND2X1 NAND2X1_22 ( .A(_392_), .B(_396_), .Y(_319__14_) );
INVX1 INVX1_43 ( .A(w_C_15_), .Y(_400_) );
OR2X2 OR2X2_12 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_401_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_402_) );
NAND3X1 NAND3X1_20 ( .A(_400_), .B(_402_), .C(_401_), .Y(_403_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_397_) );
AND2X2 AND2X2_20 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_398_) );
OAI21X1 OAI21X1_16 ( .A(_397_), .B(_398_), .C(w_C_15_), .Y(_399_) );
NAND2X1 NAND2X1_24 ( .A(_399_), .B(_403_), .Y(_319__15_) );
INVX1 INVX1_44 ( .A(w_C_16_), .Y(_407_) );
OR2X2 OR2X2_13 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_408_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_409_) );
NAND3X1 NAND3X1_21 ( .A(_407_), .B(_409_), .C(_408_), .Y(_410_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_404_) );
AND2X2 AND2X2_21 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_405_) );
OAI21X1 OAI21X1_17 ( .A(_404_), .B(_405_), .C(w_C_16_), .Y(_406_) );
NAND2X1 NAND2X1_26 ( .A(_406_), .B(_410_), .Y(_319__16_) );
INVX1 INVX1_45 ( .A(w_C_17_), .Y(_414_) );
OR2X2 OR2X2_14 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_415_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_416_) );
NAND3X1 NAND3X1_22 ( .A(_414_), .B(_416_), .C(_415_), .Y(_417_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_411_) );
AND2X2 AND2X2_22 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_412_) );
OAI21X1 OAI21X1_18 ( .A(_411_), .B(_412_), .C(w_C_17_), .Y(_413_) );
NAND2X1 NAND2X1_28 ( .A(_413_), .B(_417_), .Y(_319__17_) );
INVX1 INVX1_46 ( .A(w_C_18_), .Y(_421_) );
OR2X2 OR2X2_15 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_422_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_423_) );
NAND3X1 NAND3X1_23 ( .A(_421_), .B(_423_), .C(_422_), .Y(_424_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_418_) );
AND2X2 AND2X2_23 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_419_) );
OAI21X1 OAI21X1_19 ( .A(_418_), .B(_419_), .C(w_C_18_), .Y(_420_) );
NAND2X1 NAND2X1_30 ( .A(_420_), .B(_424_), .Y(_319__18_) );
INVX1 INVX1_47 ( .A(w_C_19_), .Y(_428_) );
OR2X2 OR2X2_16 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_429_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_430_) );
NAND3X1 NAND3X1_24 ( .A(_428_), .B(_430_), .C(_429_), .Y(_431_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_425_) );
AND2X2 AND2X2_24 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_426_) );
OAI21X1 OAI21X1_20 ( .A(_425_), .B(_426_), .C(w_C_19_), .Y(_427_) );
NAND2X1 NAND2X1_32 ( .A(_427_), .B(_431_), .Y(_319__19_) );
INVX1 INVX1_48 ( .A(w_C_20_), .Y(_435_) );
OR2X2 OR2X2_17 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_436_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_437_) );
NAND3X1 NAND3X1_25 ( .A(_435_), .B(_437_), .C(_436_), .Y(_438_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_432_) );
AND2X2 AND2X2_25 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_433_) );
OAI21X1 OAI21X1_21 ( .A(_432_), .B(_433_), .C(w_C_20_), .Y(_434_) );
NAND2X1 NAND2X1_34 ( .A(_434_), .B(_438_), .Y(_319__20_) );
INVX1 INVX1_49 ( .A(w_C_21_), .Y(_442_) );
OR2X2 OR2X2_18 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_443_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_444_) );
NAND3X1 NAND3X1_26 ( .A(_442_), .B(_444_), .C(_443_), .Y(_445_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_439_) );
AND2X2 AND2X2_26 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_440_) );
OAI21X1 OAI21X1_22 ( .A(_439_), .B(_440_), .C(w_C_21_), .Y(_441_) );
NAND2X1 NAND2X1_36 ( .A(_441_), .B(_445_), .Y(_319__21_) );
INVX1 INVX1_50 ( .A(w_C_22_), .Y(_449_) );
OR2X2 OR2X2_19 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_450_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_451_) );
NAND3X1 NAND3X1_27 ( .A(_449_), .B(_451_), .C(_450_), .Y(_452_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_446_) );
AND2X2 AND2X2_27 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_447_) );
OAI21X1 OAI21X1_23 ( .A(_446_), .B(_447_), .C(w_C_22_), .Y(_448_) );
NAND2X1 NAND2X1_38 ( .A(_448_), .B(_452_), .Y(_319__22_) );
INVX1 INVX1_51 ( .A(w_C_23_), .Y(_456_) );
OR2X2 OR2X2_20 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_457_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_458_) );
NAND3X1 NAND3X1_28 ( .A(_456_), .B(_458_), .C(_457_), .Y(_459_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_453_) );
AND2X2 AND2X2_28 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_454_) );
OAI21X1 OAI21X1_24 ( .A(_453_), .B(_454_), .C(w_C_23_), .Y(_455_) );
NAND2X1 NAND2X1_40 ( .A(_455_), .B(_459_), .Y(_319__23_) );
INVX1 INVX1_52 ( .A(w_C_24_), .Y(_463_) );
OR2X2 OR2X2_21 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_464_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_465_) );
NAND3X1 NAND3X1_29 ( .A(_463_), .B(_465_), .C(_464_), .Y(_466_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_460_) );
AND2X2 AND2X2_29 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_461_) );
OAI21X1 OAI21X1_25 ( .A(_460_), .B(_461_), .C(w_C_24_), .Y(_462_) );
NAND2X1 NAND2X1_42 ( .A(_462_), .B(_466_), .Y(_319__24_) );
INVX1 INVX1_53 ( .A(w_C_25_), .Y(_470_) );
OR2X2 OR2X2_22 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_471_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_472_) );
NAND3X1 NAND3X1_30 ( .A(_470_), .B(_472_), .C(_471_), .Y(_473_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_467_) );
AND2X2 AND2X2_30 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_468_) );
OAI21X1 OAI21X1_26 ( .A(_467_), .B(_468_), .C(w_C_25_), .Y(_469_) );
NAND2X1 NAND2X1_44 ( .A(_469_), .B(_473_), .Y(_319__25_) );
INVX1 INVX1_54 ( .A(w_C_26_), .Y(_477_) );
OR2X2 OR2X2_23 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_478_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_479_) );
NAND3X1 NAND3X1_31 ( .A(_477_), .B(_479_), .C(_478_), .Y(_480_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_474_) );
AND2X2 AND2X2_31 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_475_) );
OAI21X1 OAI21X1_27 ( .A(_474_), .B(_475_), .C(w_C_26_), .Y(_476_) );
NAND2X1 NAND2X1_46 ( .A(_476_), .B(_480_), .Y(_319__26_) );
INVX1 INVX1_55 ( .A(w_C_27_), .Y(_484_) );
OR2X2 OR2X2_24 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_485_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_486_) );
NAND3X1 NAND3X1_32 ( .A(_484_), .B(_486_), .C(_485_), .Y(_487_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_481_) );
AND2X2 AND2X2_32 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_482_) );
OAI21X1 OAI21X1_28 ( .A(_481_), .B(_482_), .C(w_C_27_), .Y(_483_) );
NAND2X1 NAND2X1_48 ( .A(_483_), .B(_487_), .Y(_319__27_) );
INVX1 INVX1_56 ( .A(w_C_28_), .Y(_491_) );
OR2X2 OR2X2_25 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_492_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_493_) );
NAND3X1 NAND3X1_33 ( .A(_491_), .B(_493_), .C(_492_), .Y(_494_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_488_) );
AND2X2 AND2X2_33 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_489_) );
OAI21X1 OAI21X1_29 ( .A(_488_), .B(_489_), .C(w_C_28_), .Y(_490_) );
NAND2X1 NAND2X1_50 ( .A(_490_), .B(_494_), .Y(_319__28_) );
INVX1 INVX1_57 ( .A(w_C_29_), .Y(_498_) );
OR2X2 OR2X2_26 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_499_) );
NAND2X1 NAND2X1_51 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_500_) );
NAND3X1 NAND3X1_34 ( .A(_498_), .B(_500_), .C(_499_), .Y(_501_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_495_) );
AND2X2 AND2X2_34 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_496_) );
OAI21X1 OAI21X1_30 ( .A(_495_), .B(_496_), .C(w_C_29_), .Y(_497_) );
NAND2X1 NAND2X1_52 ( .A(_497_), .B(_501_), .Y(_319__29_) );
INVX1 INVX1_58 ( .A(w_C_30_), .Y(_505_) );
OR2X2 OR2X2_27 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_506_) );
NAND2X1 NAND2X1_53 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_507_) );
NAND3X1 NAND3X1_35 ( .A(_505_), .B(_507_), .C(_506_), .Y(_508_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_502_) );
AND2X2 AND2X2_35 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_503_) );
OAI21X1 OAI21X1_31 ( .A(_502_), .B(_503_), .C(w_C_30_), .Y(_504_) );
NAND2X1 NAND2X1_54 ( .A(_504_), .B(_508_), .Y(_319__30_) );
INVX1 INVX1_59 ( .A(w_C_31_), .Y(_512_) );
OR2X2 OR2X2_28 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_513_) );
NAND2X1 NAND2X1_55 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_514_) );
NAND3X1 NAND3X1_36 ( .A(_512_), .B(_514_), .C(_513_), .Y(_515_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_509_) );
AND2X2 AND2X2_36 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_510_) );
OAI21X1 OAI21X1_32 ( .A(_509_), .B(_510_), .C(w_C_31_), .Y(_511_) );
NAND2X1 NAND2X1_56 ( .A(_511_), .B(_515_), .Y(_319__31_) );
INVX1 INVX1_60 ( .A(w_C_32_), .Y(_519_) );
OR2X2 OR2X2_29 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_520_) );
NAND2X1 NAND2X1_57 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_521_) );
NAND3X1 NAND3X1_37 ( .A(_519_), .B(_521_), .C(_520_), .Y(_522_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_516_) );
AND2X2 AND2X2_37 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_517_) );
OAI21X1 OAI21X1_33 ( .A(_516_), .B(_517_), .C(w_C_32_), .Y(_518_) );
NAND2X1 NAND2X1_58 ( .A(_518_), .B(_522_), .Y(_319__32_) );
INVX1 INVX1_61 ( .A(w_C_33_), .Y(_526_) );
OR2X2 OR2X2_30 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_527_) );
NAND2X1 NAND2X1_59 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_528_) );
NAND3X1 NAND3X1_38 ( .A(_526_), .B(_528_), .C(_527_), .Y(_529_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_523_) );
AND2X2 AND2X2_38 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_524_) );
OAI21X1 OAI21X1_34 ( .A(_523_), .B(_524_), .C(w_C_33_), .Y(_525_) );
NAND2X1 NAND2X1_60 ( .A(_525_), .B(_529_), .Y(_319__33_) );
INVX1 INVX1_62 ( .A(w_C_34_), .Y(_533_) );
OR2X2 OR2X2_31 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_534_) );
NAND2X1 NAND2X1_61 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_535_) );
NAND3X1 NAND3X1_39 ( .A(_533_), .B(_535_), .C(_534_), .Y(_536_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_530_) );
AND2X2 AND2X2_39 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_531_) );
OAI21X1 OAI21X1_35 ( .A(_530_), .B(_531_), .C(w_C_34_), .Y(_532_) );
NAND2X1 NAND2X1_62 ( .A(_532_), .B(_536_), .Y(_319__34_) );
INVX1 INVX1_63 ( .A(w_C_35_), .Y(_540_) );
OR2X2 OR2X2_32 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_541_) );
NAND2X1 NAND2X1_63 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_542_) );
NAND3X1 NAND3X1_40 ( .A(_540_), .B(_542_), .C(_541_), .Y(_543_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_537_) );
AND2X2 AND2X2_40 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_538_) );
OAI21X1 OAI21X1_36 ( .A(_537_), .B(_538_), .C(w_C_35_), .Y(_539_) );
NAND2X1 NAND2X1_64 ( .A(_539_), .B(_543_), .Y(_319__35_) );
INVX1 INVX1_64 ( .A(w_C_36_), .Y(_547_) );
OR2X2 OR2X2_33 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_548_) );
NAND2X1 NAND2X1_65 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_549_) );
NAND3X1 NAND3X1_41 ( .A(_547_), .B(_549_), .C(_548_), .Y(_550_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_544_) );
AND2X2 AND2X2_41 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_545_) );
OAI21X1 OAI21X1_37 ( .A(_544_), .B(_545_), .C(w_C_36_), .Y(_546_) );
NAND2X1 NAND2X1_66 ( .A(_546_), .B(_550_), .Y(_319__36_) );
INVX1 INVX1_65 ( .A(w_C_37_), .Y(_554_) );
OR2X2 OR2X2_34 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_555_) );
NAND2X1 NAND2X1_67 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_556_) );
NAND3X1 NAND3X1_42 ( .A(_554_), .B(_556_), .C(_555_), .Y(_557_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_551_) );
AND2X2 AND2X2_42 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_552_) );
OAI21X1 OAI21X1_38 ( .A(_551_), .B(_552_), .C(w_C_37_), .Y(_553_) );
NAND2X1 NAND2X1_68 ( .A(_553_), .B(_557_), .Y(_319__37_) );
INVX1 INVX1_66 ( .A(w_C_38_), .Y(_561_) );
OR2X2 OR2X2_35 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_562_) );
NAND2X1 NAND2X1_69 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_563_) );
NAND3X1 NAND3X1_43 ( .A(_561_), .B(_563_), .C(_562_), .Y(_564_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_558_) );
AND2X2 AND2X2_43 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_559_) );
OAI21X1 OAI21X1_39 ( .A(_558_), .B(_559_), .C(w_C_38_), .Y(_560_) );
NAND2X1 NAND2X1_70 ( .A(_560_), .B(_564_), .Y(_319__38_) );
INVX1 INVX1_67 ( .A(w_C_39_), .Y(_568_) );
OR2X2 OR2X2_36 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_569_) );
NAND2X1 NAND2X1_71 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_570_) );
NAND3X1 NAND3X1_44 ( .A(_568_), .B(_570_), .C(_569_), .Y(_571_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_565_) );
AND2X2 AND2X2_44 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_566_) );
OAI21X1 OAI21X1_40 ( .A(_565_), .B(_566_), .C(w_C_39_), .Y(_567_) );
NAND2X1 NAND2X1_72 ( .A(_567_), .B(_571_), .Y(_319__39_) );
INVX1 INVX1_68 ( .A(w_C_40_), .Y(_575_) );
OR2X2 OR2X2_37 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_576_) );
NAND2X1 NAND2X1_73 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_577_) );
NAND3X1 NAND3X1_45 ( .A(_575_), .B(_577_), .C(_576_), .Y(_578_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_572_) );
AND2X2 AND2X2_45 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_573_) );
OAI21X1 OAI21X1_41 ( .A(_572_), .B(_573_), .C(w_C_40_), .Y(_574_) );
NAND2X1 NAND2X1_74 ( .A(_574_), .B(_578_), .Y(_319__40_) );
INVX1 INVX1_69 ( .A(w_C_41_), .Y(_582_) );
OR2X2 OR2X2_38 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_583_) );
NAND2X1 NAND2X1_75 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_584_) );
NAND3X1 NAND3X1_46 ( .A(_582_), .B(_584_), .C(_583_), .Y(_585_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_579_) );
AND2X2 AND2X2_46 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_580_) );
OAI21X1 OAI21X1_42 ( .A(_579_), .B(_580_), .C(w_C_41_), .Y(_581_) );
NAND2X1 NAND2X1_76 ( .A(_581_), .B(_585_), .Y(_319__41_) );
INVX1 INVX1_70 ( .A(w_C_42_), .Y(_589_) );
OR2X2 OR2X2_39 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_590_) );
NAND2X1 NAND2X1_77 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_591_) );
NAND3X1 NAND3X1_47 ( .A(_589_), .B(_591_), .C(_590_), .Y(_592_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_586_) );
AND2X2 AND2X2_47 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_587_) );
OAI21X1 OAI21X1_43 ( .A(_586_), .B(_587_), .C(w_C_42_), .Y(_588_) );
NAND2X1 NAND2X1_78 ( .A(_588_), .B(_592_), .Y(_319__42_) );
INVX1 INVX1_71 ( .A(w_C_43_), .Y(_596_) );
OR2X2 OR2X2_40 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_597_) );
NAND2X1 NAND2X1_79 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_598_) );
NAND3X1 NAND3X1_48 ( .A(_596_), .B(_598_), .C(_597_), .Y(_599_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_593_) );
AND2X2 AND2X2_48 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_594_) );
OAI21X1 OAI21X1_44 ( .A(_593_), .B(_594_), .C(w_C_43_), .Y(_595_) );
NAND2X1 NAND2X1_80 ( .A(_595_), .B(_599_), .Y(_319__43_) );
INVX1 INVX1_72 ( .A(w_C_44_), .Y(_603_) );
OR2X2 OR2X2_41 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_604_) );
NAND2X1 NAND2X1_81 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_605_) );
NAND3X1 NAND3X1_49 ( .A(_603_), .B(_605_), .C(_604_), .Y(_606_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_600_) );
AND2X2 AND2X2_49 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_601_) );
OAI21X1 OAI21X1_45 ( .A(_600_), .B(_601_), .C(w_C_44_), .Y(_602_) );
NAND2X1 NAND2X1_82 ( .A(_602_), .B(_606_), .Y(_319__44_) );
INVX1 INVX1_73 ( .A(w_C_45_), .Y(_610_) );
OR2X2 OR2X2_42 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_611_) );
NAND2X1 NAND2X1_83 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_612_) );
NAND3X1 NAND3X1_50 ( .A(_610_), .B(_612_), .C(_611_), .Y(_613_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_607_) );
AND2X2 AND2X2_50 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_608_) );
OAI21X1 OAI21X1_46 ( .A(_607_), .B(_608_), .C(w_C_45_), .Y(_609_) );
NAND2X1 NAND2X1_84 ( .A(_609_), .B(_613_), .Y(_319__45_) );
INVX1 INVX1_74 ( .A(w_C_46_), .Y(_617_) );
OR2X2 OR2X2_43 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_618_) );
NAND2X1 NAND2X1_85 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_619_) );
NAND3X1 NAND3X1_51 ( .A(_617_), .B(_619_), .C(_618_), .Y(_620_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_614_) );
AND2X2 AND2X2_51 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_615_) );
OAI21X1 OAI21X1_47 ( .A(_614_), .B(_615_), .C(w_C_46_), .Y(_616_) );
NAND2X1 NAND2X1_86 ( .A(_616_), .B(_620_), .Y(_319__46_) );
INVX1 INVX1_75 ( .A(w_C_47_), .Y(_624_) );
OR2X2 OR2X2_44 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_625_) );
NAND2X1 NAND2X1_87 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_626_) );
NAND3X1 NAND3X1_52 ( .A(_624_), .B(_626_), .C(_625_), .Y(_627_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_621_) );
AND2X2 AND2X2_52 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_622_) );
OAI21X1 OAI21X1_48 ( .A(_621_), .B(_622_), .C(w_C_47_), .Y(_623_) );
NAND2X1 NAND2X1_88 ( .A(_623_), .B(_627_), .Y(_319__47_) );
INVX1 INVX1_76 ( .A(w_C_48_), .Y(_631_) );
OR2X2 OR2X2_45 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_632_) );
NAND2X1 NAND2X1_89 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_633_) );
NAND3X1 NAND3X1_53 ( .A(_631_), .B(_633_), .C(_632_), .Y(_634_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_628_) );
AND2X2 AND2X2_53 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_629_) );
OAI21X1 OAI21X1_49 ( .A(_628_), .B(_629_), .C(w_C_48_), .Y(_630_) );
NAND2X1 NAND2X1_90 ( .A(_630_), .B(_634_), .Y(_319__48_) );
INVX1 INVX1_77 ( .A(w_C_49_), .Y(_638_) );
OR2X2 OR2X2_46 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_639_) );
NAND2X1 NAND2X1_91 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_640_) );
NAND3X1 NAND3X1_54 ( .A(_638_), .B(_640_), .C(_639_), .Y(_641_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_635_) );
AND2X2 AND2X2_54 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_636_) );
OAI21X1 OAI21X1_50 ( .A(_635_), .B(_636_), .C(w_C_49_), .Y(_637_) );
NAND2X1 NAND2X1_92 ( .A(_637_), .B(_641_), .Y(_319__49_) );
INVX1 INVX1_78 ( .A(w_C_50_), .Y(_645_) );
OR2X2 OR2X2_47 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_646_) );
NAND2X1 NAND2X1_93 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_647_) );
NAND3X1 NAND3X1_55 ( .A(_645_), .B(_647_), .C(_646_), .Y(_648_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_642_) );
AND2X2 AND2X2_55 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_643_) );
OAI21X1 OAI21X1_51 ( .A(_642_), .B(_643_), .C(w_C_50_), .Y(_644_) );
NAND2X1 NAND2X1_94 ( .A(_644_), .B(_648_), .Y(_319__50_) );
INVX1 INVX1_79 ( .A(w_C_51_), .Y(_652_) );
OR2X2 OR2X2_48 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_653_) );
NAND2X1 NAND2X1_95 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_654_) );
NAND3X1 NAND3X1_56 ( .A(_652_), .B(_654_), .C(_653_), .Y(_655_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_649_) );
AND2X2 AND2X2_56 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_650_) );
OAI21X1 OAI21X1_52 ( .A(_649_), .B(_650_), .C(w_C_51_), .Y(_651_) );
NAND2X1 NAND2X1_96 ( .A(_651_), .B(_655_), .Y(_319__51_) );
INVX1 INVX1_80 ( .A(w_C_52_), .Y(_659_) );
OR2X2 OR2X2_49 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_660_) );
NAND2X1 NAND2X1_97 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_661_) );
NAND3X1 NAND3X1_57 ( .A(_659_), .B(_661_), .C(_660_), .Y(_662_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_656_) );
AND2X2 AND2X2_57 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_657_) );
OAI21X1 OAI21X1_53 ( .A(_656_), .B(_657_), .C(w_C_52_), .Y(_658_) );
NAND2X1 NAND2X1_98 ( .A(_658_), .B(_662_), .Y(_319__52_) );
INVX1 INVX1_81 ( .A(gnd), .Y(_666_) );
OR2X2 OR2X2_50 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_667_) );
NAND2X1 NAND2X1_99 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_668_) );
NAND3X1 NAND3X1_58 ( .A(_666_), .B(_668_), .C(_667_), .Y(_669_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_663_) );
AND2X2 AND2X2_58 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_664_) );
OAI21X1 OAI21X1_54 ( .A(_663_), .B(_664_), .C(gnd), .Y(_665_) );
NAND2X1 NAND2X1_100 ( .A(_665_), .B(_669_), .Y(_319__0_) );
INVX1 INVX1_82 ( .A(w_C_1_), .Y(_673_) );
OR2X2 OR2X2_51 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_674_) );
NAND2X1 NAND2X1_101 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_675_) );
NAND3X1 NAND3X1_59 ( .A(_673_), .B(_675_), .C(_674_), .Y(_676_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_670_) );
AND2X2 AND2X2_59 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_671_) );
OAI21X1 OAI21X1_55 ( .A(_670_), .B(_671_), .C(w_C_1_), .Y(_672_) );
NAND2X1 NAND2X1_102 ( .A(_672_), .B(_676_), .Y(_319__1_) );
INVX1 INVX1_83 ( .A(w_C_2_), .Y(_680_) );
OR2X2 OR2X2_52 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_681_) );
NAND2X1 NAND2X1_103 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_682_) );
NAND3X1 NAND3X1_60 ( .A(_680_), .B(_682_), .C(_681_), .Y(_683_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_677_) );
AND2X2 AND2X2_60 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_678_) );
OAI21X1 OAI21X1_56 ( .A(_677_), .B(_678_), .C(w_C_2_), .Y(_679_) );
NAND2X1 NAND2X1_104 ( .A(_679_), .B(_683_), .Y(_319__2_) );
INVX1 INVX1_84 ( .A(w_C_3_), .Y(_687_) );
OR2X2 OR2X2_53 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_688_) );
NAND2X1 NAND2X1_105 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_689_) );
NAND3X1 NAND3X1_61 ( .A(_687_), .B(_689_), .C(_688_), .Y(_690_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_684_) );
AND2X2 AND2X2_61 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_685_) );
OAI21X1 OAI21X1_57 ( .A(_684_), .B(_685_), .C(w_C_3_), .Y(_686_) );
NAND2X1 NAND2X1_106 ( .A(_686_), .B(_690_), .Y(_319__3_) );
INVX1 INVX1_85 ( .A(i_add2[26]), .Y(_154_) );
INVX1 INVX1_86 ( .A(i_add1[26]), .Y(_155_) );
NOR2X1 NOR2X1_66 ( .A(_154_), .B(_155_), .Y(_156_) );
INVX1 INVX1_87 ( .A(_156_), .Y(_157_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_158_) );
INVX1 INVX1_88 ( .A(_158_), .Y(_159_) );
NOR2X1 NOR2X1_68 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_160_) );
INVX1 INVX1_89 ( .A(_160_), .Y(_161_) );
NAND3X1 NAND3X1_62 ( .A(_159_), .B(_161_), .C(_152_), .Y(_162_) );
AND2X2 AND2X2_62 ( .A(_162_), .B(_157_), .Y(_163_) );
INVX1 INVX1_90 ( .A(_163_), .Y(w_C_27_) );
AND2X2 AND2X2_63 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_164_) );
INVX1 INVX1_91 ( .A(_164_), .Y(_165_) );
NAND3X1 NAND3X1_63 ( .A(_157_), .B(_165_), .C(_162_), .Y(_166_) );
OAI21X1 OAI21X1_58 ( .A(i_add2[27]), .B(i_add1[27]), .C(_166_), .Y(_167_) );
INVX1 INVX1_92 ( .A(_167_), .Y(w_C_28_) );
INVX1 INVX1_93 ( .A(i_add2[28]), .Y(_168_) );
INVX1 INVX1_94 ( .A(i_add1[28]), .Y(_169_) );
NOR2X1 NOR2X1_69 ( .A(_168_), .B(_169_), .Y(_170_) );
INVX1 INVX1_95 ( .A(_170_), .Y(_171_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_172_) );
INVX1 INVX1_96 ( .A(_172_), .Y(_173_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_174_) );
INVX1 INVX1_97 ( .A(_174_), .Y(_175_) );
NAND3X1 NAND3X1_64 ( .A(_173_), .B(_175_), .C(_166_), .Y(_176_) );
AND2X2 AND2X2_64 ( .A(_176_), .B(_171_), .Y(_177_) );
INVX1 INVX1_98 ( .A(_177_), .Y(w_C_29_) );
AND2X2 AND2X2_65 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_178_) );
INVX1 INVX1_99 ( .A(_178_), .Y(_179_) );
NAND3X1 NAND3X1_65 ( .A(_171_), .B(_179_), .C(_176_), .Y(_180_) );
OAI21X1 OAI21X1_59 ( .A(i_add2[29]), .B(i_add1[29]), .C(_180_), .Y(_181_) );
INVX1 INVX1_100 ( .A(_181_), .Y(w_C_30_) );
INVX1 INVX1_101 ( .A(i_add2[30]), .Y(_182_) );
INVX1 INVX1_102 ( .A(i_add1[30]), .Y(_183_) );
NOR2X1 NOR2X1_72 ( .A(_182_), .B(_183_), .Y(_184_) );
INVX1 INVX1_103 ( .A(_184_), .Y(_185_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_186_) );
INVX1 INVX1_104 ( .A(_186_), .Y(_187_) );
NOR2X1 NOR2X1_74 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_188_) );
INVX1 INVX1_105 ( .A(_188_), .Y(_189_) );
NAND3X1 NAND3X1_66 ( .A(_187_), .B(_189_), .C(_180_), .Y(_190_) );
AND2X2 AND2X2_66 ( .A(_190_), .B(_185_), .Y(_191_) );
INVX1 INVX1_106 ( .A(_191_), .Y(w_C_31_) );
AND2X2 AND2X2_67 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_192_) );
INVX1 INVX1_107 ( .A(_192_), .Y(_193_) );
NAND3X1 NAND3X1_67 ( .A(_185_), .B(_193_), .C(_190_), .Y(_194_) );
OAI21X1 OAI21X1_60 ( .A(i_add2[31]), .B(i_add1[31]), .C(_194_), .Y(_195_) );
INVX1 INVX1_108 ( .A(_195_), .Y(w_C_32_) );
INVX1 INVX1_109 ( .A(i_add2[32]), .Y(_196_) );
INVX1 INVX1_110 ( .A(i_add1[32]), .Y(_197_) );
NOR2X1 NOR2X1_75 ( .A(_196_), .B(_197_), .Y(_198_) );
INVX1 INVX1_111 ( .A(_198_), .Y(_199_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_200_) );
INVX1 INVX1_112 ( .A(_200_), .Y(_201_) );
NOR2X1 NOR2X1_77 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_202_) );
INVX1 INVX1_113 ( .A(_202_), .Y(_203_) );
NAND3X1 NAND3X1_68 ( .A(_201_), .B(_203_), .C(_194_), .Y(_204_) );
AND2X2 AND2X2_68 ( .A(_204_), .B(_199_), .Y(_205_) );
INVX1 INVX1_114 ( .A(_205_), .Y(w_C_33_) );
AND2X2 AND2X2_69 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_206_) );
INVX1 INVX1_115 ( .A(_206_), .Y(_207_) );
NAND3X1 NAND3X1_69 ( .A(_199_), .B(_207_), .C(_204_), .Y(_208_) );
OAI21X1 OAI21X1_61 ( .A(i_add2[33]), .B(i_add1[33]), .C(_208_), .Y(_209_) );
INVX1 INVX1_116 ( .A(_209_), .Y(w_C_34_) );
INVX1 INVX1_117 ( .A(i_add2[34]), .Y(_210_) );
INVX1 INVX1_118 ( .A(i_add1[34]), .Y(_211_) );
NOR2X1 NOR2X1_78 ( .A(_210_), .B(_211_), .Y(_212_) );
INVX1 INVX1_119 ( .A(_212_), .Y(_213_) );
NOR2X1 NOR2X1_79 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_214_) );
INVX1 INVX1_120 ( .A(_214_), .Y(_215_) );
NOR2X1 NOR2X1_80 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_216_) );
INVX1 INVX1_121 ( .A(_216_), .Y(_217_) );
NAND3X1 NAND3X1_70 ( .A(_215_), .B(_217_), .C(_208_), .Y(_218_) );
AND2X2 AND2X2_70 ( .A(_218_), .B(_213_), .Y(_219_) );
INVX1 INVX1_122 ( .A(_219_), .Y(w_C_35_) );
AND2X2 AND2X2_71 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_220_) );
INVX1 INVX1_123 ( .A(_220_), .Y(_221_) );
NAND3X1 NAND3X1_71 ( .A(_213_), .B(_221_), .C(_218_), .Y(_222_) );
OAI21X1 OAI21X1_62 ( .A(i_add2[35]), .B(i_add1[35]), .C(_222_), .Y(_223_) );
INVX1 INVX1_124 ( .A(_223_), .Y(w_C_36_) );
INVX1 INVX1_125 ( .A(i_add2[36]), .Y(_224_) );
INVX1 INVX1_126 ( .A(i_add1[36]), .Y(_225_) );
NOR2X1 NOR2X1_81 ( .A(_224_), .B(_225_), .Y(_226_) );
INVX1 INVX1_127 ( .A(_226_), .Y(_227_) );
NOR2X1 NOR2X1_82 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_228_) );
INVX1 INVX1_128 ( .A(_228_), .Y(_229_) );
NOR2X1 NOR2X1_83 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_230_) );
INVX1 INVX1_129 ( .A(_230_), .Y(_231_) );
NAND3X1 NAND3X1_72 ( .A(_229_), .B(_231_), .C(_222_), .Y(_232_) );
AND2X2 AND2X2_72 ( .A(_232_), .B(_227_), .Y(_233_) );
INVX1 INVX1_130 ( .A(_233_), .Y(w_C_37_) );
AND2X2 AND2X2_73 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_234_) );
INVX1 INVX1_131 ( .A(_234_), .Y(_235_) );
NAND3X1 NAND3X1_73 ( .A(_227_), .B(_235_), .C(_232_), .Y(_236_) );
OAI21X1 OAI21X1_63 ( .A(i_add2[37]), .B(i_add1[37]), .C(_236_), .Y(_237_) );
INVX1 INVX1_132 ( .A(_237_), .Y(w_C_38_) );
INVX1 INVX1_133 ( .A(i_add2[38]), .Y(_238_) );
INVX1 INVX1_134 ( .A(i_add1[38]), .Y(_239_) );
NOR2X1 NOR2X1_84 ( .A(_238_), .B(_239_), .Y(_240_) );
INVX1 INVX1_135 ( .A(_240_), .Y(_241_) );
NOR2X1 NOR2X1_85 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_242_) );
INVX1 INVX1_136 ( .A(_242_), .Y(_243_) );
NOR2X1 NOR2X1_86 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_244_) );
INVX1 INVX1_137 ( .A(_244_), .Y(_245_) );
NAND3X1 NAND3X1_74 ( .A(_243_), .B(_245_), .C(_236_), .Y(_246_) );
AND2X2 AND2X2_74 ( .A(_246_), .B(_241_), .Y(_247_) );
INVX1 INVX1_138 ( .A(_247_), .Y(w_C_39_) );
AND2X2 AND2X2_75 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_248_) );
INVX1 INVX1_139 ( .A(_248_), .Y(_249_) );
NAND3X1 NAND3X1_75 ( .A(_241_), .B(_249_), .C(_246_), .Y(_250_) );
OAI21X1 OAI21X1_64 ( .A(i_add2[39]), .B(i_add1[39]), .C(_250_), .Y(_251_) );
INVX1 INVX1_140 ( .A(_251_), .Y(w_C_40_) );
INVX1 INVX1_141 ( .A(i_add2[40]), .Y(_252_) );
INVX1 INVX1_142 ( .A(i_add1[40]), .Y(_253_) );
NOR2X1 NOR2X1_87 ( .A(_252_), .B(_253_), .Y(_254_) );
INVX1 INVX1_143 ( .A(_254_), .Y(_255_) );
NOR2X1 NOR2X1_88 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_256_) );
INVX1 INVX1_144 ( .A(_256_), .Y(_257_) );
NOR2X1 NOR2X1_89 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_258_) );
INVX1 INVX1_145 ( .A(_258_), .Y(_259_) );
NAND3X1 NAND3X1_76 ( .A(_257_), .B(_259_), .C(_250_), .Y(_260_) );
AND2X2 AND2X2_76 ( .A(_260_), .B(_255_), .Y(_261_) );
INVX1 INVX1_146 ( .A(_261_), .Y(w_C_41_) );
AND2X2 AND2X2_77 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_262_) );
INVX1 INVX1_147 ( .A(_262_), .Y(_263_) );
NAND3X1 NAND3X1_77 ( .A(_255_), .B(_263_), .C(_260_), .Y(_264_) );
OAI21X1 OAI21X1_65 ( .A(i_add2[41]), .B(i_add1[41]), .C(_264_), .Y(_265_) );
INVX1 INVX1_148 ( .A(_265_), .Y(w_C_42_) );
NAND2X1 NAND2X1_107 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_266_) );
NOR2X1 NOR2X1_90 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_267_) );
OAI21X1 OAI21X1_66 ( .A(_267_), .B(_265_), .C(_266_), .Y(w_C_43_) );
OR2X2 OR2X2_54 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_268_) );
NOR2X1 NOR2X1_91 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_269_) );
INVX1 INVX1_149 ( .A(_269_), .Y(_270_) );
INVX1 INVX1_150 ( .A(_267_), .Y(_271_) );
NAND3X1 NAND3X1_78 ( .A(_270_), .B(_271_), .C(_264_), .Y(_272_) );
NAND2X1 NAND2X1_108 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_273_) );
NAND3X1 NAND3X1_79 ( .A(_266_), .B(_273_), .C(_272_), .Y(_274_) );
AND2X2 AND2X2_78 ( .A(_274_), .B(_268_), .Y(w_C_44_) );
INVX1 INVX1_151 ( .A(i_add2[44]), .Y(_275_) );
INVX1 INVX1_152 ( .A(i_add1[44]), .Y(_276_) );
NAND2X1 NAND2X1_109 ( .A(_275_), .B(_276_), .Y(_277_) );
NAND3X1 NAND3X1_80 ( .A(_268_), .B(_277_), .C(_274_), .Y(_278_) );
OAI21X1 OAI21X1_67 ( .A(_275_), .B(_276_), .C(_278_), .Y(w_C_45_) );
INVX1 INVX1_153 ( .A(i_add2[45]), .Y(_279_) );
INVX1 INVX1_154 ( .A(i_add1[45]), .Y(_280_) );
NAND2X1 NAND2X1_110 ( .A(_279_), .B(_280_), .Y(_281_) );
NAND2X1 NAND2X1_111 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_282_) );
NAND2X1 NAND2X1_112 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_283_) );
NAND3X1 NAND3X1_81 ( .A(_282_), .B(_283_), .C(_278_), .Y(_284_) );
AND2X2 AND2X2_79 ( .A(_284_), .B(_281_), .Y(w_C_46_) );
INVX1 INVX1_155 ( .A(i_add2[46]), .Y(_285_) );
INVX1 INVX1_156 ( .A(i_add1[46]), .Y(_286_) );
NAND2X1 NAND2X1_113 ( .A(_285_), .B(_286_), .Y(_287_) );
NAND3X1 NAND3X1_82 ( .A(_281_), .B(_287_), .C(_284_), .Y(_288_) );
OAI21X1 OAI21X1_68 ( .A(_285_), .B(_286_), .C(_288_), .Y(w_C_47_) );
INVX1 INVX1_157 ( .A(i_add2[47]), .Y(_289_) );
INVX1 INVX1_158 ( .A(i_add1[47]), .Y(_290_) );
OAI21X1 OAI21X1_69 ( .A(i_add2[47]), .B(i_add1[47]), .C(w_C_47_), .Y(_291_) );
OAI21X1 OAI21X1_70 ( .A(_289_), .B(_290_), .C(_291_), .Y(w_C_48_) );
NOR2X1 NOR2X1_92 ( .A(_289_), .B(_290_), .Y(_292_) );
INVX1 INVX1_159 ( .A(_292_), .Y(_293_) );
AND2X2 AND2X2_80 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_294_) );
INVX1 INVX1_160 ( .A(_294_), .Y(_295_) );
NAND3X1 NAND3X1_83 ( .A(_293_), .B(_295_), .C(_291_), .Y(_296_) );
OAI21X1 OAI21X1_71 ( .A(i_add2[48]), .B(i_add1[48]), .C(_296_), .Y(_297_) );
INVX1 INVX1_161 ( .A(_297_), .Y(w_C_49_) );
NAND2X1 NAND2X1_114 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_298_) );
NOR2X1 NOR2X1_93 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_299_) );
OAI21X1 OAI21X1_72 ( .A(_299_), .B(_297_), .C(_298_), .Y(w_C_50_) );
NAND2X1 NAND2X1_115 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_300_) );
INVX1 INVX1_162 ( .A(_299_), .Y(_301_) );
NOR2X1 NOR2X1_94 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_302_) );
INVX1 INVX1_163 ( .A(_302_), .Y(_303_) );
NOR2X1 NOR2X1_95 ( .A(_285_), .B(_286_), .Y(_304_) );
INVX1 INVX1_164 ( .A(_304_), .Y(_305_) );
NAND3X1 NAND3X1_84 ( .A(_305_), .B(_293_), .C(_288_), .Y(_306_) );
NOR2X1 NOR2X1_96 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_307_) );
INVX1 INVX1_165 ( .A(_307_), .Y(_308_) );
NAND3X1 NAND3X1_85 ( .A(_303_), .B(_308_), .C(_306_), .Y(_309_) );
NAND3X1 NAND3X1_86 ( .A(_295_), .B(_298_), .C(_309_), .Y(_310_) );
OR2X2 OR2X2_55 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_311_) );
NAND3X1 NAND3X1_87 ( .A(_301_), .B(_311_), .C(_310_), .Y(_312_) );
NAND2X1 NAND2X1_116 ( .A(_300_), .B(_312_), .Y(w_C_51_) );
OR2X2 OR2X2_56 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_313_) );
NAND2X1 NAND2X1_117 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_314_) );
NAND3X1 NAND3X1_88 ( .A(_300_), .B(_314_), .C(_312_), .Y(_315_) );
AND2X2 AND2X2_81 ( .A(_315_), .B(_313_), .Y(w_C_52_) );
NAND2X1 NAND2X1_118 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_316_) );
OR2X2 OR2X2_57 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_317_) );
NAND3X1 NAND3X1_89 ( .A(_313_), .B(_317_), .C(_315_), .Y(_318_) );
NAND2X1 NAND2X1_119 ( .A(_316_), .B(_318_), .Y(w_C_53_) );
NAND2X1 NAND2X1_120 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_166 ( .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_121 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_122 ( .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_73 ( .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_167 ( .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_123 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_58 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_59 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_90 ( .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_124 ( .A(_4_), .B(_7_), .Y(w_C_3_) );
NAND2X1 NAND2X1_125 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
NAND3X1 NAND3X1_91 ( .A(_4_), .B(_8_), .C(_7_), .Y(_9_) );
OAI21X1 OAI21X1_74 ( .A(i_add2[3]), .B(i_add1[3]), .C(_9_), .Y(_10_) );
INVX1 INVX1_168 ( .A(_10_), .Y(w_C_4_) );
NAND2X1 NAND2X1_126 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
OR2X2 OR2X2_60 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_12_) );
OR2X2 OR2X2_61 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
NAND3X1 NAND3X1_92 ( .A(_12_), .B(_13_), .C(_9_), .Y(_14_) );
NAND2X1 NAND2X1_127 ( .A(_11_), .B(_14_), .Y(w_C_5_) );
NAND2X1 NAND2X1_128 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_15_) );
NAND3X1 NAND3X1_93 ( .A(_11_), .B(_15_), .C(_14_), .Y(_16_) );
OAI21X1 OAI21X1_75 ( .A(i_add2[5]), .B(i_add1[5]), .C(_16_), .Y(_17_) );
INVX1 INVX1_169 ( .A(_17_), .Y(w_C_6_) );
INVX1 INVX1_170 ( .A(i_add2[6]), .Y(_18_) );
INVX1 INVX1_171 ( .A(i_add1[6]), .Y(_19_) );
NOR2X1 NOR2X1_97 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_20_) );
INVX1 INVX1_172 ( .A(_20_), .Y(_21_) );
NOR2X1 NOR2X1_98 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_173 ( .A(_22_), .Y(_23_) );
NAND3X1 NAND3X1_94 ( .A(_21_), .B(_23_), .C(_16_), .Y(_24_) );
OAI21X1 OAI21X1_76 ( .A(_18_), .B(_19_), .C(_24_), .Y(w_C_7_) );
NOR2X1 NOR2X1_99 ( .A(_18_), .B(_19_), .Y(_25_) );
INVX1 INVX1_174 ( .A(_25_), .Y(_26_) );
AND2X2 AND2X2_82 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_27_) );
INVX1 INVX1_175 ( .A(_27_), .Y(_28_) );
NAND3X1 NAND3X1_95 ( .A(_26_), .B(_28_), .C(_24_), .Y(_29_) );
OAI21X1 OAI21X1_77 ( .A(i_add2[7]), .B(i_add1[7]), .C(_29_), .Y(_30_) );
INVX1 INVX1_176 ( .A(_30_), .Y(w_C_8_) );
INVX1 INVX1_177 ( .A(i_add2[8]), .Y(_31_) );
INVX1 INVX1_178 ( .A(i_add1[8]), .Y(_32_) );
NOR2X1 NOR2X1_100 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_33_) );
INVX1 INVX1_179 ( .A(_33_), .Y(_34_) );
NOR2X1 NOR2X1_101 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_35_) );
INVX1 INVX1_180 ( .A(_35_), .Y(_36_) );
NAND3X1 NAND3X1_96 ( .A(_34_), .B(_36_), .C(_29_), .Y(_37_) );
OAI21X1 OAI21X1_78 ( .A(_31_), .B(_32_), .C(_37_), .Y(w_C_9_) );
NOR2X1 NOR2X1_102 ( .A(_31_), .B(_32_), .Y(_38_) );
INVX1 INVX1_181 ( .A(_38_), .Y(_39_) );
AND2X2 AND2X2_83 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_40_) );
INVX1 INVX1_182 ( .A(_40_), .Y(_41_) );
NAND3X1 NAND3X1_97 ( .A(_39_), .B(_41_), .C(_37_), .Y(_42_) );
OAI21X1 OAI21X1_79 ( .A(i_add2[9]), .B(i_add1[9]), .C(_42_), .Y(_43_) );
INVX1 INVX1_183 ( .A(_43_), .Y(w_C_10_) );
INVX1 INVX1_184 ( .A(i_add2[10]), .Y(_44_) );
INVX1 INVX1_185 ( .A(i_add1[10]), .Y(_45_) );
NOR2X1 NOR2X1_103 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_46_) );
INVX1 INVX1_186 ( .A(_46_), .Y(_47_) );
NOR2X1 NOR2X1_104 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_48_) );
INVX1 INVX1_187 ( .A(_48_), .Y(_49_) );
NAND3X1 NAND3X1_98 ( .A(_47_), .B(_49_), .C(_42_), .Y(_50_) );
OAI21X1 OAI21X1_80 ( .A(_44_), .B(_45_), .C(_50_), .Y(w_C_11_) );
NOR2X1 NOR2X1_105 ( .A(_44_), .B(_45_), .Y(_51_) );
INVX1 INVX1_188 ( .A(_51_), .Y(_52_) );
AND2X2 AND2X2_84 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_53_) );
INVX1 INVX1_189 ( .A(_53_), .Y(_54_) );
NAND3X1 NAND3X1_99 ( .A(_52_), .B(_54_), .C(_50_), .Y(_55_) );
OAI21X1 OAI21X1_81 ( .A(i_add2[11]), .B(i_add1[11]), .C(_55_), .Y(_56_) );
INVX1 INVX1_190 ( .A(_56_), .Y(w_C_12_) );
INVX1 INVX1_191 ( .A(i_add2[12]), .Y(_57_) );
INVX1 INVX1_192 ( .A(i_add1[12]), .Y(_58_) );
NOR2X1 NOR2X1_106 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_59_) );
INVX1 INVX1_193 ( .A(_59_), .Y(_60_) );
NOR2X1 NOR2X1_107 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_61_) );
INVX1 INVX1_194 ( .A(_61_), .Y(_62_) );
NAND3X1 NAND3X1_100 ( .A(_60_), .B(_62_), .C(_55_), .Y(_63_) );
OAI21X1 OAI21X1_82 ( .A(_57_), .B(_58_), .C(_63_), .Y(w_C_13_) );
NOR2X1 NOR2X1_108 ( .A(_57_), .B(_58_), .Y(_64_) );
INVX1 INVX1_195 ( .A(_64_), .Y(_65_) );
AND2X2 AND2X2_85 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_66_) );
INVX1 INVX1_196 ( .A(_66_), .Y(_67_) );
NAND3X1 NAND3X1_101 ( .A(_65_), .B(_67_), .C(_63_), .Y(_68_) );
OAI21X1 OAI21X1_83 ( .A(i_add2[13]), .B(i_add1[13]), .C(_68_), .Y(_69_) );
INVX1 INVX1_197 ( .A(_69_), .Y(w_C_14_) );
INVX1 INVX1_198 ( .A(i_add2[14]), .Y(_70_) );
INVX1 INVX1_199 ( .A(i_add1[14]), .Y(_71_) );
NOR2X1 NOR2X1_109 ( .A(_70_), .B(_71_), .Y(_72_) );
INVX1 INVX1_200 ( .A(_72_), .Y(_73_) );
NOR2X1 NOR2X1_110 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_74_) );
INVX1 INVX1_201 ( .A(_74_), .Y(_75_) );
NOR2X1 NOR2X1_111 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_76_) );
INVX1 INVX1_202 ( .A(_76_), .Y(_77_) );
NAND3X1 NAND3X1_102 ( .A(_75_), .B(_77_), .C(_68_), .Y(_78_) );
AND2X2 AND2X2_86 ( .A(_78_), .B(_73_), .Y(_79_) );
INVX1 INVX1_203 ( .A(_79_), .Y(w_C_15_) );
AND2X2 AND2X2_87 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_80_) );
INVX1 INVX1_204 ( .A(_80_), .Y(_81_) );
NAND3X1 NAND3X1_103 ( .A(_73_), .B(_81_), .C(_78_), .Y(_82_) );
OAI21X1 OAI21X1_84 ( .A(i_add2[15]), .B(i_add1[15]), .C(_82_), .Y(_83_) );
INVX1 INVX1_205 ( .A(_83_), .Y(w_C_16_) );
INVX1 INVX1_206 ( .A(i_add2[16]), .Y(_84_) );
INVX1 INVX1_207 ( .A(i_add1[16]), .Y(_85_) );
NOR2X1 NOR2X1_112 ( .A(_84_), .B(_85_), .Y(_86_) );
INVX1 INVX1_208 ( .A(_86_), .Y(_87_) );
NOR2X1 NOR2X1_113 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_88_) );
INVX1 INVX1_209 ( .A(_88_), .Y(_89_) );
NOR2X1 NOR2X1_114 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_90_) );
INVX1 INVX1_210 ( .A(_90_), .Y(_91_) );
NAND3X1 NAND3X1_104 ( .A(_89_), .B(_91_), .C(_82_), .Y(_92_) );
AND2X2 AND2X2_88 ( .A(_92_), .B(_87_), .Y(_93_) );
INVX1 INVX1_211 ( .A(_93_), .Y(w_C_17_) );
AND2X2 AND2X2_89 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_94_) );
INVX1 INVX1_212 ( .A(_94_), .Y(_95_) );
NAND3X1 NAND3X1_105 ( .A(_87_), .B(_95_), .C(_92_), .Y(_96_) );
OAI21X1 OAI21X1_85 ( .A(i_add2[17]), .B(i_add1[17]), .C(_96_), .Y(_97_) );
INVX1 INVX1_213 ( .A(_97_), .Y(w_C_18_) );
INVX1 INVX1_214 ( .A(i_add2[18]), .Y(_98_) );
BUFX2 BUFX2_55 ( .A(w_C_53_), .Y(_319__53_) );
BUFX2 BUFX2_56 ( .A(gnd), .Y(w_C_0_) );
endmodule
