module carry_lookahead_adder_5bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];

OR2X2 OR2X2_1 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_40_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_41_) );
NAND3X1 NAND3X1_1 ( .A(_39_), .B(_41_), .C(_40_), .Y(_42_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_36_) );
AND2X2 AND2X2_1 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_37_) );
OAI21X1 OAI21X1_1 ( .A(_36_), .B(_37_), .C(w_C_2_), .Y(_38_) );
NAND2X1 NAND2X1_2 ( .A(_38_), .B(_42_), .Y(_14__2_) );
INVX1 INVX1_1 ( .A(w_C_3_), .Y(_46_) );
OR2X2 OR2X2_2 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_47_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_48_) );
NAND3X1 NAND3X1_2 ( .A(_46_), .B(_48_), .C(_47_), .Y(_49_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_43_) );
AND2X2 AND2X2_2 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_44_) );
OAI21X1 OAI21X1_2 ( .A(_43_), .B(_44_), .C(w_C_3_), .Y(_45_) );
NAND2X1 NAND2X1_4 ( .A(_45_), .B(_49_), .Y(_14__3_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_2 ( .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_1_) );
OR2X2 OR2X2_3 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_2_) );
OR2X2 OR2X2_4 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_3_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_4_) );
NAND2X1 NAND2X1_8 ( .A(_0_), .B(_4_), .Y(_5_) );
NAND3X1 NAND3X1_3 ( .A(_2_), .B(_3_), .C(_5_), .Y(_6_) );
NAND2X1 NAND2X1_9 ( .A(_1_), .B(_6_), .Y(w_C_3_) );
OR2X2 OR2X2_5 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_7_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
NAND3X1 NAND3X1_4 ( .A(_1_), .B(_8_), .C(_6_), .Y(_9_) );
AND2X2 AND2X2_3 ( .A(_9_), .B(_7_), .Y(w_C_4_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_10_) );
OR2X2 OR2X2_6 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
NAND3X1 NAND3X1_5 ( .A(_7_), .B(_11_), .C(_9_), .Y(_12_) );
NAND2X1 NAND2X1_12 ( .A(_10_), .B(_12_), .Y(w_C_5_) );
OAI21X1 OAI21X1_3 ( .A(i_add2[1]), .B(i_add1[1]), .C(_5_), .Y(_13_) );
INVX1 INVX1_3 ( .A(_13_), .Y(w_C_2_) );
BUFX2 BUFX2_1 ( .A(_14__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_14__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_14__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_14__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_14__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(w_C_5_), .Y(o_result[5]) );
INVX1 INVX1_4 ( .A(w_C_4_), .Y(_18_) );
OR2X2 OR2X2_7 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_19_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_20_) );
NAND3X1 NAND3X1_6 ( .A(_18_), .B(_20_), .C(_19_), .Y(_21_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_15_) );
AND2X2 AND2X2_4 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_16_) );
OAI21X1 OAI21X1_4 ( .A(_15_), .B(_16_), .C(w_C_4_), .Y(_17_) );
NAND2X1 NAND2X1_14 ( .A(_17_), .B(_21_), .Y(_14__4_) );
INVX1 INVX1_5 ( .A(1'b0), .Y(_25_) );
OR2X2 OR2X2_8 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_26_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_27_) );
NAND3X1 NAND3X1_7 ( .A(_25_), .B(_27_), .C(_26_), .Y(_28_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_22_) );
AND2X2 AND2X2_5 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_23_) );
OAI21X1 OAI21X1_5 ( .A(_22_), .B(_23_), .C(1'b0), .Y(_24_) );
NAND2X1 NAND2X1_16 ( .A(_24_), .B(_28_), .Y(_14__0_) );
INVX1 INVX1_6 ( .A(w_C_1_), .Y(_32_) );
OR2X2 OR2X2_9 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_33_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_34_) );
NAND3X1 NAND3X1_8 ( .A(_32_), .B(_34_), .C(_33_), .Y(_35_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_29_) );
AND2X2 AND2X2_6 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_30_) );
OAI21X1 OAI21X1_6 ( .A(_29_), .B(_30_), .C(w_C_1_), .Y(_31_) );
NAND2X1 NAND2X1_18 ( .A(_31_), .B(_35_), .Y(_14__1_) );
INVX1 INVX1_7 ( .A(w_C_2_), .Y(_39_) );
BUFX2 BUFX2_7 ( .A(w_C_5_), .Y(_14__5_) );
BUFX2 BUFX2_8 ( .A(1'b0), .Y(w_C_0_) );
endmodule
