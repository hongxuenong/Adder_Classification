module csa_60bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term1[45], i_add_term1[46], i_add_term1[47], i_add_term1[48], i_add_term1[49], i_add_term1[50], i_add_term1[51], i_add_term1[52], i_add_term1[53], i_add_term1[54], i_add_term1[55], i_add_term1[56], i_add_term1[57], i_add_term1[58], i_add_term1[59], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], i_add_term2[45], i_add_term2[46], i_add_term2[47], i_add_term2[48], i_add_term2[49], i_add_term2[50], i_add_term2[51], i_add_term2[52], i_add_term2[53], i_add_term2[54], i_add_term2[55], i_add_term2[56], i_add_term2[57], i_add_term2[58], i_add_term2[59], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], sum[45], sum[46], sum[47], sum[48], sum[49], sum[50], sum[51], sum[52], sum[53], sum[54], sum[55], sum[56], sum[57], sum[58], sum[59], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term1[45];
input i_add_term1[46];
input i_add_term1[47];
input i_add_term1[48];
input i_add_term1[49];
input i_add_term1[50];
input i_add_term1[51];
input i_add_term1[52];
input i_add_term1[53];
input i_add_term1[54];
input i_add_term1[55];
input i_add_term1[56];
input i_add_term1[57];
input i_add_term1[58];
input i_add_term1[59];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
input i_add_term2[45];
input i_add_term2[46];
input i_add_term2[47];
input i_add_term2[48];
input i_add_term2[49];
input i_add_term2[50];
input i_add_term2[51];
input i_add_term2[52];
input i_add_term2[53];
input i_add_term2[54];
input i_add_term2[55];
input i_add_term2[56];
input i_add_term2[57];
input i_add_term2[58];
input i_add_term2[59];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output sum[45];
output sum[46];
output sum[47];
output sum[48];
output sum[49];
output sum[50];
output sum[51];
output sum[52];
output sum[53];
output sum[54];
output sum[55];
output sum[56];
output sum[57];
output sum[58];
output sum[59];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_14_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .A(_0__54_), .Y(sum[54]) );
BUFX2 BUFX2_57 ( .A(_0__55_), .Y(sum[55]) );
BUFX2 BUFX2_58 ( .A(_0__56_), .Y(sum[56]) );
BUFX2 BUFX2_59 ( .A(_0__57_), .Y(sum[57]) );
BUFX2 BUFX2_60 ( .A(_0__58_), .Y(sum[58]) );
BUFX2 BUFX2_61 ( .A(_0__59_), .Y(sum[59]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_85_) );
NAND2X1 NAND2X1_1 ( .A(_2_), .B(rca_inst_cout), .Y(_86_) );
OAI21X1 OAI21X1_1 ( .A(rca_inst_cout), .B(_85_), .C(_86_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3__0_), .Y(_87_) );
NAND2X1 NAND2X1_2 ( .A(_4__0_), .B(rca_inst_cout), .Y(_88_) );
OAI21X1 OAI21X1_2 ( .A(rca_inst_cout), .B(_87_), .C(_88_), .Y(_0__4_) );
INVX1 INVX1_3 ( .A(_3__1_), .Y(_89_) );
NAND2X1 NAND2X1_3 ( .A(rca_inst_cout), .B(_4__1_), .Y(_90_) );
OAI21X1 OAI21X1_3 ( .A(rca_inst_cout), .B(_89_), .C(_90_), .Y(_0__5_) );
INVX1 INVX1_4 ( .A(_3__2_), .Y(_91_) );
NAND2X1 NAND2X1_4 ( .A(rca_inst_cout), .B(_4__2_), .Y(_92_) );
OAI21X1 OAI21X1_4 ( .A(rca_inst_cout), .B(_91_), .C(_92_), .Y(_0__6_) );
INVX1 INVX1_5 ( .A(_3__3_), .Y(_93_) );
NAND2X1 NAND2X1_5 ( .A(rca_inst_cout), .B(_4__3_), .Y(_94_) );
OAI21X1 OAI21X1_5 ( .A(rca_inst_cout), .B(_93_), .C(_94_), .Y(_0__7_) );
INVX1 INVX1_6 ( .A(1'b0), .Y(_98_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_99_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_100_) );
NAND3X1 NAND3X1_1 ( .A(_98_), .B(_100_), .C(_99_), .Y(_101_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_95_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_96_) );
OAI21X1 OAI21X1_6 ( .A(_95_), .B(_96_), .C(1'b0), .Y(_97_) );
NAND2X1 NAND2X1_7 ( .A(_97_), .B(_101_), .Y(_3__0_) );
OAI21X1 OAI21X1_7 ( .A(_98_), .B(_95_), .C(_100_), .Y(_5__1_) );
INVX1 INVX1_7 ( .A(_5__3_), .Y(_105_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_106_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_107_) );
NAND3X1 NAND3X1_2 ( .A(_105_), .B(_107_), .C(_106_), .Y(_108_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_102_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_103_) );
OAI21X1 OAI21X1_8 ( .A(_102_), .B(_103_), .C(_5__3_), .Y(_104_) );
NAND2X1 NAND2X1_9 ( .A(_104_), .B(_108_), .Y(_3__3_) );
OAI21X1 OAI21X1_9 ( .A(_105_), .B(_102_), .C(_107_), .Y(_1_) );
INVX1 INVX1_8 ( .A(_5__1_), .Y(_112_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_113_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_114_) );
NAND3X1 NAND3X1_3 ( .A(_112_), .B(_114_), .C(_113_), .Y(_115_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_109_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_110_) );
OAI21X1 OAI21X1_10 ( .A(_109_), .B(_110_), .C(_5__1_), .Y(_111_) );
NAND2X1 NAND2X1_11 ( .A(_111_), .B(_115_), .Y(_3__1_) );
OAI21X1 OAI21X1_11 ( .A(_112_), .B(_109_), .C(_114_), .Y(_5__2_) );
INVX1 INVX1_9 ( .A(_5__2_), .Y(_119_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_120_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_121_) );
NAND3X1 NAND3X1_4 ( .A(_119_), .B(_121_), .C(_120_), .Y(_122_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_116_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_117_) );
OAI21X1 OAI21X1_12 ( .A(_116_), .B(_117_), .C(_5__2_), .Y(_118_) );
NAND2X1 NAND2X1_13 ( .A(_118_), .B(_122_), .Y(_3__2_) );
OAI21X1 OAI21X1_13 ( .A(_119_), .B(_116_), .C(_121_), .Y(_5__3_) );
INVX1 INVX1_10 ( .A(1'b1), .Y(_126_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_127_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_128_) );
NAND3X1 NAND3X1_5 ( .A(_126_), .B(_128_), .C(_127_), .Y(_129_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_123_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_124_) );
OAI21X1 OAI21X1_14 ( .A(_123_), .B(_124_), .C(1'b1), .Y(_125_) );
NAND2X1 NAND2X1_15 ( .A(_125_), .B(_129_), .Y(_4__0_) );
OAI21X1 OAI21X1_15 ( .A(_126_), .B(_123_), .C(_128_), .Y(_6__1_) );
INVX1 INVX1_11 ( .A(_6__3_), .Y(_133_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_134_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_135_) );
NAND3X1 NAND3X1_6 ( .A(_133_), .B(_135_), .C(_134_), .Y(_136_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_130_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_131_) );
OAI21X1 OAI21X1_16 ( .A(_130_), .B(_131_), .C(_6__3_), .Y(_132_) );
NAND2X1 NAND2X1_17 ( .A(_132_), .B(_136_), .Y(_4__3_) );
OAI21X1 OAI21X1_17 ( .A(_133_), .B(_130_), .C(_135_), .Y(_2_) );
INVX1 INVX1_12 ( .A(_6__1_), .Y(_140_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_141_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_142_) );
NAND3X1 NAND3X1_7 ( .A(_140_), .B(_142_), .C(_141_), .Y(_143_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_137_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_138_) );
OAI21X1 OAI21X1_18 ( .A(_137_), .B(_138_), .C(_6__1_), .Y(_139_) );
NAND2X1 NAND2X1_19 ( .A(_139_), .B(_143_), .Y(_4__1_) );
OAI21X1 OAI21X1_19 ( .A(_140_), .B(_137_), .C(_142_), .Y(_6__2_) );
INVX1 INVX1_13 ( .A(_6__2_), .Y(_147_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_148_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_149_) );
NAND3X1 NAND3X1_8 ( .A(_147_), .B(_149_), .C(_148_), .Y(_150_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_144_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_145_) );
OAI21X1 OAI21X1_20 ( .A(_144_), .B(_145_), .C(_6__2_), .Y(_146_) );
NAND2X1 NAND2X1_21 ( .A(_146_), .B(_150_), .Y(_4__2_) );
OAI21X1 OAI21X1_21 ( .A(_147_), .B(_144_), .C(_149_), .Y(_6__3_) );
INVX1 INVX1_14 ( .A(_7_), .Y(_151_) );
NAND2X1 NAND2X1_22 ( .A(_8_), .B(w_cout_1_), .Y(_152_) );
OAI21X1 OAI21X1_22 ( .A(w_cout_1_), .B(_151_), .C(_152_), .Y(w_cout_2_) );
INVX1 INVX1_15 ( .A(_9__0_), .Y(_153_) );
NAND2X1 NAND2X1_23 ( .A(_10__0_), .B(w_cout_1_), .Y(_154_) );
OAI21X1 OAI21X1_23 ( .A(w_cout_1_), .B(_153_), .C(_154_), .Y(_0__8_) );
INVX1 INVX1_16 ( .A(_9__1_), .Y(_155_) );
NAND2X1 NAND2X1_24 ( .A(w_cout_1_), .B(_10__1_), .Y(_156_) );
OAI21X1 OAI21X1_24 ( .A(w_cout_1_), .B(_155_), .C(_156_), .Y(_0__9_) );
INVX1 INVX1_17 ( .A(_9__2_), .Y(_157_) );
NAND2X1 NAND2X1_25 ( .A(w_cout_1_), .B(_10__2_), .Y(_158_) );
OAI21X1 OAI21X1_25 ( .A(w_cout_1_), .B(_157_), .C(_158_), .Y(_0__10_) );
INVX1 INVX1_18 ( .A(_9__3_), .Y(_159_) );
NAND2X1 NAND2X1_26 ( .A(w_cout_1_), .B(_10__3_), .Y(_160_) );
OAI21X1 OAI21X1_26 ( .A(w_cout_1_), .B(_159_), .C(_160_), .Y(_0__11_) );
INVX1 INVX1_19 ( .A(1'b0), .Y(_164_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_165_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_166_) );
NAND3X1 NAND3X1_9 ( .A(_164_), .B(_166_), .C(_165_), .Y(_167_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_161_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_162_) );
OAI21X1 OAI21X1_27 ( .A(_161_), .B(_162_), .C(1'b0), .Y(_163_) );
NAND2X1 NAND2X1_28 ( .A(_163_), .B(_167_), .Y(_9__0_) );
OAI21X1 OAI21X1_28 ( .A(_164_), .B(_161_), .C(_166_), .Y(_11__1_) );
INVX1 INVX1_20 ( .A(_11__3_), .Y(_171_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_172_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_173_) );
NAND3X1 NAND3X1_10 ( .A(_171_), .B(_173_), .C(_172_), .Y(_174_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_168_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_169_) );
OAI21X1 OAI21X1_29 ( .A(_168_), .B(_169_), .C(_11__3_), .Y(_170_) );
NAND2X1 NAND2X1_30 ( .A(_170_), .B(_174_), .Y(_9__3_) );
OAI21X1 OAI21X1_30 ( .A(_171_), .B(_168_), .C(_173_), .Y(_7_) );
INVX1 INVX1_21 ( .A(_11__1_), .Y(_178_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_179_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_180_) );
NAND3X1 NAND3X1_11 ( .A(_178_), .B(_180_), .C(_179_), .Y(_181_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_175_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_176_) );
OAI21X1 OAI21X1_31 ( .A(_175_), .B(_176_), .C(_11__1_), .Y(_177_) );
NAND2X1 NAND2X1_32 ( .A(_177_), .B(_181_), .Y(_9__1_) );
OAI21X1 OAI21X1_32 ( .A(_178_), .B(_175_), .C(_180_), .Y(_11__2_) );
INVX1 INVX1_22 ( .A(_11__2_), .Y(_185_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_186_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_187_) );
NAND3X1 NAND3X1_12 ( .A(_185_), .B(_187_), .C(_186_), .Y(_188_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_182_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_183_) );
OAI21X1 OAI21X1_33 ( .A(_182_), .B(_183_), .C(_11__2_), .Y(_184_) );
NAND2X1 NAND2X1_34 ( .A(_184_), .B(_188_), .Y(_9__2_) );
OAI21X1 OAI21X1_34 ( .A(_185_), .B(_182_), .C(_187_), .Y(_11__3_) );
INVX1 INVX1_23 ( .A(1'b1), .Y(_192_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_193_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_194_) );
NAND3X1 NAND3X1_13 ( .A(_192_), .B(_194_), .C(_193_), .Y(_195_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_189_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_190_) );
OAI21X1 OAI21X1_35 ( .A(_189_), .B(_190_), .C(1'b1), .Y(_191_) );
NAND2X1 NAND2X1_36 ( .A(_191_), .B(_195_), .Y(_10__0_) );
OAI21X1 OAI21X1_36 ( .A(_192_), .B(_189_), .C(_194_), .Y(_12__1_) );
INVX1 INVX1_24 ( .A(_12__3_), .Y(_199_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_200_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_201_) );
NAND3X1 NAND3X1_14 ( .A(_199_), .B(_201_), .C(_200_), .Y(_202_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_196_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_197_) );
OAI21X1 OAI21X1_37 ( .A(_196_), .B(_197_), .C(_12__3_), .Y(_198_) );
NAND2X1 NAND2X1_38 ( .A(_198_), .B(_202_), .Y(_10__3_) );
OAI21X1 OAI21X1_38 ( .A(_199_), .B(_196_), .C(_201_), .Y(_8_) );
INVX1 INVX1_25 ( .A(_12__1_), .Y(_206_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_207_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_208_) );
NAND3X1 NAND3X1_15 ( .A(_206_), .B(_208_), .C(_207_), .Y(_209_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_203_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_204_) );
OAI21X1 OAI21X1_39 ( .A(_203_), .B(_204_), .C(_12__1_), .Y(_205_) );
NAND2X1 NAND2X1_40 ( .A(_205_), .B(_209_), .Y(_10__1_) );
OAI21X1 OAI21X1_40 ( .A(_206_), .B(_203_), .C(_208_), .Y(_12__2_) );
INVX1 INVX1_26 ( .A(_12__2_), .Y(_213_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_214_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_215_) );
NAND3X1 NAND3X1_16 ( .A(_213_), .B(_215_), .C(_214_), .Y(_216_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_210_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_211_) );
OAI21X1 OAI21X1_41 ( .A(_210_), .B(_211_), .C(_12__2_), .Y(_212_) );
NAND2X1 NAND2X1_42 ( .A(_212_), .B(_216_), .Y(_10__2_) );
OAI21X1 OAI21X1_42 ( .A(_213_), .B(_210_), .C(_215_), .Y(_12__3_) );
INVX1 INVX1_27 ( .A(_13_), .Y(_217_) );
NAND2X1 NAND2X1_43 ( .A(_14_), .B(w_cout_2_), .Y(_218_) );
OAI21X1 OAI21X1_43 ( .A(w_cout_2_), .B(_217_), .C(_218_), .Y(w_cout_3_) );
INVX1 INVX1_28 ( .A(_15__0_), .Y(_219_) );
NAND2X1 NAND2X1_44 ( .A(_16__0_), .B(w_cout_2_), .Y(_220_) );
OAI21X1 OAI21X1_44 ( .A(w_cout_2_), .B(_219_), .C(_220_), .Y(_0__12_) );
INVX1 INVX1_29 ( .A(_15__1_), .Y(_221_) );
NAND2X1 NAND2X1_45 ( .A(w_cout_2_), .B(_16__1_), .Y(_222_) );
OAI21X1 OAI21X1_45 ( .A(w_cout_2_), .B(_221_), .C(_222_), .Y(_0__13_) );
INVX1 INVX1_30 ( .A(_15__2_), .Y(_223_) );
NAND2X1 NAND2X1_46 ( .A(w_cout_2_), .B(_16__2_), .Y(_224_) );
OAI21X1 OAI21X1_46 ( .A(w_cout_2_), .B(_223_), .C(_224_), .Y(_0__14_) );
INVX1 INVX1_31 ( .A(_15__3_), .Y(_225_) );
NAND2X1 NAND2X1_47 ( .A(w_cout_2_), .B(_16__3_), .Y(_226_) );
OAI21X1 OAI21X1_47 ( .A(w_cout_2_), .B(_225_), .C(_226_), .Y(_0__15_) );
INVX1 INVX1_32 ( .A(1'b0), .Y(_230_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_231_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_232_) );
NAND3X1 NAND3X1_17 ( .A(_230_), .B(_232_), .C(_231_), .Y(_233_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_227_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_228_) );
OAI21X1 OAI21X1_48 ( .A(_227_), .B(_228_), .C(1'b0), .Y(_229_) );
NAND2X1 NAND2X1_49 ( .A(_229_), .B(_233_), .Y(_15__0_) );
OAI21X1 OAI21X1_49 ( .A(_230_), .B(_227_), .C(_232_), .Y(_17__1_) );
INVX1 INVX1_33 ( .A(_17__3_), .Y(_237_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_238_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_239_) );
NAND3X1 NAND3X1_18 ( .A(_237_), .B(_239_), .C(_238_), .Y(_240_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_234_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_235_) );
OAI21X1 OAI21X1_50 ( .A(_234_), .B(_235_), .C(_17__3_), .Y(_236_) );
NAND2X1 NAND2X1_51 ( .A(_236_), .B(_240_), .Y(_15__3_) );
OAI21X1 OAI21X1_51 ( .A(_237_), .B(_234_), .C(_239_), .Y(_13_) );
INVX1 INVX1_34 ( .A(_17__1_), .Y(_244_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_245_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_246_) );
NAND3X1 NAND3X1_19 ( .A(_244_), .B(_246_), .C(_245_), .Y(_247_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_241_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_242_) );
OAI21X1 OAI21X1_52 ( .A(_241_), .B(_242_), .C(_17__1_), .Y(_243_) );
NAND2X1 NAND2X1_53 ( .A(_243_), .B(_247_), .Y(_15__1_) );
OAI21X1 OAI21X1_53 ( .A(_244_), .B(_241_), .C(_246_), .Y(_17__2_) );
INVX1 INVX1_35 ( .A(_17__2_), .Y(_251_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_252_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_253_) );
NAND3X1 NAND3X1_20 ( .A(_251_), .B(_253_), .C(_252_), .Y(_254_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_248_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_249_) );
OAI21X1 OAI21X1_54 ( .A(_248_), .B(_249_), .C(_17__2_), .Y(_250_) );
NAND2X1 NAND2X1_55 ( .A(_250_), .B(_254_), .Y(_15__2_) );
OAI21X1 OAI21X1_55 ( .A(_251_), .B(_248_), .C(_253_), .Y(_17__3_) );
INVX1 INVX1_36 ( .A(1'b1), .Y(_258_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_259_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_260_) );
NAND3X1 NAND3X1_21 ( .A(_258_), .B(_260_), .C(_259_), .Y(_261_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_255_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_256_) );
OAI21X1 OAI21X1_56 ( .A(_255_), .B(_256_), .C(1'b1), .Y(_257_) );
NAND2X1 NAND2X1_57 ( .A(_257_), .B(_261_), .Y(_16__0_) );
OAI21X1 OAI21X1_57 ( .A(_258_), .B(_255_), .C(_260_), .Y(_18__1_) );
INVX1 INVX1_37 ( .A(_18__3_), .Y(_265_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_266_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_267_) );
NAND3X1 NAND3X1_22 ( .A(_265_), .B(_267_), .C(_266_), .Y(_268_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_262_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_263_) );
OAI21X1 OAI21X1_58 ( .A(_262_), .B(_263_), .C(_18__3_), .Y(_264_) );
NAND2X1 NAND2X1_59 ( .A(_264_), .B(_268_), .Y(_16__3_) );
OAI21X1 OAI21X1_59 ( .A(_265_), .B(_262_), .C(_267_), .Y(_14_) );
INVX1 INVX1_38 ( .A(_18__1_), .Y(_272_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_273_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_274_) );
NAND3X1 NAND3X1_23 ( .A(_272_), .B(_274_), .C(_273_), .Y(_275_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_269_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_270_) );
OAI21X1 OAI21X1_60 ( .A(_269_), .B(_270_), .C(_18__1_), .Y(_271_) );
NAND2X1 NAND2X1_61 ( .A(_271_), .B(_275_), .Y(_16__1_) );
OAI21X1 OAI21X1_61 ( .A(_272_), .B(_269_), .C(_274_), .Y(_18__2_) );
INVX1 INVX1_39 ( .A(_18__2_), .Y(_279_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_280_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_281_) );
NAND3X1 NAND3X1_24 ( .A(_279_), .B(_281_), .C(_280_), .Y(_282_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_276_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_277_) );
OAI21X1 OAI21X1_62 ( .A(_276_), .B(_277_), .C(_18__2_), .Y(_278_) );
NAND2X1 NAND2X1_63 ( .A(_278_), .B(_282_), .Y(_16__2_) );
OAI21X1 OAI21X1_63 ( .A(_279_), .B(_276_), .C(_281_), .Y(_18__3_) );
INVX1 INVX1_40 ( .A(_19_), .Y(_283_) );
NAND2X1 NAND2X1_64 ( .A(_20_), .B(w_cout_3_), .Y(_284_) );
OAI21X1 OAI21X1_64 ( .A(w_cout_3_), .B(_283_), .C(_284_), .Y(w_cout_4_) );
INVX1 INVX1_41 ( .A(_21__0_), .Y(_285_) );
NAND2X1 NAND2X1_65 ( .A(_22__0_), .B(w_cout_3_), .Y(_286_) );
OAI21X1 OAI21X1_65 ( .A(w_cout_3_), .B(_285_), .C(_286_), .Y(_0__16_) );
INVX1 INVX1_42 ( .A(_21__1_), .Y(_287_) );
NAND2X1 NAND2X1_66 ( .A(w_cout_3_), .B(_22__1_), .Y(_288_) );
OAI21X1 OAI21X1_66 ( .A(w_cout_3_), .B(_287_), .C(_288_), .Y(_0__17_) );
INVX1 INVX1_43 ( .A(_21__2_), .Y(_289_) );
NAND2X1 NAND2X1_67 ( .A(w_cout_3_), .B(_22__2_), .Y(_290_) );
OAI21X1 OAI21X1_67 ( .A(w_cout_3_), .B(_289_), .C(_290_), .Y(_0__18_) );
INVX1 INVX1_44 ( .A(_21__3_), .Y(_291_) );
NAND2X1 NAND2X1_68 ( .A(w_cout_3_), .B(_22__3_), .Y(_292_) );
OAI21X1 OAI21X1_68 ( .A(w_cout_3_), .B(_291_), .C(_292_), .Y(_0__19_) );
INVX1 INVX1_45 ( .A(1'b0), .Y(_296_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_297_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_298_) );
NAND3X1 NAND3X1_25 ( .A(_296_), .B(_298_), .C(_297_), .Y(_299_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_293_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_294_) );
OAI21X1 OAI21X1_69 ( .A(_293_), .B(_294_), .C(1'b0), .Y(_295_) );
NAND2X1 NAND2X1_70 ( .A(_295_), .B(_299_), .Y(_21__0_) );
OAI21X1 OAI21X1_70 ( .A(_296_), .B(_293_), .C(_298_), .Y(_23__1_) );
INVX1 INVX1_46 ( .A(_23__3_), .Y(_303_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_304_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_305_) );
NAND3X1 NAND3X1_26 ( .A(_303_), .B(_305_), .C(_304_), .Y(_306_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_300_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_301_) );
OAI21X1 OAI21X1_71 ( .A(_300_), .B(_301_), .C(_23__3_), .Y(_302_) );
NAND2X1 NAND2X1_72 ( .A(_302_), .B(_306_), .Y(_21__3_) );
OAI21X1 OAI21X1_72 ( .A(_303_), .B(_300_), .C(_305_), .Y(_19_) );
INVX1 INVX1_47 ( .A(_23__1_), .Y(_310_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_311_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_312_) );
NAND3X1 NAND3X1_27 ( .A(_310_), .B(_312_), .C(_311_), .Y(_313_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_307_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_308_) );
OAI21X1 OAI21X1_73 ( .A(_307_), .B(_308_), .C(_23__1_), .Y(_309_) );
NAND2X1 NAND2X1_74 ( .A(_309_), .B(_313_), .Y(_21__1_) );
OAI21X1 OAI21X1_74 ( .A(_310_), .B(_307_), .C(_312_), .Y(_23__2_) );
INVX1 INVX1_48 ( .A(_23__2_), .Y(_317_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_318_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_319_) );
NAND3X1 NAND3X1_28 ( .A(_317_), .B(_319_), .C(_318_), .Y(_320_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_314_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_315_) );
OAI21X1 OAI21X1_75 ( .A(_314_), .B(_315_), .C(_23__2_), .Y(_316_) );
NAND2X1 NAND2X1_76 ( .A(_316_), .B(_320_), .Y(_21__2_) );
OAI21X1 OAI21X1_76 ( .A(_317_), .B(_314_), .C(_319_), .Y(_23__3_) );
INVX1 INVX1_49 ( .A(1'b1), .Y(_324_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_325_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_326_) );
NAND3X1 NAND3X1_29 ( .A(_324_), .B(_326_), .C(_325_), .Y(_327_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_321_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_322_) );
OAI21X1 OAI21X1_77 ( .A(_321_), .B(_322_), .C(1'b1), .Y(_323_) );
NAND2X1 NAND2X1_78 ( .A(_323_), .B(_327_), .Y(_22__0_) );
OAI21X1 OAI21X1_78 ( .A(_324_), .B(_321_), .C(_326_), .Y(_24__1_) );
INVX1 INVX1_50 ( .A(_24__3_), .Y(_331_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_332_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_333_) );
NAND3X1 NAND3X1_30 ( .A(_331_), .B(_333_), .C(_332_), .Y(_334_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_328_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_329_) );
OAI21X1 OAI21X1_79 ( .A(_328_), .B(_329_), .C(_24__3_), .Y(_330_) );
NAND2X1 NAND2X1_80 ( .A(_330_), .B(_334_), .Y(_22__3_) );
OAI21X1 OAI21X1_80 ( .A(_331_), .B(_328_), .C(_333_), .Y(_20_) );
INVX1 INVX1_51 ( .A(_24__1_), .Y(_338_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_339_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_340_) );
NAND3X1 NAND3X1_31 ( .A(_338_), .B(_340_), .C(_339_), .Y(_341_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_335_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_336_) );
OAI21X1 OAI21X1_81 ( .A(_335_), .B(_336_), .C(_24__1_), .Y(_337_) );
NAND2X1 NAND2X1_82 ( .A(_337_), .B(_341_), .Y(_22__1_) );
OAI21X1 OAI21X1_82 ( .A(_338_), .B(_335_), .C(_340_), .Y(_24__2_) );
INVX1 INVX1_52 ( .A(_24__2_), .Y(_345_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_346_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_347_) );
NAND3X1 NAND3X1_32 ( .A(_345_), .B(_347_), .C(_346_), .Y(_348_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_342_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_343_) );
OAI21X1 OAI21X1_83 ( .A(_342_), .B(_343_), .C(_24__2_), .Y(_344_) );
NAND2X1 NAND2X1_84 ( .A(_344_), .B(_348_), .Y(_22__2_) );
OAI21X1 OAI21X1_84 ( .A(_345_), .B(_342_), .C(_347_), .Y(_24__3_) );
INVX1 INVX1_53 ( .A(_25_), .Y(_349_) );
NAND2X1 NAND2X1_85 ( .A(_26_), .B(w_cout_4_), .Y(_350_) );
OAI21X1 OAI21X1_85 ( .A(w_cout_4_), .B(_349_), .C(_350_), .Y(w_cout_5_) );
INVX1 INVX1_54 ( .A(_27__0_), .Y(_351_) );
NAND2X1 NAND2X1_86 ( .A(_28__0_), .B(w_cout_4_), .Y(_352_) );
OAI21X1 OAI21X1_86 ( .A(w_cout_4_), .B(_351_), .C(_352_), .Y(_0__20_) );
INVX1 INVX1_55 ( .A(_27__1_), .Y(_353_) );
NAND2X1 NAND2X1_87 ( .A(w_cout_4_), .B(_28__1_), .Y(_354_) );
OAI21X1 OAI21X1_87 ( .A(w_cout_4_), .B(_353_), .C(_354_), .Y(_0__21_) );
INVX1 INVX1_56 ( .A(_27__2_), .Y(_355_) );
NAND2X1 NAND2X1_88 ( .A(w_cout_4_), .B(_28__2_), .Y(_356_) );
OAI21X1 OAI21X1_88 ( .A(w_cout_4_), .B(_355_), .C(_356_), .Y(_0__22_) );
INVX1 INVX1_57 ( .A(_27__3_), .Y(_357_) );
NAND2X1 NAND2X1_89 ( .A(w_cout_4_), .B(_28__3_), .Y(_358_) );
OAI21X1 OAI21X1_89 ( .A(w_cout_4_), .B(_357_), .C(_358_), .Y(_0__23_) );
INVX1 INVX1_58 ( .A(1'b0), .Y(_362_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_363_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_364_) );
NAND3X1 NAND3X1_33 ( .A(_362_), .B(_364_), .C(_363_), .Y(_365_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_359_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_360_) );
OAI21X1 OAI21X1_90 ( .A(_359_), .B(_360_), .C(1'b0), .Y(_361_) );
NAND2X1 NAND2X1_91 ( .A(_361_), .B(_365_), .Y(_27__0_) );
OAI21X1 OAI21X1_91 ( .A(_362_), .B(_359_), .C(_364_), .Y(_29__1_) );
INVX1 INVX1_59 ( .A(_29__3_), .Y(_369_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_370_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_371_) );
NAND3X1 NAND3X1_34 ( .A(_369_), .B(_371_), .C(_370_), .Y(_372_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_366_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_367_) );
OAI21X1 OAI21X1_92 ( .A(_366_), .B(_367_), .C(_29__3_), .Y(_368_) );
NAND2X1 NAND2X1_93 ( .A(_368_), .B(_372_), .Y(_27__3_) );
OAI21X1 OAI21X1_93 ( .A(_369_), .B(_366_), .C(_371_), .Y(_25_) );
INVX1 INVX1_60 ( .A(_29__1_), .Y(_376_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_377_) );
NAND2X1 NAND2X1_94 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_378_) );
NAND3X1 NAND3X1_35 ( .A(_376_), .B(_378_), .C(_377_), .Y(_379_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_373_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_374_) );
OAI21X1 OAI21X1_94 ( .A(_373_), .B(_374_), .C(_29__1_), .Y(_375_) );
NAND2X1 NAND2X1_95 ( .A(_375_), .B(_379_), .Y(_27__1_) );
OAI21X1 OAI21X1_95 ( .A(_376_), .B(_373_), .C(_378_), .Y(_29__2_) );
INVX1 INVX1_61 ( .A(_29__2_), .Y(_383_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_384_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_385_) );
NAND3X1 NAND3X1_36 ( .A(_383_), .B(_385_), .C(_384_), .Y(_386_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_380_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_381_) );
OAI21X1 OAI21X1_96 ( .A(_380_), .B(_381_), .C(_29__2_), .Y(_382_) );
NAND2X1 NAND2X1_97 ( .A(_382_), .B(_386_), .Y(_27__2_) );
OAI21X1 OAI21X1_97 ( .A(_383_), .B(_380_), .C(_385_), .Y(_29__3_) );
INVX1 INVX1_62 ( .A(1'b1), .Y(_390_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_391_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_392_) );
NAND3X1 NAND3X1_37 ( .A(_390_), .B(_392_), .C(_391_), .Y(_393_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_387_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_388_) );
OAI21X1 OAI21X1_98 ( .A(_387_), .B(_388_), .C(1'b1), .Y(_389_) );
NAND2X1 NAND2X1_99 ( .A(_389_), .B(_393_), .Y(_28__0_) );
OAI21X1 OAI21X1_99 ( .A(_390_), .B(_387_), .C(_392_), .Y(_30__1_) );
INVX1 INVX1_63 ( .A(_30__3_), .Y(_397_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_398_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_399_) );
NAND3X1 NAND3X1_38 ( .A(_397_), .B(_399_), .C(_398_), .Y(_400_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_394_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_395_) );
OAI21X1 OAI21X1_100 ( .A(_394_), .B(_395_), .C(_30__3_), .Y(_396_) );
NAND2X1 NAND2X1_101 ( .A(_396_), .B(_400_), .Y(_28__3_) );
OAI21X1 OAI21X1_101 ( .A(_397_), .B(_394_), .C(_399_), .Y(_26_) );
INVX1 INVX1_64 ( .A(_30__1_), .Y(_404_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_405_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_406_) );
NAND3X1 NAND3X1_39 ( .A(_404_), .B(_406_), .C(_405_), .Y(_407_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_401_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_402_) );
OAI21X1 OAI21X1_102 ( .A(_401_), .B(_402_), .C(_30__1_), .Y(_403_) );
NAND2X1 NAND2X1_103 ( .A(_403_), .B(_407_), .Y(_28__1_) );
OAI21X1 OAI21X1_103 ( .A(_404_), .B(_401_), .C(_406_), .Y(_30__2_) );
INVX1 INVX1_65 ( .A(_30__2_), .Y(_411_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_412_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_413_) );
NAND3X1 NAND3X1_40 ( .A(_411_), .B(_413_), .C(_412_), .Y(_414_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_408_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_409_) );
OAI21X1 OAI21X1_104 ( .A(_408_), .B(_409_), .C(_30__2_), .Y(_410_) );
NAND2X1 NAND2X1_105 ( .A(_410_), .B(_414_), .Y(_28__2_) );
OAI21X1 OAI21X1_105 ( .A(_411_), .B(_408_), .C(_413_), .Y(_30__3_) );
INVX1 INVX1_66 ( .A(_31_), .Y(_415_) );
NAND2X1 NAND2X1_106 ( .A(_32_), .B(w_cout_5_), .Y(_416_) );
OAI21X1 OAI21X1_106 ( .A(w_cout_5_), .B(_415_), .C(_416_), .Y(w_cout_6_) );
INVX1 INVX1_67 ( .A(_33__0_), .Y(_417_) );
NAND2X1 NAND2X1_107 ( .A(_34__0_), .B(w_cout_5_), .Y(_418_) );
OAI21X1 OAI21X1_107 ( .A(w_cout_5_), .B(_417_), .C(_418_), .Y(_0__24_) );
INVX1 INVX1_68 ( .A(_33__1_), .Y(_419_) );
NAND2X1 NAND2X1_108 ( .A(w_cout_5_), .B(_34__1_), .Y(_420_) );
OAI21X1 OAI21X1_108 ( .A(w_cout_5_), .B(_419_), .C(_420_), .Y(_0__25_) );
INVX1 INVX1_69 ( .A(_33__2_), .Y(_421_) );
NAND2X1 NAND2X1_109 ( .A(w_cout_5_), .B(_34__2_), .Y(_422_) );
OAI21X1 OAI21X1_109 ( .A(w_cout_5_), .B(_421_), .C(_422_), .Y(_0__26_) );
INVX1 INVX1_70 ( .A(_33__3_), .Y(_423_) );
NAND2X1 NAND2X1_110 ( .A(w_cout_5_), .B(_34__3_), .Y(_424_) );
OAI21X1 OAI21X1_110 ( .A(w_cout_5_), .B(_423_), .C(_424_), .Y(_0__27_) );
INVX1 INVX1_71 ( .A(1'b0), .Y(_428_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_429_) );
NAND2X1 NAND2X1_111 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_430_) );
NAND3X1 NAND3X1_41 ( .A(_428_), .B(_430_), .C(_429_), .Y(_431_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_425_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_426_) );
OAI21X1 OAI21X1_111 ( .A(_425_), .B(_426_), .C(1'b0), .Y(_427_) );
NAND2X1 NAND2X1_112 ( .A(_427_), .B(_431_), .Y(_33__0_) );
OAI21X1 OAI21X1_112 ( .A(_428_), .B(_425_), .C(_430_), .Y(_35__1_) );
INVX1 INVX1_72 ( .A(_35__3_), .Y(_435_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_436_) );
NAND2X1 NAND2X1_113 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_437_) );
NAND3X1 NAND3X1_42 ( .A(_435_), .B(_437_), .C(_436_), .Y(_438_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_432_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_433_) );
OAI21X1 OAI21X1_113 ( .A(_432_), .B(_433_), .C(_35__3_), .Y(_434_) );
NAND2X1 NAND2X1_114 ( .A(_434_), .B(_438_), .Y(_33__3_) );
OAI21X1 OAI21X1_114 ( .A(_435_), .B(_432_), .C(_437_), .Y(_31_) );
INVX1 INVX1_73 ( .A(_35__1_), .Y(_442_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_443_) );
NAND2X1 NAND2X1_115 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_444_) );
NAND3X1 NAND3X1_43 ( .A(_442_), .B(_444_), .C(_443_), .Y(_445_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_439_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_440_) );
OAI21X1 OAI21X1_115 ( .A(_439_), .B(_440_), .C(_35__1_), .Y(_441_) );
NAND2X1 NAND2X1_116 ( .A(_441_), .B(_445_), .Y(_33__1_) );
OAI21X1 OAI21X1_116 ( .A(_442_), .B(_439_), .C(_444_), .Y(_35__2_) );
INVX1 INVX1_74 ( .A(_35__2_), .Y(_449_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_450_) );
NAND2X1 NAND2X1_117 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_451_) );
NAND3X1 NAND3X1_44 ( .A(_449_), .B(_451_), .C(_450_), .Y(_452_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_446_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_447_) );
OAI21X1 OAI21X1_117 ( .A(_446_), .B(_447_), .C(_35__2_), .Y(_448_) );
NAND2X1 NAND2X1_118 ( .A(_448_), .B(_452_), .Y(_33__2_) );
OAI21X1 OAI21X1_118 ( .A(_449_), .B(_446_), .C(_451_), .Y(_35__3_) );
INVX1 INVX1_75 ( .A(1'b1), .Y(_456_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_457_) );
NAND2X1 NAND2X1_119 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_458_) );
NAND3X1 NAND3X1_45 ( .A(_456_), .B(_458_), .C(_457_), .Y(_459_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_453_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_454_) );
OAI21X1 OAI21X1_119 ( .A(_453_), .B(_454_), .C(1'b1), .Y(_455_) );
NAND2X1 NAND2X1_120 ( .A(_455_), .B(_459_), .Y(_34__0_) );
OAI21X1 OAI21X1_120 ( .A(_456_), .B(_453_), .C(_458_), .Y(_36__1_) );
INVX1 INVX1_76 ( .A(_36__3_), .Y(_463_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_464_) );
NAND2X1 NAND2X1_121 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_465_) );
NAND3X1 NAND3X1_46 ( .A(_463_), .B(_465_), .C(_464_), .Y(_466_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_460_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_461_) );
OAI21X1 OAI21X1_121 ( .A(_460_), .B(_461_), .C(_36__3_), .Y(_462_) );
NAND2X1 NAND2X1_122 ( .A(_462_), .B(_466_), .Y(_34__3_) );
OAI21X1 OAI21X1_122 ( .A(_463_), .B(_460_), .C(_465_), .Y(_32_) );
INVX1 INVX1_77 ( .A(_36__1_), .Y(_470_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_471_) );
NAND2X1 NAND2X1_123 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_472_) );
NAND3X1 NAND3X1_47 ( .A(_470_), .B(_472_), .C(_471_), .Y(_473_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_467_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_468_) );
OAI21X1 OAI21X1_123 ( .A(_467_), .B(_468_), .C(_36__1_), .Y(_469_) );
NAND2X1 NAND2X1_124 ( .A(_469_), .B(_473_), .Y(_34__1_) );
OAI21X1 OAI21X1_124 ( .A(_470_), .B(_467_), .C(_472_), .Y(_36__2_) );
INVX1 INVX1_78 ( .A(_36__2_), .Y(_477_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_478_) );
NAND2X1 NAND2X1_125 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_479_) );
NAND3X1 NAND3X1_48 ( .A(_477_), .B(_479_), .C(_478_), .Y(_480_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_474_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_475_) );
OAI21X1 OAI21X1_125 ( .A(_474_), .B(_475_), .C(_36__2_), .Y(_476_) );
NAND2X1 NAND2X1_126 ( .A(_476_), .B(_480_), .Y(_34__2_) );
OAI21X1 OAI21X1_126 ( .A(_477_), .B(_474_), .C(_479_), .Y(_36__3_) );
INVX1 INVX1_79 ( .A(_37_), .Y(_481_) );
NAND2X1 NAND2X1_127 ( .A(_38_), .B(w_cout_6_), .Y(_482_) );
OAI21X1 OAI21X1_127 ( .A(w_cout_6_), .B(_481_), .C(_482_), .Y(w_cout_7_) );
INVX1 INVX1_80 ( .A(_39__0_), .Y(_483_) );
NAND2X1 NAND2X1_128 ( .A(_40__0_), .B(w_cout_6_), .Y(_484_) );
OAI21X1 OAI21X1_128 ( .A(w_cout_6_), .B(_483_), .C(_484_), .Y(_0__28_) );
INVX1 INVX1_81 ( .A(_39__1_), .Y(_485_) );
NAND2X1 NAND2X1_129 ( .A(w_cout_6_), .B(_40__1_), .Y(_486_) );
OAI21X1 OAI21X1_129 ( .A(w_cout_6_), .B(_485_), .C(_486_), .Y(_0__29_) );
INVX1 INVX1_82 ( .A(_39__2_), .Y(_487_) );
NAND2X1 NAND2X1_130 ( .A(w_cout_6_), .B(_40__2_), .Y(_488_) );
OAI21X1 OAI21X1_130 ( .A(w_cout_6_), .B(_487_), .C(_488_), .Y(_0__30_) );
INVX1 INVX1_83 ( .A(_39__3_), .Y(_489_) );
NAND2X1 NAND2X1_131 ( .A(w_cout_6_), .B(_40__3_), .Y(_490_) );
OAI21X1 OAI21X1_131 ( .A(w_cout_6_), .B(_489_), .C(_490_), .Y(_0__31_) );
INVX1 INVX1_84 ( .A(1'b0), .Y(_494_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_495_) );
NAND2X1 NAND2X1_132 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_496_) );
NAND3X1 NAND3X1_49 ( .A(_494_), .B(_496_), .C(_495_), .Y(_497_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_491_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_492_) );
OAI21X1 OAI21X1_132 ( .A(_491_), .B(_492_), .C(1'b0), .Y(_493_) );
NAND2X1 NAND2X1_133 ( .A(_493_), .B(_497_), .Y(_39__0_) );
OAI21X1 OAI21X1_133 ( .A(_494_), .B(_491_), .C(_496_), .Y(_41__1_) );
INVX1 INVX1_85 ( .A(_41__3_), .Y(_501_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_502_) );
NAND2X1 NAND2X1_134 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_503_) );
NAND3X1 NAND3X1_50 ( .A(_501_), .B(_503_), .C(_502_), .Y(_504_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_498_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_499_) );
OAI21X1 OAI21X1_134 ( .A(_498_), .B(_499_), .C(_41__3_), .Y(_500_) );
NAND2X1 NAND2X1_135 ( .A(_500_), .B(_504_), .Y(_39__3_) );
OAI21X1 OAI21X1_135 ( .A(_501_), .B(_498_), .C(_503_), .Y(_37_) );
INVX1 INVX1_86 ( .A(_41__1_), .Y(_508_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_509_) );
NAND2X1 NAND2X1_136 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_510_) );
NAND3X1 NAND3X1_51 ( .A(_508_), .B(_510_), .C(_509_), .Y(_511_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_505_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_506_) );
OAI21X1 OAI21X1_136 ( .A(_505_), .B(_506_), .C(_41__1_), .Y(_507_) );
NAND2X1 NAND2X1_137 ( .A(_507_), .B(_511_), .Y(_39__1_) );
OAI21X1 OAI21X1_137 ( .A(_508_), .B(_505_), .C(_510_), .Y(_41__2_) );
INVX1 INVX1_87 ( .A(_41__2_), .Y(_515_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_516_) );
NAND2X1 NAND2X1_138 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_517_) );
NAND3X1 NAND3X1_52 ( .A(_515_), .B(_517_), .C(_516_), .Y(_518_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_512_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_513_) );
OAI21X1 OAI21X1_138 ( .A(_512_), .B(_513_), .C(_41__2_), .Y(_514_) );
NAND2X1 NAND2X1_139 ( .A(_514_), .B(_518_), .Y(_39__2_) );
OAI21X1 OAI21X1_139 ( .A(_515_), .B(_512_), .C(_517_), .Y(_41__3_) );
INVX1 INVX1_88 ( .A(1'b1), .Y(_522_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_523_) );
NAND2X1 NAND2X1_140 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_524_) );
NAND3X1 NAND3X1_53 ( .A(_522_), .B(_524_), .C(_523_), .Y(_525_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_519_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_520_) );
OAI21X1 OAI21X1_140 ( .A(_519_), .B(_520_), .C(1'b1), .Y(_521_) );
NAND2X1 NAND2X1_141 ( .A(_521_), .B(_525_), .Y(_40__0_) );
OAI21X1 OAI21X1_141 ( .A(_522_), .B(_519_), .C(_524_), .Y(_42__1_) );
INVX1 INVX1_89 ( .A(_42__3_), .Y(_529_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_530_) );
NAND2X1 NAND2X1_142 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_531_) );
NAND3X1 NAND3X1_54 ( .A(_529_), .B(_531_), .C(_530_), .Y(_532_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_526_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_527_) );
OAI21X1 OAI21X1_142 ( .A(_526_), .B(_527_), .C(_42__3_), .Y(_528_) );
NAND2X1 NAND2X1_143 ( .A(_528_), .B(_532_), .Y(_40__3_) );
OAI21X1 OAI21X1_143 ( .A(_529_), .B(_526_), .C(_531_), .Y(_38_) );
INVX1 INVX1_90 ( .A(_42__1_), .Y(_536_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_537_) );
NAND2X1 NAND2X1_144 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_538_) );
NAND3X1 NAND3X1_55 ( .A(_536_), .B(_538_), .C(_537_), .Y(_539_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_533_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_534_) );
OAI21X1 OAI21X1_144 ( .A(_533_), .B(_534_), .C(_42__1_), .Y(_535_) );
NAND2X1 NAND2X1_145 ( .A(_535_), .B(_539_), .Y(_40__1_) );
OAI21X1 OAI21X1_145 ( .A(_536_), .B(_533_), .C(_538_), .Y(_42__2_) );
INVX1 INVX1_91 ( .A(_42__2_), .Y(_543_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_544_) );
NAND2X1 NAND2X1_146 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_545_) );
NAND3X1 NAND3X1_56 ( .A(_543_), .B(_545_), .C(_544_), .Y(_546_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_540_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_541_) );
OAI21X1 OAI21X1_146 ( .A(_540_), .B(_541_), .C(_42__2_), .Y(_542_) );
NAND2X1 NAND2X1_147 ( .A(_542_), .B(_546_), .Y(_40__2_) );
OAI21X1 OAI21X1_147 ( .A(_543_), .B(_540_), .C(_545_), .Y(_42__3_) );
INVX1 INVX1_92 ( .A(_43_), .Y(_547_) );
NAND2X1 NAND2X1_148 ( .A(_44_), .B(w_cout_7_), .Y(_548_) );
OAI21X1 OAI21X1_148 ( .A(w_cout_7_), .B(_547_), .C(_548_), .Y(w_cout_8_) );
INVX1 INVX1_93 ( .A(_45__0_), .Y(_549_) );
NAND2X1 NAND2X1_149 ( .A(_46__0_), .B(w_cout_7_), .Y(_550_) );
OAI21X1 OAI21X1_149 ( .A(w_cout_7_), .B(_549_), .C(_550_), .Y(_0__32_) );
INVX1 INVX1_94 ( .A(_45__1_), .Y(_551_) );
NAND2X1 NAND2X1_150 ( .A(w_cout_7_), .B(_46__1_), .Y(_552_) );
OAI21X1 OAI21X1_150 ( .A(w_cout_7_), .B(_551_), .C(_552_), .Y(_0__33_) );
INVX1 INVX1_95 ( .A(_45__2_), .Y(_553_) );
NAND2X1 NAND2X1_151 ( .A(w_cout_7_), .B(_46__2_), .Y(_554_) );
OAI21X1 OAI21X1_151 ( .A(w_cout_7_), .B(_553_), .C(_554_), .Y(_0__34_) );
INVX1 INVX1_96 ( .A(_45__3_), .Y(_555_) );
NAND2X1 NAND2X1_152 ( .A(w_cout_7_), .B(_46__3_), .Y(_556_) );
OAI21X1 OAI21X1_152 ( .A(w_cout_7_), .B(_555_), .C(_556_), .Y(_0__35_) );
INVX1 INVX1_97 ( .A(1'b0), .Y(_560_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_561_) );
NAND2X1 NAND2X1_153 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_562_) );
NAND3X1 NAND3X1_57 ( .A(_560_), .B(_562_), .C(_561_), .Y(_563_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_557_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_558_) );
OAI21X1 OAI21X1_153 ( .A(_557_), .B(_558_), .C(1'b0), .Y(_559_) );
NAND2X1 NAND2X1_154 ( .A(_559_), .B(_563_), .Y(_45__0_) );
OAI21X1 OAI21X1_154 ( .A(_560_), .B(_557_), .C(_562_), .Y(_47__1_) );
INVX1 INVX1_98 ( .A(_47__3_), .Y(_567_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_568_) );
NAND2X1 NAND2X1_155 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_569_) );
NAND3X1 NAND3X1_58 ( .A(_567_), .B(_569_), .C(_568_), .Y(_570_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_564_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_565_) );
OAI21X1 OAI21X1_155 ( .A(_564_), .B(_565_), .C(_47__3_), .Y(_566_) );
NAND2X1 NAND2X1_156 ( .A(_566_), .B(_570_), .Y(_45__3_) );
OAI21X1 OAI21X1_156 ( .A(_567_), .B(_564_), .C(_569_), .Y(_43_) );
INVX1 INVX1_99 ( .A(_47__1_), .Y(_574_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_575_) );
NAND2X1 NAND2X1_157 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_576_) );
NAND3X1 NAND3X1_59 ( .A(_574_), .B(_576_), .C(_575_), .Y(_577_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_571_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_572_) );
OAI21X1 OAI21X1_157 ( .A(_571_), .B(_572_), .C(_47__1_), .Y(_573_) );
NAND2X1 NAND2X1_158 ( .A(_573_), .B(_577_), .Y(_45__1_) );
OAI21X1 OAI21X1_158 ( .A(_574_), .B(_571_), .C(_576_), .Y(_47__2_) );
INVX1 INVX1_100 ( .A(_47__2_), .Y(_581_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_582_) );
NAND2X1 NAND2X1_159 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_583_) );
NAND3X1 NAND3X1_60 ( .A(_581_), .B(_583_), .C(_582_), .Y(_584_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_578_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_579_) );
OAI21X1 OAI21X1_159 ( .A(_578_), .B(_579_), .C(_47__2_), .Y(_580_) );
NAND2X1 NAND2X1_160 ( .A(_580_), .B(_584_), .Y(_45__2_) );
OAI21X1 OAI21X1_160 ( .A(_581_), .B(_578_), .C(_583_), .Y(_47__3_) );
INVX1 INVX1_101 ( .A(1'b1), .Y(_588_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_589_) );
NAND2X1 NAND2X1_161 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_590_) );
NAND3X1 NAND3X1_61 ( .A(_588_), .B(_590_), .C(_589_), .Y(_591_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_585_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_586_) );
OAI21X1 OAI21X1_161 ( .A(_585_), .B(_586_), .C(1'b1), .Y(_587_) );
NAND2X1 NAND2X1_162 ( .A(_587_), .B(_591_), .Y(_46__0_) );
OAI21X1 OAI21X1_162 ( .A(_588_), .B(_585_), .C(_590_), .Y(_48__1_) );
INVX1 INVX1_102 ( .A(_48__3_), .Y(_595_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_596_) );
NAND2X1 NAND2X1_163 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_597_) );
NAND3X1 NAND3X1_62 ( .A(_595_), .B(_597_), .C(_596_), .Y(_598_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_592_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_593_) );
OAI21X1 OAI21X1_163 ( .A(_592_), .B(_593_), .C(_48__3_), .Y(_594_) );
NAND2X1 NAND2X1_164 ( .A(_594_), .B(_598_), .Y(_46__3_) );
OAI21X1 OAI21X1_164 ( .A(_595_), .B(_592_), .C(_597_), .Y(_44_) );
INVX1 INVX1_103 ( .A(_48__1_), .Y(_602_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_603_) );
NAND2X1 NAND2X1_165 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_604_) );
NAND3X1 NAND3X1_63 ( .A(_602_), .B(_604_), .C(_603_), .Y(_605_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_599_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_600_) );
OAI21X1 OAI21X1_165 ( .A(_599_), .B(_600_), .C(_48__1_), .Y(_601_) );
NAND2X1 NAND2X1_166 ( .A(_601_), .B(_605_), .Y(_46__1_) );
OAI21X1 OAI21X1_166 ( .A(_602_), .B(_599_), .C(_604_), .Y(_48__2_) );
INVX1 INVX1_104 ( .A(_48__2_), .Y(_609_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_610_) );
NAND2X1 NAND2X1_167 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_611_) );
NAND3X1 NAND3X1_64 ( .A(_609_), .B(_611_), .C(_610_), .Y(_612_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_606_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_607_) );
OAI21X1 OAI21X1_167 ( .A(_606_), .B(_607_), .C(_48__2_), .Y(_608_) );
NAND2X1 NAND2X1_168 ( .A(_608_), .B(_612_), .Y(_46__2_) );
OAI21X1 OAI21X1_168 ( .A(_609_), .B(_606_), .C(_611_), .Y(_48__3_) );
INVX1 INVX1_105 ( .A(_49_), .Y(_613_) );
NAND2X1 NAND2X1_169 ( .A(_50_), .B(w_cout_8_), .Y(_614_) );
OAI21X1 OAI21X1_169 ( .A(w_cout_8_), .B(_613_), .C(_614_), .Y(w_cout_9_) );
INVX1 INVX1_106 ( .A(_51__0_), .Y(_615_) );
NAND2X1 NAND2X1_170 ( .A(_52__0_), .B(w_cout_8_), .Y(_616_) );
OAI21X1 OAI21X1_170 ( .A(w_cout_8_), .B(_615_), .C(_616_), .Y(_0__36_) );
INVX1 INVX1_107 ( .A(_51__1_), .Y(_617_) );
NAND2X1 NAND2X1_171 ( .A(w_cout_8_), .B(_52__1_), .Y(_618_) );
OAI21X1 OAI21X1_171 ( .A(w_cout_8_), .B(_617_), .C(_618_), .Y(_0__37_) );
INVX1 INVX1_108 ( .A(_51__2_), .Y(_619_) );
NAND2X1 NAND2X1_172 ( .A(w_cout_8_), .B(_52__2_), .Y(_620_) );
OAI21X1 OAI21X1_172 ( .A(w_cout_8_), .B(_619_), .C(_620_), .Y(_0__38_) );
INVX1 INVX1_109 ( .A(_51__3_), .Y(_621_) );
NAND2X1 NAND2X1_173 ( .A(w_cout_8_), .B(_52__3_), .Y(_622_) );
OAI21X1 OAI21X1_173 ( .A(w_cout_8_), .B(_621_), .C(_622_), .Y(_0__39_) );
INVX1 INVX1_110 ( .A(1'b0), .Y(_626_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_627_) );
NAND2X1 NAND2X1_174 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_628_) );
NAND3X1 NAND3X1_65 ( .A(_626_), .B(_628_), .C(_627_), .Y(_629_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_623_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_624_) );
OAI21X1 OAI21X1_174 ( .A(_623_), .B(_624_), .C(1'b0), .Y(_625_) );
NAND2X1 NAND2X1_175 ( .A(_625_), .B(_629_), .Y(_51__0_) );
OAI21X1 OAI21X1_175 ( .A(_626_), .B(_623_), .C(_628_), .Y(_53__1_) );
INVX1 INVX1_111 ( .A(_53__3_), .Y(_633_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_634_) );
NAND2X1 NAND2X1_176 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_635_) );
NAND3X1 NAND3X1_66 ( .A(_633_), .B(_635_), .C(_634_), .Y(_636_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_630_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_631_) );
OAI21X1 OAI21X1_176 ( .A(_630_), .B(_631_), .C(_53__3_), .Y(_632_) );
NAND2X1 NAND2X1_177 ( .A(_632_), .B(_636_), .Y(_51__3_) );
OAI21X1 OAI21X1_177 ( .A(_633_), .B(_630_), .C(_635_), .Y(_49_) );
INVX1 INVX1_112 ( .A(_53__1_), .Y(_640_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_641_) );
NAND2X1 NAND2X1_178 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_642_) );
NAND3X1 NAND3X1_67 ( .A(_640_), .B(_642_), .C(_641_), .Y(_643_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_637_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_638_) );
OAI21X1 OAI21X1_178 ( .A(_637_), .B(_638_), .C(_53__1_), .Y(_639_) );
NAND2X1 NAND2X1_179 ( .A(_639_), .B(_643_), .Y(_51__1_) );
OAI21X1 OAI21X1_179 ( .A(_640_), .B(_637_), .C(_642_), .Y(_53__2_) );
INVX1 INVX1_113 ( .A(_53__2_), .Y(_647_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_648_) );
NAND2X1 NAND2X1_180 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_649_) );
NAND3X1 NAND3X1_68 ( .A(_647_), .B(_649_), .C(_648_), .Y(_650_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_644_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_645_) );
OAI21X1 OAI21X1_180 ( .A(_644_), .B(_645_), .C(_53__2_), .Y(_646_) );
NAND2X1 NAND2X1_181 ( .A(_646_), .B(_650_), .Y(_51__2_) );
OAI21X1 OAI21X1_181 ( .A(_647_), .B(_644_), .C(_649_), .Y(_53__3_) );
INVX1 INVX1_114 ( .A(1'b1), .Y(_654_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_655_) );
NAND2X1 NAND2X1_182 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_656_) );
NAND3X1 NAND3X1_69 ( .A(_654_), .B(_656_), .C(_655_), .Y(_657_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_651_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_652_) );
OAI21X1 OAI21X1_182 ( .A(_651_), .B(_652_), .C(1'b1), .Y(_653_) );
NAND2X1 NAND2X1_183 ( .A(_653_), .B(_657_), .Y(_52__0_) );
OAI21X1 OAI21X1_183 ( .A(_654_), .B(_651_), .C(_656_), .Y(_54__1_) );
INVX1 INVX1_115 ( .A(_54__3_), .Y(_661_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_662_) );
NAND2X1 NAND2X1_184 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_663_) );
NAND3X1 NAND3X1_70 ( .A(_661_), .B(_663_), .C(_662_), .Y(_664_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_658_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_659_) );
OAI21X1 OAI21X1_184 ( .A(_658_), .B(_659_), .C(_54__3_), .Y(_660_) );
NAND2X1 NAND2X1_185 ( .A(_660_), .B(_664_), .Y(_52__3_) );
OAI21X1 OAI21X1_185 ( .A(_661_), .B(_658_), .C(_663_), .Y(_50_) );
INVX1 INVX1_116 ( .A(_54__1_), .Y(_668_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_669_) );
NAND2X1 NAND2X1_186 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_670_) );
NAND3X1 NAND3X1_71 ( .A(_668_), .B(_670_), .C(_669_), .Y(_671_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_665_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_666_) );
OAI21X1 OAI21X1_186 ( .A(_665_), .B(_666_), .C(_54__1_), .Y(_667_) );
NAND2X1 NAND2X1_187 ( .A(_667_), .B(_671_), .Y(_52__1_) );
OAI21X1 OAI21X1_187 ( .A(_668_), .B(_665_), .C(_670_), .Y(_54__2_) );
INVX1 INVX1_117 ( .A(_54__2_), .Y(_675_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_676_) );
NAND2X1 NAND2X1_188 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_677_) );
NAND3X1 NAND3X1_72 ( .A(_675_), .B(_677_), .C(_676_), .Y(_678_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_672_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_673_) );
OAI21X1 OAI21X1_188 ( .A(_672_), .B(_673_), .C(_54__2_), .Y(_674_) );
NAND2X1 NAND2X1_189 ( .A(_674_), .B(_678_), .Y(_52__2_) );
OAI21X1 OAI21X1_189 ( .A(_675_), .B(_672_), .C(_677_), .Y(_54__3_) );
INVX1 INVX1_118 ( .A(_55_), .Y(_679_) );
NAND2X1 NAND2X1_190 ( .A(_56_), .B(w_cout_9_), .Y(_680_) );
OAI21X1 OAI21X1_190 ( .A(w_cout_9_), .B(_679_), .C(_680_), .Y(w_cout_10_) );
INVX1 INVX1_119 ( .A(_57__0_), .Y(_681_) );
NAND2X1 NAND2X1_191 ( .A(_58__0_), .B(w_cout_9_), .Y(_682_) );
OAI21X1 OAI21X1_191 ( .A(w_cout_9_), .B(_681_), .C(_682_), .Y(_0__40_) );
INVX1 INVX1_120 ( .A(_57__1_), .Y(_683_) );
NAND2X1 NAND2X1_192 ( .A(w_cout_9_), .B(_58__1_), .Y(_684_) );
OAI21X1 OAI21X1_192 ( .A(w_cout_9_), .B(_683_), .C(_684_), .Y(_0__41_) );
INVX1 INVX1_121 ( .A(_57__2_), .Y(_685_) );
NAND2X1 NAND2X1_193 ( .A(w_cout_9_), .B(_58__2_), .Y(_686_) );
OAI21X1 OAI21X1_193 ( .A(w_cout_9_), .B(_685_), .C(_686_), .Y(_0__42_) );
INVX1 INVX1_122 ( .A(_57__3_), .Y(_687_) );
NAND2X1 NAND2X1_194 ( .A(w_cout_9_), .B(_58__3_), .Y(_688_) );
OAI21X1 OAI21X1_194 ( .A(w_cout_9_), .B(_687_), .C(_688_), .Y(_0__43_) );
INVX1 INVX1_123 ( .A(1'b0), .Y(_692_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_693_) );
NAND2X1 NAND2X1_195 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_694_) );
NAND3X1 NAND3X1_73 ( .A(_692_), .B(_694_), .C(_693_), .Y(_695_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_689_) );
AND2X2 AND2X2_73 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_690_) );
OAI21X1 OAI21X1_195 ( .A(_689_), .B(_690_), .C(1'b0), .Y(_691_) );
NAND2X1 NAND2X1_196 ( .A(_691_), .B(_695_), .Y(_57__0_) );
OAI21X1 OAI21X1_196 ( .A(_692_), .B(_689_), .C(_694_), .Y(_59__1_) );
INVX1 INVX1_124 ( .A(_59__3_), .Y(_699_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_700_) );
NAND2X1 NAND2X1_197 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_701_) );
NAND3X1 NAND3X1_74 ( .A(_699_), .B(_701_), .C(_700_), .Y(_702_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_696_) );
AND2X2 AND2X2_74 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_697_) );
OAI21X1 OAI21X1_197 ( .A(_696_), .B(_697_), .C(_59__3_), .Y(_698_) );
NAND2X1 NAND2X1_198 ( .A(_698_), .B(_702_), .Y(_57__3_) );
OAI21X1 OAI21X1_198 ( .A(_699_), .B(_696_), .C(_701_), .Y(_55_) );
INVX1 INVX1_125 ( .A(_59__1_), .Y(_706_) );
OR2X2 OR2X2_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_707_) );
NAND2X1 NAND2X1_199 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_708_) );
NAND3X1 NAND3X1_75 ( .A(_706_), .B(_708_), .C(_707_), .Y(_709_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_703_) );
AND2X2 AND2X2_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_704_) );
OAI21X1 OAI21X1_199 ( .A(_703_), .B(_704_), .C(_59__1_), .Y(_705_) );
NAND2X1 NAND2X1_200 ( .A(_705_), .B(_709_), .Y(_57__1_) );
OAI21X1 OAI21X1_200 ( .A(_706_), .B(_703_), .C(_708_), .Y(_59__2_) );
INVX1 INVX1_126 ( .A(_59__2_), .Y(_713_) );
OR2X2 OR2X2_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_714_) );
NAND2X1 NAND2X1_201 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_715_) );
NAND3X1 NAND3X1_76 ( .A(_713_), .B(_715_), .C(_714_), .Y(_716_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_710_) );
AND2X2 AND2X2_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_711_) );
OAI21X1 OAI21X1_201 ( .A(_710_), .B(_711_), .C(_59__2_), .Y(_712_) );
NAND2X1 NAND2X1_202 ( .A(_712_), .B(_716_), .Y(_57__2_) );
OAI21X1 OAI21X1_202 ( .A(_713_), .B(_710_), .C(_715_), .Y(_59__3_) );
INVX1 INVX1_127 ( .A(1'b1), .Y(_720_) );
OR2X2 OR2X2_77 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_721_) );
NAND2X1 NAND2X1_203 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_722_) );
NAND3X1 NAND3X1_77 ( .A(_720_), .B(_722_), .C(_721_), .Y(_723_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_717_) );
AND2X2 AND2X2_77 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_718_) );
OAI21X1 OAI21X1_203 ( .A(_717_), .B(_718_), .C(1'b1), .Y(_719_) );
NAND2X1 NAND2X1_204 ( .A(_719_), .B(_723_), .Y(_58__0_) );
OAI21X1 OAI21X1_204 ( .A(_720_), .B(_717_), .C(_722_), .Y(_60__1_) );
INVX1 INVX1_128 ( .A(_60__3_), .Y(_727_) );
OR2X2 OR2X2_78 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_728_) );
NAND2X1 NAND2X1_205 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_729_) );
NAND3X1 NAND3X1_78 ( .A(_727_), .B(_729_), .C(_728_), .Y(_730_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_724_) );
AND2X2 AND2X2_78 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_725_) );
OAI21X1 OAI21X1_205 ( .A(_724_), .B(_725_), .C(_60__3_), .Y(_726_) );
NAND2X1 NAND2X1_206 ( .A(_726_), .B(_730_), .Y(_58__3_) );
OAI21X1 OAI21X1_206 ( .A(_727_), .B(_724_), .C(_729_), .Y(_56_) );
INVX1 INVX1_129 ( .A(_60__1_), .Y(_734_) );
OR2X2 OR2X2_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_735_) );
NAND2X1 NAND2X1_207 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_736_) );
NAND3X1 NAND3X1_79 ( .A(_734_), .B(_736_), .C(_735_), .Y(_737_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_731_) );
AND2X2 AND2X2_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_732_) );
OAI21X1 OAI21X1_207 ( .A(_731_), .B(_732_), .C(_60__1_), .Y(_733_) );
NAND2X1 NAND2X1_208 ( .A(_733_), .B(_737_), .Y(_58__1_) );
OAI21X1 OAI21X1_208 ( .A(_734_), .B(_731_), .C(_736_), .Y(_60__2_) );
INVX1 INVX1_130 ( .A(_60__2_), .Y(_741_) );
OR2X2 OR2X2_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_742_) );
NAND2X1 NAND2X1_209 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_743_) );
NAND3X1 NAND3X1_80 ( .A(_741_), .B(_743_), .C(_742_), .Y(_744_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_738_) );
AND2X2 AND2X2_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_739_) );
OAI21X1 OAI21X1_209 ( .A(_738_), .B(_739_), .C(_60__2_), .Y(_740_) );
NAND2X1 NAND2X1_210 ( .A(_740_), .B(_744_), .Y(_58__2_) );
OAI21X1 OAI21X1_210 ( .A(_741_), .B(_738_), .C(_743_), .Y(_60__3_) );
INVX1 INVX1_131 ( .A(_61_), .Y(_745_) );
NAND2X1 NAND2X1_211 ( .A(_62_), .B(w_cout_10_), .Y(_746_) );
OAI21X1 OAI21X1_211 ( .A(w_cout_10_), .B(_745_), .C(_746_), .Y(w_cout_11_) );
INVX1 INVX1_132 ( .A(_63__0_), .Y(_747_) );
NAND2X1 NAND2X1_212 ( .A(_64__0_), .B(w_cout_10_), .Y(_748_) );
OAI21X1 OAI21X1_212 ( .A(w_cout_10_), .B(_747_), .C(_748_), .Y(_0__44_) );
INVX1 INVX1_133 ( .A(_63__1_), .Y(_749_) );
NAND2X1 NAND2X1_213 ( .A(w_cout_10_), .B(_64__1_), .Y(_750_) );
OAI21X1 OAI21X1_213 ( .A(w_cout_10_), .B(_749_), .C(_750_), .Y(_0__45_) );
INVX1 INVX1_134 ( .A(_63__2_), .Y(_751_) );
NAND2X1 NAND2X1_214 ( .A(w_cout_10_), .B(_64__2_), .Y(_752_) );
OAI21X1 OAI21X1_214 ( .A(w_cout_10_), .B(_751_), .C(_752_), .Y(_0__46_) );
INVX1 INVX1_135 ( .A(_63__3_), .Y(_753_) );
NAND2X1 NAND2X1_215 ( .A(w_cout_10_), .B(_64__3_), .Y(_754_) );
OAI21X1 OAI21X1_215 ( .A(w_cout_10_), .B(_753_), .C(_754_), .Y(_0__47_) );
INVX1 INVX1_136 ( .A(1'b0), .Y(_758_) );
OR2X2 OR2X2_81 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_759_) );
NAND2X1 NAND2X1_216 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_760_) );
NAND3X1 NAND3X1_81 ( .A(_758_), .B(_760_), .C(_759_), .Y(_761_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_755_) );
AND2X2 AND2X2_81 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_756_) );
OAI21X1 OAI21X1_216 ( .A(_755_), .B(_756_), .C(1'b0), .Y(_757_) );
NAND2X1 NAND2X1_217 ( .A(_757_), .B(_761_), .Y(_63__0_) );
OAI21X1 OAI21X1_217 ( .A(_758_), .B(_755_), .C(_760_), .Y(_65__1_) );
INVX1 INVX1_137 ( .A(_65__3_), .Y(_765_) );
OR2X2 OR2X2_82 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_766_) );
NAND2X1 NAND2X1_218 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_767_) );
NAND3X1 NAND3X1_82 ( .A(_765_), .B(_767_), .C(_766_), .Y(_768_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_762_) );
AND2X2 AND2X2_82 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_763_) );
OAI21X1 OAI21X1_218 ( .A(_762_), .B(_763_), .C(_65__3_), .Y(_764_) );
NAND2X1 NAND2X1_219 ( .A(_764_), .B(_768_), .Y(_63__3_) );
OAI21X1 OAI21X1_219 ( .A(_765_), .B(_762_), .C(_767_), .Y(_61_) );
INVX1 INVX1_138 ( .A(_65__1_), .Y(_772_) );
OR2X2 OR2X2_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_773_) );
NAND2X1 NAND2X1_220 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_774_) );
NAND3X1 NAND3X1_83 ( .A(_772_), .B(_774_), .C(_773_), .Y(_775_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_769_) );
AND2X2 AND2X2_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_770_) );
OAI21X1 OAI21X1_220 ( .A(_769_), .B(_770_), .C(_65__1_), .Y(_771_) );
NAND2X1 NAND2X1_221 ( .A(_771_), .B(_775_), .Y(_63__1_) );
OAI21X1 OAI21X1_221 ( .A(_772_), .B(_769_), .C(_774_), .Y(_65__2_) );
INVX1 INVX1_139 ( .A(_65__2_), .Y(_779_) );
OR2X2 OR2X2_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_780_) );
NAND2X1 NAND2X1_222 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_781_) );
NAND3X1 NAND3X1_84 ( .A(_779_), .B(_781_), .C(_780_), .Y(_782_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_776_) );
AND2X2 AND2X2_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_777_) );
OAI21X1 OAI21X1_222 ( .A(_776_), .B(_777_), .C(_65__2_), .Y(_778_) );
NAND2X1 NAND2X1_223 ( .A(_778_), .B(_782_), .Y(_63__2_) );
OAI21X1 OAI21X1_223 ( .A(_779_), .B(_776_), .C(_781_), .Y(_65__3_) );
INVX1 INVX1_140 ( .A(1'b1), .Y(_786_) );
OR2X2 OR2X2_85 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_787_) );
NAND2X1 NAND2X1_224 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_788_) );
NAND3X1 NAND3X1_85 ( .A(_786_), .B(_788_), .C(_787_), .Y(_789_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_783_) );
AND2X2 AND2X2_85 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_784_) );
OAI21X1 OAI21X1_224 ( .A(_783_), .B(_784_), .C(1'b1), .Y(_785_) );
NAND2X1 NAND2X1_225 ( .A(_785_), .B(_789_), .Y(_64__0_) );
OAI21X1 OAI21X1_225 ( .A(_786_), .B(_783_), .C(_788_), .Y(_66__1_) );
INVX1 INVX1_141 ( .A(_66__3_), .Y(_793_) );
OR2X2 OR2X2_86 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_794_) );
NAND2X1 NAND2X1_226 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_795_) );
NAND3X1 NAND3X1_86 ( .A(_793_), .B(_795_), .C(_794_), .Y(_796_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_790_) );
AND2X2 AND2X2_86 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_791_) );
OAI21X1 OAI21X1_226 ( .A(_790_), .B(_791_), .C(_66__3_), .Y(_792_) );
NAND2X1 NAND2X1_227 ( .A(_792_), .B(_796_), .Y(_64__3_) );
OAI21X1 OAI21X1_227 ( .A(_793_), .B(_790_), .C(_795_), .Y(_62_) );
INVX1 INVX1_142 ( .A(_66__1_), .Y(_800_) );
OR2X2 OR2X2_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_801_) );
NAND2X1 NAND2X1_228 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_802_) );
NAND3X1 NAND3X1_87 ( .A(_800_), .B(_802_), .C(_801_), .Y(_803_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_797_) );
AND2X2 AND2X2_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_798_) );
OAI21X1 OAI21X1_228 ( .A(_797_), .B(_798_), .C(_66__1_), .Y(_799_) );
NAND2X1 NAND2X1_229 ( .A(_799_), .B(_803_), .Y(_64__1_) );
OAI21X1 OAI21X1_229 ( .A(_800_), .B(_797_), .C(_802_), .Y(_66__2_) );
INVX1 INVX1_143 ( .A(_66__2_), .Y(_807_) );
OR2X2 OR2X2_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_808_) );
NAND2X1 NAND2X1_230 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_809_) );
NAND3X1 NAND3X1_88 ( .A(_807_), .B(_809_), .C(_808_), .Y(_810_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_804_) );
AND2X2 AND2X2_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_805_) );
OAI21X1 OAI21X1_230 ( .A(_804_), .B(_805_), .C(_66__2_), .Y(_806_) );
NAND2X1 NAND2X1_231 ( .A(_806_), .B(_810_), .Y(_64__2_) );
OAI21X1 OAI21X1_231 ( .A(_807_), .B(_804_), .C(_809_), .Y(_66__3_) );
INVX1 INVX1_144 ( .A(_67_), .Y(_811_) );
NAND2X1 NAND2X1_232 ( .A(_68_), .B(w_cout_11_), .Y(_812_) );
OAI21X1 OAI21X1_232 ( .A(w_cout_11_), .B(_811_), .C(_812_), .Y(w_cout_12_) );
INVX1 INVX1_145 ( .A(_69__0_), .Y(_813_) );
NAND2X1 NAND2X1_233 ( .A(_70__0_), .B(w_cout_11_), .Y(_814_) );
OAI21X1 OAI21X1_233 ( .A(w_cout_11_), .B(_813_), .C(_814_), .Y(_0__48_) );
INVX1 INVX1_146 ( .A(_69__1_), .Y(_815_) );
NAND2X1 NAND2X1_234 ( .A(w_cout_11_), .B(_70__1_), .Y(_816_) );
OAI21X1 OAI21X1_234 ( .A(w_cout_11_), .B(_815_), .C(_816_), .Y(_0__49_) );
INVX1 INVX1_147 ( .A(_69__2_), .Y(_817_) );
NAND2X1 NAND2X1_235 ( .A(w_cout_11_), .B(_70__2_), .Y(_818_) );
OAI21X1 OAI21X1_235 ( .A(w_cout_11_), .B(_817_), .C(_818_), .Y(_0__50_) );
INVX1 INVX1_148 ( .A(_69__3_), .Y(_819_) );
NAND2X1 NAND2X1_236 ( .A(w_cout_11_), .B(_70__3_), .Y(_820_) );
OAI21X1 OAI21X1_236 ( .A(w_cout_11_), .B(_819_), .C(_820_), .Y(_0__51_) );
INVX1 INVX1_149 ( .A(1'b0), .Y(_824_) );
OR2X2 OR2X2_89 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_825_) );
NAND2X1 NAND2X1_237 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_826_) );
NAND3X1 NAND3X1_89 ( .A(_824_), .B(_826_), .C(_825_), .Y(_827_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_821_) );
AND2X2 AND2X2_89 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_822_) );
OAI21X1 OAI21X1_237 ( .A(_821_), .B(_822_), .C(1'b0), .Y(_823_) );
NAND2X1 NAND2X1_238 ( .A(_823_), .B(_827_), .Y(_69__0_) );
OAI21X1 OAI21X1_238 ( .A(_824_), .B(_821_), .C(_826_), .Y(_71__1_) );
INVX1 INVX1_150 ( .A(_71__3_), .Y(_831_) );
OR2X2 OR2X2_90 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_832_) );
NAND2X1 NAND2X1_239 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_833_) );
NAND3X1 NAND3X1_90 ( .A(_831_), .B(_833_), .C(_832_), .Y(_834_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_828_) );
AND2X2 AND2X2_90 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_829_) );
OAI21X1 OAI21X1_239 ( .A(_828_), .B(_829_), .C(_71__3_), .Y(_830_) );
NAND2X1 NAND2X1_240 ( .A(_830_), .B(_834_), .Y(_69__3_) );
OAI21X1 OAI21X1_240 ( .A(_831_), .B(_828_), .C(_833_), .Y(_67_) );
INVX1 INVX1_151 ( .A(_71__1_), .Y(_838_) );
OR2X2 OR2X2_91 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_839_) );
NAND2X1 NAND2X1_241 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_840_) );
NAND3X1 NAND3X1_91 ( .A(_838_), .B(_840_), .C(_839_), .Y(_841_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_835_) );
AND2X2 AND2X2_91 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_836_) );
OAI21X1 OAI21X1_241 ( .A(_835_), .B(_836_), .C(_71__1_), .Y(_837_) );
NAND2X1 NAND2X1_242 ( .A(_837_), .B(_841_), .Y(_69__1_) );
OAI21X1 OAI21X1_242 ( .A(_838_), .B(_835_), .C(_840_), .Y(_71__2_) );
INVX1 INVX1_152 ( .A(_71__2_), .Y(_845_) );
OR2X2 OR2X2_92 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_846_) );
NAND2X1 NAND2X1_243 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_847_) );
NAND3X1 NAND3X1_92 ( .A(_845_), .B(_847_), .C(_846_), .Y(_848_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_842_) );
AND2X2 AND2X2_92 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_843_) );
OAI21X1 OAI21X1_243 ( .A(_842_), .B(_843_), .C(_71__2_), .Y(_844_) );
NAND2X1 NAND2X1_244 ( .A(_844_), .B(_848_), .Y(_69__2_) );
OAI21X1 OAI21X1_244 ( .A(_845_), .B(_842_), .C(_847_), .Y(_71__3_) );
INVX1 INVX1_153 ( .A(1'b1), .Y(_852_) );
OR2X2 OR2X2_93 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_853_) );
NAND2X1 NAND2X1_245 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_854_) );
NAND3X1 NAND3X1_93 ( .A(_852_), .B(_854_), .C(_853_), .Y(_855_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_849_) );
AND2X2 AND2X2_93 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_850_) );
OAI21X1 OAI21X1_245 ( .A(_849_), .B(_850_), .C(1'b1), .Y(_851_) );
NAND2X1 NAND2X1_246 ( .A(_851_), .B(_855_), .Y(_70__0_) );
OAI21X1 OAI21X1_246 ( .A(_852_), .B(_849_), .C(_854_), .Y(_72__1_) );
INVX1 INVX1_154 ( .A(_72__3_), .Y(_859_) );
OR2X2 OR2X2_94 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_860_) );
NAND2X1 NAND2X1_247 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_861_) );
NAND3X1 NAND3X1_94 ( .A(_859_), .B(_861_), .C(_860_), .Y(_862_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_856_) );
AND2X2 AND2X2_94 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_857_) );
OAI21X1 OAI21X1_247 ( .A(_856_), .B(_857_), .C(_72__3_), .Y(_858_) );
NAND2X1 NAND2X1_248 ( .A(_858_), .B(_862_), .Y(_70__3_) );
OAI21X1 OAI21X1_248 ( .A(_859_), .B(_856_), .C(_861_), .Y(_68_) );
INVX1 INVX1_155 ( .A(_72__1_), .Y(_866_) );
OR2X2 OR2X2_95 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_867_) );
NAND2X1 NAND2X1_249 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_868_) );
NAND3X1 NAND3X1_95 ( .A(_866_), .B(_868_), .C(_867_), .Y(_869_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_863_) );
AND2X2 AND2X2_95 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_864_) );
OAI21X1 OAI21X1_249 ( .A(_863_), .B(_864_), .C(_72__1_), .Y(_865_) );
NAND2X1 NAND2X1_250 ( .A(_865_), .B(_869_), .Y(_70__1_) );
OAI21X1 OAI21X1_250 ( .A(_866_), .B(_863_), .C(_868_), .Y(_72__2_) );
INVX1 INVX1_156 ( .A(_72__2_), .Y(_873_) );
OR2X2 OR2X2_96 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_874_) );
NAND2X1 NAND2X1_251 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_875_) );
NAND3X1 NAND3X1_96 ( .A(_873_), .B(_875_), .C(_874_), .Y(_876_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_870_) );
AND2X2 AND2X2_96 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_871_) );
OAI21X1 OAI21X1_251 ( .A(_870_), .B(_871_), .C(_72__2_), .Y(_872_) );
NAND2X1 NAND2X1_252 ( .A(_872_), .B(_876_), .Y(_70__2_) );
OAI21X1 OAI21X1_252 ( .A(_873_), .B(_870_), .C(_875_), .Y(_72__3_) );
INVX1 INVX1_157 ( .A(_73_), .Y(_877_) );
NAND2X1 NAND2X1_253 ( .A(_74_), .B(w_cout_12_), .Y(_878_) );
OAI21X1 OAI21X1_253 ( .A(w_cout_12_), .B(_877_), .C(_878_), .Y(w_cout_13_) );
INVX1 INVX1_158 ( .A(_75__0_), .Y(_879_) );
NAND2X1 NAND2X1_254 ( .A(_76__0_), .B(w_cout_12_), .Y(_880_) );
OAI21X1 OAI21X1_254 ( .A(w_cout_12_), .B(_879_), .C(_880_), .Y(_0__52_) );
INVX1 INVX1_159 ( .A(_75__1_), .Y(_881_) );
NAND2X1 NAND2X1_255 ( .A(w_cout_12_), .B(_76__1_), .Y(_882_) );
OAI21X1 OAI21X1_255 ( .A(w_cout_12_), .B(_881_), .C(_882_), .Y(_0__53_) );
INVX1 INVX1_160 ( .A(_75__2_), .Y(_883_) );
NAND2X1 NAND2X1_256 ( .A(w_cout_12_), .B(_76__2_), .Y(_884_) );
OAI21X1 OAI21X1_256 ( .A(w_cout_12_), .B(_883_), .C(_884_), .Y(_0__54_) );
INVX1 INVX1_161 ( .A(_75__3_), .Y(_885_) );
NAND2X1 NAND2X1_257 ( .A(w_cout_12_), .B(_76__3_), .Y(_886_) );
OAI21X1 OAI21X1_257 ( .A(w_cout_12_), .B(_885_), .C(_886_), .Y(_0__55_) );
INVX1 INVX1_162 ( .A(1'b0), .Y(_890_) );
OR2X2 OR2X2_97 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_891_) );
NAND2X1 NAND2X1_258 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_892_) );
NAND3X1 NAND3X1_97 ( .A(_890_), .B(_892_), .C(_891_), .Y(_893_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_887_) );
AND2X2 AND2X2_97 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_888_) );
OAI21X1 OAI21X1_258 ( .A(_887_), .B(_888_), .C(1'b0), .Y(_889_) );
NAND2X1 NAND2X1_259 ( .A(_889_), .B(_893_), .Y(_75__0_) );
OAI21X1 OAI21X1_259 ( .A(_890_), .B(_887_), .C(_892_), .Y(_77__1_) );
INVX1 INVX1_163 ( .A(_77__3_), .Y(_897_) );
OR2X2 OR2X2_98 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_898_) );
NAND2X1 NAND2X1_260 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_899_) );
NAND3X1 NAND3X1_98 ( .A(_897_), .B(_899_), .C(_898_), .Y(_900_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_894_) );
AND2X2 AND2X2_98 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_895_) );
OAI21X1 OAI21X1_260 ( .A(_894_), .B(_895_), .C(_77__3_), .Y(_896_) );
NAND2X1 NAND2X1_261 ( .A(_896_), .B(_900_), .Y(_75__3_) );
OAI21X1 OAI21X1_261 ( .A(_897_), .B(_894_), .C(_899_), .Y(_73_) );
INVX1 INVX1_164 ( .A(_77__1_), .Y(_904_) );
OR2X2 OR2X2_99 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_905_) );
NAND2X1 NAND2X1_262 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_906_) );
NAND3X1 NAND3X1_99 ( .A(_904_), .B(_906_), .C(_905_), .Y(_907_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_901_) );
AND2X2 AND2X2_99 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_902_) );
OAI21X1 OAI21X1_262 ( .A(_901_), .B(_902_), .C(_77__1_), .Y(_903_) );
NAND2X1 NAND2X1_263 ( .A(_903_), .B(_907_), .Y(_75__1_) );
OAI21X1 OAI21X1_263 ( .A(_904_), .B(_901_), .C(_906_), .Y(_77__2_) );
INVX1 INVX1_165 ( .A(_77__2_), .Y(_911_) );
OR2X2 OR2X2_100 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_912_) );
NAND2X1 NAND2X1_264 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_913_) );
NAND3X1 NAND3X1_100 ( .A(_911_), .B(_913_), .C(_912_), .Y(_914_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_908_) );
AND2X2 AND2X2_100 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_909_) );
OAI21X1 OAI21X1_264 ( .A(_908_), .B(_909_), .C(_77__2_), .Y(_910_) );
NAND2X1 NAND2X1_265 ( .A(_910_), .B(_914_), .Y(_75__2_) );
OAI21X1 OAI21X1_265 ( .A(_911_), .B(_908_), .C(_913_), .Y(_77__3_) );
INVX1 INVX1_166 ( .A(1'b1), .Y(_918_) );
OR2X2 OR2X2_101 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_919_) );
NAND2X1 NAND2X1_266 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_920_) );
NAND3X1 NAND3X1_101 ( .A(_918_), .B(_920_), .C(_919_), .Y(_921_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_915_) );
AND2X2 AND2X2_101 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_916_) );
OAI21X1 OAI21X1_266 ( .A(_915_), .B(_916_), .C(1'b1), .Y(_917_) );
NAND2X1 NAND2X1_267 ( .A(_917_), .B(_921_), .Y(_76__0_) );
OAI21X1 OAI21X1_267 ( .A(_918_), .B(_915_), .C(_920_), .Y(_78__1_) );
INVX1 INVX1_167 ( .A(_78__3_), .Y(_925_) );
OR2X2 OR2X2_102 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_926_) );
NAND2X1 NAND2X1_268 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_927_) );
NAND3X1 NAND3X1_102 ( .A(_925_), .B(_927_), .C(_926_), .Y(_928_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_922_) );
AND2X2 AND2X2_102 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_923_) );
OAI21X1 OAI21X1_268 ( .A(_922_), .B(_923_), .C(_78__3_), .Y(_924_) );
NAND2X1 NAND2X1_269 ( .A(_924_), .B(_928_), .Y(_76__3_) );
OAI21X1 OAI21X1_269 ( .A(_925_), .B(_922_), .C(_927_), .Y(_74_) );
INVX1 INVX1_168 ( .A(_78__1_), .Y(_932_) );
OR2X2 OR2X2_103 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_933_) );
NAND2X1 NAND2X1_270 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_934_) );
NAND3X1 NAND3X1_103 ( .A(_932_), .B(_934_), .C(_933_), .Y(_935_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_929_) );
AND2X2 AND2X2_103 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_930_) );
OAI21X1 OAI21X1_270 ( .A(_929_), .B(_930_), .C(_78__1_), .Y(_931_) );
NAND2X1 NAND2X1_271 ( .A(_931_), .B(_935_), .Y(_76__1_) );
OAI21X1 OAI21X1_271 ( .A(_932_), .B(_929_), .C(_934_), .Y(_78__2_) );
INVX1 INVX1_169 ( .A(_78__2_), .Y(_939_) );
OR2X2 OR2X2_104 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_940_) );
NAND2X1 NAND2X1_272 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_941_) );
NAND3X1 NAND3X1_104 ( .A(_939_), .B(_941_), .C(_940_), .Y(_942_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_936_) );
AND2X2 AND2X2_104 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_937_) );
OAI21X1 OAI21X1_272 ( .A(_936_), .B(_937_), .C(_78__2_), .Y(_938_) );
NAND2X1 NAND2X1_273 ( .A(_938_), .B(_942_), .Y(_76__2_) );
OAI21X1 OAI21X1_273 ( .A(_939_), .B(_936_), .C(_941_), .Y(_78__3_) );
INVX1 INVX1_170 ( .A(_79_), .Y(_943_) );
NAND2X1 NAND2X1_274 ( .A(_80_), .B(w_cout_13_), .Y(_944_) );
OAI21X1 OAI21X1_274 ( .A(w_cout_13_), .B(_943_), .C(_944_), .Y(w_cout_14_) );
INVX1 INVX1_171 ( .A(_81__0_), .Y(_945_) );
NAND2X1 NAND2X1_275 ( .A(_82__0_), .B(w_cout_13_), .Y(_946_) );
OAI21X1 OAI21X1_275 ( .A(w_cout_13_), .B(_945_), .C(_946_), .Y(_0__56_) );
INVX1 INVX1_172 ( .A(_81__1_), .Y(_947_) );
NAND2X1 NAND2X1_276 ( .A(w_cout_13_), .B(_82__1_), .Y(_948_) );
OAI21X1 OAI21X1_276 ( .A(w_cout_13_), .B(_947_), .C(_948_), .Y(_0__57_) );
INVX1 INVX1_173 ( .A(_81__2_), .Y(_949_) );
NAND2X1 NAND2X1_277 ( .A(w_cout_13_), .B(_82__2_), .Y(_950_) );
OAI21X1 OAI21X1_277 ( .A(w_cout_13_), .B(_949_), .C(_950_), .Y(_0__58_) );
INVX1 INVX1_174 ( .A(_81__3_), .Y(_951_) );
NAND2X1 NAND2X1_278 ( .A(w_cout_13_), .B(_82__3_), .Y(_952_) );
OAI21X1 OAI21X1_278 ( .A(w_cout_13_), .B(_951_), .C(_952_), .Y(_0__59_) );
INVX1 INVX1_175 ( .A(1'b0), .Y(_956_) );
OR2X2 OR2X2_105 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_957_) );
NAND2X1 NAND2X1_279 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_958_) );
NAND3X1 NAND3X1_105 ( .A(_956_), .B(_958_), .C(_957_), .Y(_959_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_953_) );
AND2X2 AND2X2_105 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_954_) );
OAI21X1 OAI21X1_279 ( .A(_953_), .B(_954_), .C(1'b0), .Y(_955_) );
NAND2X1 NAND2X1_280 ( .A(_955_), .B(_959_), .Y(_81__0_) );
OAI21X1 OAI21X1_280 ( .A(_956_), .B(_953_), .C(_958_), .Y(_83__1_) );
INVX1 INVX1_176 ( .A(_83__3_), .Y(_963_) );
OR2X2 OR2X2_106 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_964_) );
NAND2X1 NAND2X1_281 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_965_) );
NAND3X1 NAND3X1_106 ( .A(_963_), .B(_965_), .C(_964_), .Y(_966_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_960_) );
AND2X2 AND2X2_106 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_961_) );
OAI21X1 OAI21X1_281 ( .A(_960_), .B(_961_), .C(_83__3_), .Y(_962_) );
NAND2X1 NAND2X1_282 ( .A(_962_), .B(_966_), .Y(_81__3_) );
OAI21X1 OAI21X1_282 ( .A(_963_), .B(_960_), .C(_965_), .Y(_79_) );
INVX1 INVX1_177 ( .A(_83__1_), .Y(_970_) );
OR2X2 OR2X2_107 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_971_) );
NAND2X1 NAND2X1_283 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_972_) );
NAND3X1 NAND3X1_107 ( .A(_970_), .B(_972_), .C(_971_), .Y(_973_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_967_) );
AND2X2 AND2X2_107 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_968_) );
OAI21X1 OAI21X1_283 ( .A(_967_), .B(_968_), .C(_83__1_), .Y(_969_) );
NAND2X1 NAND2X1_284 ( .A(_969_), .B(_973_), .Y(_81__1_) );
OAI21X1 OAI21X1_284 ( .A(_970_), .B(_967_), .C(_972_), .Y(_83__2_) );
INVX1 INVX1_178 ( .A(_83__2_), .Y(_977_) );
OR2X2 OR2X2_108 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_978_) );
NAND2X1 NAND2X1_285 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_979_) );
NAND3X1 NAND3X1_108 ( .A(_977_), .B(_979_), .C(_978_), .Y(_980_) );
NOR2X1 NOR2X1_108 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_974_) );
AND2X2 AND2X2_108 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_975_) );
OAI21X1 OAI21X1_285 ( .A(_974_), .B(_975_), .C(_83__2_), .Y(_976_) );
NAND2X1 NAND2X1_286 ( .A(_976_), .B(_980_), .Y(_81__2_) );
OAI21X1 OAI21X1_286 ( .A(_977_), .B(_974_), .C(_979_), .Y(_83__3_) );
INVX1 INVX1_179 ( .A(1'b1), .Y(_984_) );
OR2X2 OR2X2_109 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_985_) );
NAND2X1 NAND2X1_287 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_986_) );
NAND3X1 NAND3X1_109 ( .A(_984_), .B(_986_), .C(_985_), .Y(_987_) );
NOR2X1 NOR2X1_109 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_981_) );
AND2X2 AND2X2_109 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_982_) );
OAI21X1 OAI21X1_287 ( .A(_981_), .B(_982_), .C(1'b1), .Y(_983_) );
NAND2X1 NAND2X1_288 ( .A(_983_), .B(_987_), .Y(_82__0_) );
OAI21X1 OAI21X1_288 ( .A(_984_), .B(_981_), .C(_986_), .Y(_84__1_) );
INVX1 INVX1_180 ( .A(_84__3_), .Y(_991_) );
OR2X2 OR2X2_110 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_992_) );
NAND2X1 NAND2X1_289 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_993_) );
NAND3X1 NAND3X1_110 ( .A(_991_), .B(_993_), .C(_992_), .Y(_994_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_988_) );
AND2X2 AND2X2_110 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_989_) );
OAI21X1 OAI21X1_289 ( .A(_988_), .B(_989_), .C(_84__3_), .Y(_990_) );
NAND2X1 NAND2X1_290 ( .A(_990_), .B(_994_), .Y(_82__3_) );
OAI21X1 OAI21X1_290 ( .A(_991_), .B(_988_), .C(_993_), .Y(_80_) );
INVX1 INVX1_181 ( .A(_84__1_), .Y(_998_) );
OR2X2 OR2X2_111 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_999_) );
NAND2X1 NAND2X1_291 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_1000_) );
NAND3X1 NAND3X1_111 ( .A(_998_), .B(_1000_), .C(_999_), .Y(_1001_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_995_) );
AND2X2 AND2X2_111 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_996_) );
OAI21X1 OAI21X1_291 ( .A(_995_), .B(_996_), .C(_84__1_), .Y(_997_) );
NAND2X1 NAND2X1_292 ( .A(_997_), .B(_1001_), .Y(_82__1_) );
OAI21X1 OAI21X1_292 ( .A(_998_), .B(_995_), .C(_1000_), .Y(_84__2_) );
INVX1 INVX1_182 ( .A(_84__2_), .Y(_1005_) );
OR2X2 OR2X2_112 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1006_) );
NAND2X1 NAND2X1_293 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1007_) );
NAND3X1 NAND3X1_112 ( .A(_1005_), .B(_1007_), .C(_1006_), .Y(_1008_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1002_) );
AND2X2 AND2X2_112 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1003_) );
OAI21X1 OAI21X1_293 ( .A(_1002_), .B(_1003_), .C(_84__2_), .Y(_1004_) );
NAND2X1 NAND2X1_294 ( .A(_1004_), .B(_1008_), .Y(_82__2_) );
OAI21X1 OAI21X1_294 ( .A(_1005_), .B(_1002_), .C(_1007_), .Y(_84__3_) );
INVX1 INVX1_183 ( .A(1'b0), .Y(_1012_) );
OR2X2 OR2X2_113 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1013_) );
NAND2X1 NAND2X1_295 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1014_) );
NAND3X1 NAND3X1_113 ( .A(_1012_), .B(_1014_), .C(_1013_), .Y(_1015_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1009_) );
AND2X2 AND2X2_113 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1010_) );
OAI21X1 OAI21X1_295 ( .A(_1009_), .B(_1010_), .C(1'b0), .Y(_1011_) );
NAND2X1 NAND2X1_296 ( .A(_1011_), .B(_1015_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_296 ( .A(_1012_), .B(_1009_), .C(_1014_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_184 ( .A(rca_inst_fa3_i_carry), .Y(_1019_) );
OR2X2 OR2X2_114 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_1020_) );
NAND2X1 NAND2X1_297 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_1021_) );
NAND3X1 NAND3X1_114 ( .A(_1019_), .B(_1021_), .C(_1020_), .Y(_1022_) );
NOR2X1 NOR2X1_114 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_1016_) );
AND2X2 AND2X2_114 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_1017_) );
OAI21X1 OAI21X1_297 ( .A(_1016_), .B(_1017_), .C(rca_inst_fa3_i_carry), .Y(_1018_) );
NAND2X1 NAND2X1_298 ( .A(_1018_), .B(_1022_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_298 ( .A(_1019_), .B(_1016_), .C(_1021_), .Y(rca_inst_cout) );
INVX1 INVX1_185 ( .A(rca_inst_fa0_o_carry), .Y(_1026_) );
OR2X2 OR2X2_115 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1027_) );
NAND2X1 NAND2X1_299 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1028_) );
NAND3X1 NAND3X1_115 ( .A(_1026_), .B(_1028_), .C(_1027_), .Y(_1029_) );
NOR2X1 NOR2X1_115 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1023_) );
AND2X2 AND2X2_115 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1024_) );
OAI21X1 OAI21X1_299 ( .A(_1023_), .B(_1024_), .C(rca_inst_fa0_o_carry), .Y(_1025_) );
NAND2X1 NAND2X1_300 ( .A(_1025_), .B(_1029_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_300 ( .A(_1026_), .B(_1023_), .C(_1028_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_186 ( .A(rca_inst_fa_1__o_carry), .Y(_1033_) );
OR2X2 OR2X2_116 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1034_) );
NAND2X1 NAND2X1_301 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1035_) );
NAND3X1 NAND3X1_116 ( .A(_1033_), .B(_1035_), .C(_1034_), .Y(_1036_) );
NOR2X1 NOR2X1_116 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1030_) );
AND2X2 AND2X2_116 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1031_) );
OAI21X1 OAI21X1_301 ( .A(_1030_), .B(_1031_), .C(rca_inst_fa_1__o_carry), .Y(_1032_) );
NAND2X1 NAND2X1_302 ( .A(_1032_), .B(_1036_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_302 ( .A(_1033_), .B(_1030_), .C(_1035_), .Y(rca_inst_fa3_i_carry) );
BUFX2 BUFX2_62 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_63 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_64 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_65 ( .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_66 ( .A(rca_inst_cout), .Y(w_cout_0_) );
endmodule
