module CSkipA_51bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term1[45], i_add_term1[46], i_add_term1[47], i_add_term1[48], i_add_term1[49], i_add_term1[50], i_add_term1[51], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], i_add_term2[45], i_add_term2[46], i_add_term2[47], i_add_term2[48], i_add_term2[49], i_add_term2[50], i_add_term2[51], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], sum[45], sum[46], sum[47], sum[48], sum[49], sum[50], sum[51], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term1[45];
input i_add_term1[46];
input i_add_term1[47];
input i_add_term1[48];
input i_add_term1[49];
input i_add_term1[50];
input i_add_term1[51];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
input i_add_term2[45];
input i_add_term2[46];
input i_add_term2[47];
input i_add_term2[48];
input i_add_term2[49];
input i_add_term2[50];
input i_add_term2[51];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output sum[45];
output sum[46];
output sum[47];
output sum[48];
output sum[49];
output sum[50];
output sum[51];
output cout;

INVX1 INVX1_1 ( .A(w_cout_11_), .Y(_408_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_409_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_410_) );
NAND3X1 NAND3X1_1 ( .A(_408_), .B(_410_), .C(_409_), .Y(_411_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_405_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_406_) );
OAI21X1 OAI21X1_1 ( .A(_405_), .B(_406_), .C(w_cout_11_), .Y(_407_) );
NAND2X1 NAND2X1_2 ( .A(_407_), .B(_411_), .Y(_0__48_) );
OAI21X1 OAI21X1_2 ( .A(_408_), .B(_405_), .C(_410_), .Y(_24__1_) );
INVX1 INVX1_2 ( .A(_24__1_), .Y(_415_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_416_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_417_) );
NAND3X1 NAND3X1_2 ( .A(_415_), .B(_417_), .C(_416_), .Y(_418_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_412_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_413_) );
OAI21X1 OAI21X1_3 ( .A(_412_), .B(_413_), .C(_24__1_), .Y(_414_) );
NAND2X1 NAND2X1_4 ( .A(_414_), .B(_418_), .Y(_0__49_) );
OAI21X1 OAI21X1_4 ( .A(_415_), .B(_412_), .C(_417_), .Y(_24__2_) );
INVX1 INVX1_3 ( .A(_24__2_), .Y(_422_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_423_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_424_) );
NAND3X1 NAND3X1_3 ( .A(_422_), .B(_424_), .C(_423_), .Y(_425_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_419_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_420_) );
OAI21X1 OAI21X1_5 ( .A(_419_), .B(_420_), .C(_24__2_), .Y(_421_) );
NAND2X1 NAND2X1_6 ( .A(_421_), .B(_425_), .Y(_0__50_) );
OAI21X1 OAI21X1_6 ( .A(_422_), .B(_419_), .C(_424_), .Y(_24__3_) );
INVX1 INVX1_4 ( .A(_24__3_), .Y(_429_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_430_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_431_) );
NAND3X1 NAND3X1_4 ( .A(_429_), .B(_431_), .C(_430_), .Y(_432_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_426_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_427_) );
OAI21X1 OAI21X1_7 ( .A(_426_), .B(_427_), .C(_24__3_), .Y(_428_) );
NAND2X1 NAND2X1_8 ( .A(_428_), .B(_432_), .Y(_0__51_) );
OAI21X1 OAI21X1_8 ( .A(_429_), .B(_426_), .C(_431_), .Y(_23_) );
INVX1 INVX1_5 ( .A(1'b0), .Y(_436_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_437_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_438_) );
NAND3X1 NAND3X1_5 ( .A(_436_), .B(_438_), .C(_437_), .Y(_439_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_433_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_434_) );
OAI21X1 OAI21X1_9 ( .A(_433_), .B(_434_), .C(1'b0), .Y(_435_) );
NAND2X1 NAND2X1_10 ( .A(_435_), .B(_439_), .Y(_0__0_) );
OAI21X1 OAI21X1_10 ( .A(_436_), .B(_433_), .C(_438_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_6 ( .A(rca_inst_w_CARRY_1_), .Y(_443_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_444_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_445_) );
NAND3X1 NAND3X1_6 ( .A(_443_), .B(_445_), .C(_444_), .Y(_446_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_440_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_441_) );
OAI21X1 OAI21X1_11 ( .A(_440_), .B(_441_), .C(rca_inst_w_CARRY_1_), .Y(_442_) );
NAND2X1 NAND2X1_12 ( .A(_442_), .B(_446_), .Y(_0__1_) );
OAI21X1 OAI21X1_12 ( .A(_443_), .B(_440_), .C(_445_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_7 ( .A(rca_inst_w_CARRY_2_), .Y(_450_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_451_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_452_) );
NAND3X1 NAND3X1_7 ( .A(_450_), .B(_452_), .C(_451_), .Y(_453_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_447_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_448_) );
OAI21X1 OAI21X1_13 ( .A(_447_), .B(_448_), .C(rca_inst_w_CARRY_2_), .Y(_449_) );
NAND2X1 NAND2X1_14 ( .A(_449_), .B(_453_), .Y(_0__2_) );
OAI21X1 OAI21X1_14 ( .A(_450_), .B(_447_), .C(_452_), .Y(rca_inst_w_CARRY_3_) );
INVX1 INVX1_8 ( .A(rca_inst_w_CARRY_3_), .Y(_457_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_458_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_459_) );
NAND3X1 NAND3X1_8 ( .A(_457_), .B(_459_), .C(_458_), .Y(_460_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_454_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_455_) );
OAI21X1 OAI21X1_15 ( .A(_454_), .B(_455_), .C(rca_inst_w_CARRY_3_), .Y(_456_) );
NAND2X1 NAND2X1_16 ( .A(_456_), .B(_460_), .Y(_0__3_) );
OAI21X1 OAI21X1_16 ( .A(_457_), .B(_454_), .C(_459_), .Y(cout0) );
INVX1 INVX1_9 ( .A(cout0), .Y(_461_) );
OAI21X1 OAI21X1_17 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .C(1'b0), .Y(_462_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_463_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_464_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_465_) );
NAND3X1 NAND3X1_9 ( .A(_463_), .B(_464_), .C(_465_), .Y(_466_) );
OAI21X1 OAI21X1_18 ( .A(_462_), .B(_466_), .C(_461_), .Y(skip0_cin_next) );
BUFX2 BUFX2_1 ( .A(w_cout_12_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
INVX1 INVX1_10 ( .A(_1_), .Y(_25_) );
OAI21X1 OAI21X1_19 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .C(1'b0), .Y(_26_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_27_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_28_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_29_) );
NAND3X1 NAND3X1_10 ( .A(_27_), .B(_28_), .C(_29_), .Y(_30_) );
OAI21X1 OAI21X1_20 ( .A(_26_), .B(_30_), .C(_25_), .Y(w_cout_1_) );
INVX1 INVX1_11 ( .A(_3_), .Y(_31_) );
OAI21X1 OAI21X1_21 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .C(1'b0), .Y(_32_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_33_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_34_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_35_) );
NAND3X1 NAND3X1_11 ( .A(_33_), .B(_34_), .C(_35_), .Y(_36_) );
OAI21X1 OAI21X1_22 ( .A(_32_), .B(_36_), .C(_31_), .Y(w_cout_2_) );
INVX1 INVX1_12 ( .A(_5_), .Y(_37_) );
OAI21X1 OAI21X1_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .C(1'b0), .Y(_38_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_39_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_40_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_41_) );
NAND3X1 NAND3X1_12 ( .A(_39_), .B(_40_), .C(_41_), .Y(_42_) );
OAI21X1 OAI21X1_24 ( .A(_38_), .B(_42_), .C(_37_), .Y(w_cout_3_) );
INVX1 INVX1_13 ( .A(_7_), .Y(_43_) );
OAI21X1 OAI21X1_25 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .C(1'b0), .Y(_44_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_45_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_46_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_47_) );
NAND3X1 NAND3X1_13 ( .A(_45_), .B(_46_), .C(_47_), .Y(_48_) );
OAI21X1 OAI21X1_26 ( .A(_44_), .B(_48_), .C(_43_), .Y(w_cout_4_) );
INVX1 INVX1_14 ( .A(_9_), .Y(_49_) );
OAI21X1 OAI21X1_27 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .C(1'b0), .Y(_50_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_51_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_52_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_53_) );
NAND3X1 NAND3X1_14 ( .A(_51_), .B(_52_), .C(_53_), .Y(_54_) );
OAI21X1 OAI21X1_28 ( .A(_50_), .B(_54_), .C(_49_), .Y(w_cout_5_) );
INVX1 INVX1_15 ( .A(_11_), .Y(_55_) );
OAI21X1 OAI21X1_29 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .C(1'b0), .Y(_56_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_57_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_58_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_59_) );
NAND3X1 NAND3X1_15 ( .A(_57_), .B(_58_), .C(_59_), .Y(_60_) );
OAI21X1 OAI21X1_30 ( .A(_56_), .B(_60_), .C(_55_), .Y(w_cout_6_) );
INVX1 INVX1_16 ( .A(_13_), .Y(_61_) );
OAI21X1 OAI21X1_31 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .C(1'b0), .Y(_62_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_63_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_64_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_65_) );
NAND3X1 NAND3X1_16 ( .A(_63_), .B(_64_), .C(_65_), .Y(_66_) );
OAI21X1 OAI21X1_32 ( .A(_62_), .B(_66_), .C(_61_), .Y(w_cout_7_) );
INVX1 INVX1_17 ( .A(_15_), .Y(_67_) );
OAI21X1 OAI21X1_33 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .C(1'b0), .Y(_68_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_69_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_70_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_71_) );
NAND3X1 NAND3X1_17 ( .A(_69_), .B(_70_), .C(_71_), .Y(_72_) );
OAI21X1 OAI21X1_34 ( .A(_68_), .B(_72_), .C(_67_), .Y(w_cout_8_) );
INVX1 INVX1_18 ( .A(_17_), .Y(_73_) );
OAI21X1 OAI21X1_35 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .C(1'b0), .Y(_74_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_75_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_76_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_77_) );
NAND3X1 NAND3X1_18 ( .A(_75_), .B(_76_), .C(_77_), .Y(_78_) );
OAI21X1 OAI21X1_36 ( .A(_74_), .B(_78_), .C(_73_), .Y(w_cout_9_) );
INVX1 INVX1_19 ( .A(_19_), .Y(_79_) );
OAI21X1 OAI21X1_37 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .C(1'b0), .Y(_80_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_81_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_82_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_83_) );
NAND3X1 NAND3X1_19 ( .A(_81_), .B(_82_), .C(_83_), .Y(_84_) );
OAI21X1 OAI21X1_38 ( .A(_80_), .B(_84_), .C(_79_), .Y(w_cout_10_) );
INVX1 INVX1_20 ( .A(_21_), .Y(_85_) );
OAI21X1 OAI21X1_39 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .C(1'b0), .Y(_86_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_87_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_88_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_89_) );
NAND3X1 NAND3X1_20 ( .A(_87_), .B(_88_), .C(_89_), .Y(_90_) );
OAI21X1 OAI21X1_40 ( .A(_86_), .B(_90_), .C(_85_), .Y(w_cout_11_) );
INVX1 INVX1_21 ( .A(_23_), .Y(_91_) );
OAI21X1 OAI21X1_41 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .C(1'b0), .Y(_92_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_93_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_94_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_95_) );
NAND3X1 NAND3X1_21 ( .A(_93_), .B(_94_), .C(_95_), .Y(_96_) );
OAI21X1 OAI21X1_42 ( .A(_92_), .B(_96_), .C(_91_), .Y(w_cout_12_) );
INVX1 INVX1_22 ( .A(skip0_cin_next), .Y(_100_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_101_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_102_) );
NAND3X1 NAND3X1_22 ( .A(_100_), .B(_102_), .C(_101_), .Y(_103_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_97_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_98_) );
OAI21X1 OAI21X1_43 ( .A(_97_), .B(_98_), .C(skip0_cin_next), .Y(_99_) );
NAND2X1 NAND2X1_18 ( .A(_99_), .B(_103_), .Y(_0__4_) );
OAI21X1 OAI21X1_44 ( .A(_100_), .B(_97_), .C(_102_), .Y(_2__1_) );
INVX1 INVX1_23 ( .A(_2__1_), .Y(_107_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_108_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_109_) );
NAND3X1 NAND3X1_23 ( .A(_107_), .B(_109_), .C(_108_), .Y(_110_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_104_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_105_) );
OAI21X1 OAI21X1_45 ( .A(_104_), .B(_105_), .C(_2__1_), .Y(_106_) );
NAND2X1 NAND2X1_20 ( .A(_106_), .B(_110_), .Y(_0__5_) );
OAI21X1 OAI21X1_46 ( .A(_107_), .B(_104_), .C(_109_), .Y(_2__2_) );
INVX1 INVX1_24 ( .A(_2__2_), .Y(_114_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_115_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_116_) );
NAND3X1 NAND3X1_24 ( .A(_114_), .B(_116_), .C(_115_), .Y(_117_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_111_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_112_) );
OAI21X1 OAI21X1_47 ( .A(_111_), .B(_112_), .C(_2__2_), .Y(_113_) );
NAND2X1 NAND2X1_22 ( .A(_113_), .B(_117_), .Y(_0__6_) );
OAI21X1 OAI21X1_48 ( .A(_114_), .B(_111_), .C(_116_), .Y(_2__3_) );
INVX1 INVX1_25 ( .A(_2__3_), .Y(_121_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_122_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_123_) );
NAND3X1 NAND3X1_25 ( .A(_121_), .B(_123_), .C(_122_), .Y(_124_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_118_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_119_) );
OAI21X1 OAI21X1_49 ( .A(_118_), .B(_119_), .C(_2__3_), .Y(_120_) );
NAND2X1 NAND2X1_24 ( .A(_120_), .B(_124_), .Y(_0__7_) );
OAI21X1 OAI21X1_50 ( .A(_121_), .B(_118_), .C(_123_), .Y(_1_) );
INVX1 INVX1_26 ( .A(w_cout_1_), .Y(_128_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_129_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_130_) );
NAND3X1 NAND3X1_26 ( .A(_128_), .B(_130_), .C(_129_), .Y(_131_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_125_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_126_) );
OAI21X1 OAI21X1_51 ( .A(_125_), .B(_126_), .C(w_cout_1_), .Y(_127_) );
NAND2X1 NAND2X1_26 ( .A(_127_), .B(_131_), .Y(_0__8_) );
OAI21X1 OAI21X1_52 ( .A(_128_), .B(_125_), .C(_130_), .Y(_4__1_) );
INVX1 INVX1_27 ( .A(_4__1_), .Y(_135_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_136_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_137_) );
NAND3X1 NAND3X1_27 ( .A(_135_), .B(_137_), .C(_136_), .Y(_138_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_132_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_133_) );
OAI21X1 OAI21X1_53 ( .A(_132_), .B(_133_), .C(_4__1_), .Y(_134_) );
NAND2X1 NAND2X1_28 ( .A(_134_), .B(_138_), .Y(_0__9_) );
OAI21X1 OAI21X1_54 ( .A(_135_), .B(_132_), .C(_137_), .Y(_4__2_) );
INVX1 INVX1_28 ( .A(_4__2_), .Y(_142_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_143_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_144_) );
NAND3X1 NAND3X1_28 ( .A(_142_), .B(_144_), .C(_143_), .Y(_145_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_139_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_140_) );
OAI21X1 OAI21X1_55 ( .A(_139_), .B(_140_), .C(_4__2_), .Y(_141_) );
NAND2X1 NAND2X1_30 ( .A(_141_), .B(_145_), .Y(_0__10_) );
OAI21X1 OAI21X1_56 ( .A(_142_), .B(_139_), .C(_144_), .Y(_4__3_) );
INVX1 INVX1_29 ( .A(_4__3_), .Y(_149_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_150_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_151_) );
NAND3X1 NAND3X1_29 ( .A(_149_), .B(_151_), .C(_150_), .Y(_152_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_146_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_147_) );
OAI21X1 OAI21X1_57 ( .A(_146_), .B(_147_), .C(_4__3_), .Y(_148_) );
NAND2X1 NAND2X1_32 ( .A(_148_), .B(_152_), .Y(_0__11_) );
OAI21X1 OAI21X1_58 ( .A(_149_), .B(_146_), .C(_151_), .Y(_3_) );
INVX1 INVX1_30 ( .A(w_cout_2_), .Y(_156_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_157_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_158_) );
NAND3X1 NAND3X1_30 ( .A(_156_), .B(_158_), .C(_157_), .Y(_159_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_153_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_154_) );
OAI21X1 OAI21X1_59 ( .A(_153_), .B(_154_), .C(w_cout_2_), .Y(_155_) );
NAND2X1 NAND2X1_34 ( .A(_155_), .B(_159_), .Y(_0__12_) );
OAI21X1 OAI21X1_60 ( .A(_156_), .B(_153_), .C(_158_), .Y(_6__1_) );
INVX1 INVX1_31 ( .A(_6__1_), .Y(_163_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_164_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_165_) );
NAND3X1 NAND3X1_31 ( .A(_163_), .B(_165_), .C(_164_), .Y(_166_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_160_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_161_) );
OAI21X1 OAI21X1_61 ( .A(_160_), .B(_161_), .C(_6__1_), .Y(_162_) );
NAND2X1 NAND2X1_36 ( .A(_162_), .B(_166_), .Y(_0__13_) );
OAI21X1 OAI21X1_62 ( .A(_163_), .B(_160_), .C(_165_), .Y(_6__2_) );
INVX1 INVX1_32 ( .A(_6__2_), .Y(_170_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_171_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_172_) );
NAND3X1 NAND3X1_32 ( .A(_170_), .B(_172_), .C(_171_), .Y(_173_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_167_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_168_) );
OAI21X1 OAI21X1_63 ( .A(_167_), .B(_168_), .C(_6__2_), .Y(_169_) );
NAND2X1 NAND2X1_38 ( .A(_169_), .B(_173_), .Y(_0__14_) );
OAI21X1 OAI21X1_64 ( .A(_170_), .B(_167_), .C(_172_), .Y(_6__3_) );
INVX1 INVX1_33 ( .A(_6__3_), .Y(_177_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_178_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_179_) );
NAND3X1 NAND3X1_33 ( .A(_177_), .B(_179_), .C(_178_), .Y(_180_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_174_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_175_) );
OAI21X1 OAI21X1_65 ( .A(_174_), .B(_175_), .C(_6__3_), .Y(_176_) );
NAND2X1 NAND2X1_40 ( .A(_176_), .B(_180_), .Y(_0__15_) );
OAI21X1 OAI21X1_66 ( .A(_177_), .B(_174_), .C(_179_), .Y(_5_) );
INVX1 INVX1_34 ( .A(w_cout_3_), .Y(_184_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_185_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_186_) );
NAND3X1 NAND3X1_34 ( .A(_184_), .B(_186_), .C(_185_), .Y(_187_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_181_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_182_) );
OAI21X1 OAI21X1_67 ( .A(_181_), .B(_182_), .C(w_cout_3_), .Y(_183_) );
NAND2X1 NAND2X1_42 ( .A(_183_), .B(_187_), .Y(_0__16_) );
OAI21X1 OAI21X1_68 ( .A(_184_), .B(_181_), .C(_186_), .Y(_8__1_) );
INVX1 INVX1_35 ( .A(_8__1_), .Y(_191_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_192_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_193_) );
NAND3X1 NAND3X1_35 ( .A(_191_), .B(_193_), .C(_192_), .Y(_194_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_188_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_189_) );
OAI21X1 OAI21X1_69 ( .A(_188_), .B(_189_), .C(_8__1_), .Y(_190_) );
NAND2X1 NAND2X1_44 ( .A(_190_), .B(_194_), .Y(_0__17_) );
OAI21X1 OAI21X1_70 ( .A(_191_), .B(_188_), .C(_193_), .Y(_8__2_) );
INVX1 INVX1_36 ( .A(_8__2_), .Y(_198_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_199_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_200_) );
NAND3X1 NAND3X1_36 ( .A(_198_), .B(_200_), .C(_199_), .Y(_201_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_195_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_196_) );
OAI21X1 OAI21X1_71 ( .A(_195_), .B(_196_), .C(_8__2_), .Y(_197_) );
NAND2X1 NAND2X1_46 ( .A(_197_), .B(_201_), .Y(_0__18_) );
OAI21X1 OAI21X1_72 ( .A(_198_), .B(_195_), .C(_200_), .Y(_8__3_) );
INVX1 INVX1_37 ( .A(_8__3_), .Y(_205_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_206_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_207_) );
NAND3X1 NAND3X1_37 ( .A(_205_), .B(_207_), .C(_206_), .Y(_208_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_202_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_203_) );
OAI21X1 OAI21X1_73 ( .A(_202_), .B(_203_), .C(_8__3_), .Y(_204_) );
NAND2X1 NAND2X1_48 ( .A(_204_), .B(_208_), .Y(_0__19_) );
OAI21X1 OAI21X1_74 ( .A(_205_), .B(_202_), .C(_207_), .Y(_7_) );
INVX1 INVX1_38 ( .A(w_cout_4_), .Y(_212_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_213_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_214_) );
NAND3X1 NAND3X1_38 ( .A(_212_), .B(_214_), .C(_213_), .Y(_215_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_209_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_210_) );
OAI21X1 OAI21X1_75 ( .A(_209_), .B(_210_), .C(w_cout_4_), .Y(_211_) );
NAND2X1 NAND2X1_50 ( .A(_211_), .B(_215_), .Y(_0__20_) );
OAI21X1 OAI21X1_76 ( .A(_212_), .B(_209_), .C(_214_), .Y(_10__1_) );
INVX1 INVX1_39 ( .A(_10__1_), .Y(_219_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_220_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_221_) );
NAND3X1 NAND3X1_39 ( .A(_219_), .B(_221_), .C(_220_), .Y(_222_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_216_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_217_) );
OAI21X1 OAI21X1_77 ( .A(_216_), .B(_217_), .C(_10__1_), .Y(_218_) );
NAND2X1 NAND2X1_52 ( .A(_218_), .B(_222_), .Y(_0__21_) );
OAI21X1 OAI21X1_78 ( .A(_219_), .B(_216_), .C(_221_), .Y(_10__2_) );
INVX1 INVX1_40 ( .A(_10__2_), .Y(_226_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_227_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_228_) );
NAND3X1 NAND3X1_40 ( .A(_226_), .B(_228_), .C(_227_), .Y(_229_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_223_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_224_) );
OAI21X1 OAI21X1_79 ( .A(_223_), .B(_224_), .C(_10__2_), .Y(_225_) );
NAND2X1 NAND2X1_54 ( .A(_225_), .B(_229_), .Y(_0__22_) );
OAI21X1 OAI21X1_80 ( .A(_226_), .B(_223_), .C(_228_), .Y(_10__3_) );
INVX1 INVX1_41 ( .A(_10__3_), .Y(_233_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_234_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_235_) );
NAND3X1 NAND3X1_41 ( .A(_233_), .B(_235_), .C(_234_), .Y(_236_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_230_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_231_) );
OAI21X1 OAI21X1_81 ( .A(_230_), .B(_231_), .C(_10__3_), .Y(_232_) );
NAND2X1 NAND2X1_56 ( .A(_232_), .B(_236_), .Y(_0__23_) );
OAI21X1 OAI21X1_82 ( .A(_233_), .B(_230_), .C(_235_), .Y(_9_) );
INVX1 INVX1_42 ( .A(w_cout_5_), .Y(_240_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_241_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_242_) );
NAND3X1 NAND3X1_42 ( .A(_240_), .B(_242_), .C(_241_), .Y(_243_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_237_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_238_) );
OAI21X1 OAI21X1_83 ( .A(_237_), .B(_238_), .C(w_cout_5_), .Y(_239_) );
NAND2X1 NAND2X1_58 ( .A(_239_), .B(_243_), .Y(_0__24_) );
OAI21X1 OAI21X1_84 ( .A(_240_), .B(_237_), .C(_242_), .Y(_12__1_) );
INVX1 INVX1_43 ( .A(_12__1_), .Y(_247_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_248_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_249_) );
NAND3X1 NAND3X1_43 ( .A(_247_), .B(_249_), .C(_248_), .Y(_250_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_244_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_245_) );
OAI21X1 OAI21X1_85 ( .A(_244_), .B(_245_), .C(_12__1_), .Y(_246_) );
NAND2X1 NAND2X1_60 ( .A(_246_), .B(_250_), .Y(_0__25_) );
OAI21X1 OAI21X1_86 ( .A(_247_), .B(_244_), .C(_249_), .Y(_12__2_) );
INVX1 INVX1_44 ( .A(_12__2_), .Y(_254_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_255_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_256_) );
NAND3X1 NAND3X1_44 ( .A(_254_), .B(_256_), .C(_255_), .Y(_257_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_251_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_252_) );
OAI21X1 OAI21X1_87 ( .A(_251_), .B(_252_), .C(_12__2_), .Y(_253_) );
NAND2X1 NAND2X1_62 ( .A(_253_), .B(_257_), .Y(_0__26_) );
OAI21X1 OAI21X1_88 ( .A(_254_), .B(_251_), .C(_256_), .Y(_12__3_) );
INVX1 INVX1_45 ( .A(_12__3_), .Y(_261_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_262_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_263_) );
NAND3X1 NAND3X1_45 ( .A(_261_), .B(_263_), .C(_262_), .Y(_264_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_258_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_259_) );
OAI21X1 OAI21X1_89 ( .A(_258_), .B(_259_), .C(_12__3_), .Y(_260_) );
NAND2X1 NAND2X1_64 ( .A(_260_), .B(_264_), .Y(_0__27_) );
OAI21X1 OAI21X1_90 ( .A(_261_), .B(_258_), .C(_263_), .Y(_11_) );
INVX1 INVX1_46 ( .A(w_cout_6_), .Y(_268_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_269_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_270_) );
NAND3X1 NAND3X1_46 ( .A(_268_), .B(_270_), .C(_269_), .Y(_271_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_265_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_266_) );
OAI21X1 OAI21X1_91 ( .A(_265_), .B(_266_), .C(w_cout_6_), .Y(_267_) );
NAND2X1 NAND2X1_66 ( .A(_267_), .B(_271_), .Y(_0__28_) );
OAI21X1 OAI21X1_92 ( .A(_268_), .B(_265_), .C(_270_), .Y(_14__1_) );
INVX1 INVX1_47 ( .A(_14__1_), .Y(_275_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_276_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_277_) );
NAND3X1 NAND3X1_47 ( .A(_275_), .B(_277_), .C(_276_), .Y(_278_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_272_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_273_) );
OAI21X1 OAI21X1_93 ( .A(_272_), .B(_273_), .C(_14__1_), .Y(_274_) );
NAND2X1 NAND2X1_68 ( .A(_274_), .B(_278_), .Y(_0__29_) );
OAI21X1 OAI21X1_94 ( .A(_275_), .B(_272_), .C(_277_), .Y(_14__2_) );
INVX1 INVX1_48 ( .A(_14__2_), .Y(_282_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_283_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_284_) );
NAND3X1 NAND3X1_48 ( .A(_282_), .B(_284_), .C(_283_), .Y(_285_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_279_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_280_) );
OAI21X1 OAI21X1_95 ( .A(_279_), .B(_280_), .C(_14__2_), .Y(_281_) );
NAND2X1 NAND2X1_70 ( .A(_281_), .B(_285_), .Y(_0__30_) );
OAI21X1 OAI21X1_96 ( .A(_282_), .B(_279_), .C(_284_), .Y(_14__3_) );
INVX1 INVX1_49 ( .A(_14__3_), .Y(_289_) );
OR2X2 OR2X2_75 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_290_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_291_) );
NAND3X1 NAND3X1_49 ( .A(_289_), .B(_291_), .C(_290_), .Y(_292_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_286_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_287_) );
OAI21X1 OAI21X1_97 ( .A(_286_), .B(_287_), .C(_14__3_), .Y(_288_) );
NAND2X1 NAND2X1_72 ( .A(_288_), .B(_292_), .Y(_0__31_) );
OAI21X1 OAI21X1_98 ( .A(_289_), .B(_286_), .C(_291_), .Y(_13_) );
INVX1 INVX1_50 ( .A(w_cout_7_), .Y(_296_) );
OR2X2 OR2X2_76 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_297_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_298_) );
NAND3X1 NAND3X1_50 ( .A(_296_), .B(_298_), .C(_297_), .Y(_299_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_293_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_294_) );
OAI21X1 OAI21X1_99 ( .A(_293_), .B(_294_), .C(w_cout_7_), .Y(_295_) );
NAND2X1 NAND2X1_74 ( .A(_295_), .B(_299_), .Y(_0__32_) );
OAI21X1 OAI21X1_100 ( .A(_296_), .B(_293_), .C(_298_), .Y(_16__1_) );
INVX1 INVX1_51 ( .A(_16__1_), .Y(_303_) );
OR2X2 OR2X2_77 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_304_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_305_) );
NAND3X1 NAND3X1_51 ( .A(_303_), .B(_305_), .C(_304_), .Y(_306_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_300_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_301_) );
OAI21X1 OAI21X1_101 ( .A(_300_), .B(_301_), .C(_16__1_), .Y(_302_) );
NAND2X1 NAND2X1_76 ( .A(_302_), .B(_306_), .Y(_0__33_) );
OAI21X1 OAI21X1_102 ( .A(_303_), .B(_300_), .C(_305_), .Y(_16__2_) );
INVX1 INVX1_52 ( .A(_16__2_), .Y(_310_) );
OR2X2 OR2X2_78 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_311_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_312_) );
NAND3X1 NAND3X1_52 ( .A(_310_), .B(_312_), .C(_311_), .Y(_313_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_307_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_308_) );
OAI21X1 OAI21X1_103 ( .A(_307_), .B(_308_), .C(_16__2_), .Y(_309_) );
NAND2X1 NAND2X1_78 ( .A(_309_), .B(_313_), .Y(_0__34_) );
OAI21X1 OAI21X1_104 ( .A(_310_), .B(_307_), .C(_312_), .Y(_16__3_) );
INVX1 INVX1_53 ( .A(_16__3_), .Y(_317_) );
OR2X2 OR2X2_79 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_318_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_319_) );
NAND3X1 NAND3X1_53 ( .A(_317_), .B(_319_), .C(_318_), .Y(_320_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_314_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_315_) );
OAI21X1 OAI21X1_105 ( .A(_314_), .B(_315_), .C(_16__3_), .Y(_316_) );
NAND2X1 NAND2X1_80 ( .A(_316_), .B(_320_), .Y(_0__35_) );
OAI21X1 OAI21X1_106 ( .A(_317_), .B(_314_), .C(_319_), .Y(_15_) );
INVX1 INVX1_54 ( .A(w_cout_8_), .Y(_324_) );
OR2X2 OR2X2_80 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_325_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_326_) );
NAND3X1 NAND3X1_54 ( .A(_324_), .B(_326_), .C(_325_), .Y(_327_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_321_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_322_) );
OAI21X1 OAI21X1_107 ( .A(_321_), .B(_322_), .C(w_cout_8_), .Y(_323_) );
NAND2X1 NAND2X1_82 ( .A(_323_), .B(_327_), .Y(_0__36_) );
OAI21X1 OAI21X1_108 ( .A(_324_), .B(_321_), .C(_326_), .Y(_18__1_) );
INVX1 INVX1_55 ( .A(_18__1_), .Y(_331_) );
OR2X2 OR2X2_81 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_332_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_333_) );
NAND3X1 NAND3X1_55 ( .A(_331_), .B(_333_), .C(_332_), .Y(_334_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_328_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_329_) );
OAI21X1 OAI21X1_109 ( .A(_328_), .B(_329_), .C(_18__1_), .Y(_330_) );
NAND2X1 NAND2X1_84 ( .A(_330_), .B(_334_), .Y(_0__37_) );
OAI21X1 OAI21X1_110 ( .A(_331_), .B(_328_), .C(_333_), .Y(_18__2_) );
INVX1 INVX1_56 ( .A(_18__2_), .Y(_338_) );
OR2X2 OR2X2_82 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_339_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_340_) );
NAND3X1 NAND3X1_56 ( .A(_338_), .B(_340_), .C(_339_), .Y(_341_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_335_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_336_) );
OAI21X1 OAI21X1_111 ( .A(_335_), .B(_336_), .C(_18__2_), .Y(_337_) );
NAND2X1 NAND2X1_86 ( .A(_337_), .B(_341_), .Y(_0__38_) );
OAI21X1 OAI21X1_112 ( .A(_338_), .B(_335_), .C(_340_), .Y(_18__3_) );
INVX1 INVX1_57 ( .A(_18__3_), .Y(_345_) );
OR2X2 OR2X2_83 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_346_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_347_) );
NAND3X1 NAND3X1_57 ( .A(_345_), .B(_347_), .C(_346_), .Y(_348_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_342_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_343_) );
OAI21X1 OAI21X1_113 ( .A(_342_), .B(_343_), .C(_18__3_), .Y(_344_) );
NAND2X1 NAND2X1_88 ( .A(_344_), .B(_348_), .Y(_0__39_) );
OAI21X1 OAI21X1_114 ( .A(_345_), .B(_342_), .C(_347_), .Y(_17_) );
INVX1 INVX1_58 ( .A(w_cout_9_), .Y(_352_) );
OR2X2 OR2X2_84 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_353_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_354_) );
NAND3X1 NAND3X1_58 ( .A(_352_), .B(_354_), .C(_353_), .Y(_355_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_349_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_350_) );
OAI21X1 OAI21X1_115 ( .A(_349_), .B(_350_), .C(w_cout_9_), .Y(_351_) );
NAND2X1 NAND2X1_90 ( .A(_351_), .B(_355_), .Y(_0__40_) );
OAI21X1 OAI21X1_116 ( .A(_352_), .B(_349_), .C(_354_), .Y(_20__1_) );
INVX1 INVX1_59 ( .A(_20__1_), .Y(_359_) );
OR2X2 OR2X2_85 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_360_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_361_) );
NAND3X1 NAND3X1_59 ( .A(_359_), .B(_361_), .C(_360_), .Y(_362_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_356_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_357_) );
OAI21X1 OAI21X1_117 ( .A(_356_), .B(_357_), .C(_20__1_), .Y(_358_) );
NAND2X1 NAND2X1_92 ( .A(_358_), .B(_362_), .Y(_0__41_) );
OAI21X1 OAI21X1_118 ( .A(_359_), .B(_356_), .C(_361_), .Y(_20__2_) );
INVX1 INVX1_60 ( .A(_20__2_), .Y(_366_) );
OR2X2 OR2X2_86 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_367_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_368_) );
NAND3X1 NAND3X1_60 ( .A(_366_), .B(_368_), .C(_367_), .Y(_369_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_363_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_364_) );
OAI21X1 OAI21X1_119 ( .A(_363_), .B(_364_), .C(_20__2_), .Y(_365_) );
NAND2X1 NAND2X1_94 ( .A(_365_), .B(_369_), .Y(_0__42_) );
OAI21X1 OAI21X1_120 ( .A(_366_), .B(_363_), .C(_368_), .Y(_20__3_) );
INVX1 INVX1_61 ( .A(_20__3_), .Y(_373_) );
OR2X2 OR2X2_87 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_374_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_375_) );
NAND3X1 NAND3X1_61 ( .A(_373_), .B(_375_), .C(_374_), .Y(_376_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_370_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_371_) );
OAI21X1 OAI21X1_121 ( .A(_370_), .B(_371_), .C(_20__3_), .Y(_372_) );
NAND2X1 NAND2X1_96 ( .A(_372_), .B(_376_), .Y(_0__43_) );
OAI21X1 OAI21X1_122 ( .A(_373_), .B(_370_), .C(_375_), .Y(_19_) );
INVX1 INVX1_62 ( .A(w_cout_10_), .Y(_380_) );
OR2X2 OR2X2_88 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_381_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_382_) );
NAND3X1 NAND3X1_62 ( .A(_380_), .B(_382_), .C(_381_), .Y(_383_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_377_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_378_) );
OAI21X1 OAI21X1_123 ( .A(_377_), .B(_378_), .C(w_cout_10_), .Y(_379_) );
NAND2X1 NAND2X1_98 ( .A(_379_), .B(_383_), .Y(_0__44_) );
OAI21X1 OAI21X1_124 ( .A(_380_), .B(_377_), .C(_382_), .Y(_22__1_) );
INVX1 INVX1_63 ( .A(_22__1_), .Y(_387_) );
OR2X2 OR2X2_89 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_388_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_389_) );
NAND3X1 NAND3X1_63 ( .A(_387_), .B(_389_), .C(_388_), .Y(_390_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_384_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_385_) );
OAI21X1 OAI21X1_125 ( .A(_384_), .B(_385_), .C(_22__1_), .Y(_386_) );
NAND2X1 NAND2X1_100 ( .A(_386_), .B(_390_), .Y(_0__45_) );
OAI21X1 OAI21X1_126 ( .A(_387_), .B(_384_), .C(_389_), .Y(_22__2_) );
INVX1 INVX1_64 ( .A(_22__2_), .Y(_394_) );
OR2X2 OR2X2_90 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_395_) );
NAND2X1 NAND2X1_101 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_396_) );
NAND3X1 NAND3X1_64 ( .A(_394_), .B(_396_), .C(_395_), .Y(_397_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_391_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_392_) );
OAI21X1 OAI21X1_127 ( .A(_391_), .B(_392_), .C(_22__2_), .Y(_393_) );
NAND2X1 NAND2X1_102 ( .A(_393_), .B(_397_), .Y(_0__46_) );
OAI21X1 OAI21X1_128 ( .A(_394_), .B(_391_), .C(_396_), .Y(_22__3_) );
INVX1 INVX1_65 ( .A(_22__3_), .Y(_401_) );
OR2X2 OR2X2_91 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_402_) );
NAND2X1 NAND2X1_103 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_403_) );
NAND3X1 NAND3X1_65 ( .A(_401_), .B(_403_), .C(_402_), .Y(_404_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_398_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_399_) );
OAI21X1 OAI21X1_129 ( .A(_398_), .B(_399_), .C(_22__3_), .Y(_400_) );
NAND2X1 NAND2X1_104 ( .A(_400_), .B(_404_), .Y(_0__47_) );
OAI21X1 OAI21X1_130 ( .A(_401_), .B(_398_), .C(_403_), .Y(_21_) );
BUFX2 BUFX2_54 ( .A(skip0_cin_next), .Y(_2__0_) );
BUFX2 BUFX2_55 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_56 ( .A(w_cout_1_), .Y(_4__0_) );
BUFX2 BUFX2_57 ( .A(_3_), .Y(_4__4_) );
BUFX2 BUFX2_58 ( .A(w_cout_2_), .Y(_6__0_) );
BUFX2 BUFX2_59 ( .A(_5_), .Y(_6__4_) );
BUFX2 BUFX2_60 ( .A(w_cout_3_), .Y(_8__0_) );
BUFX2 BUFX2_61 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_62 ( .A(w_cout_4_), .Y(_10__0_) );
BUFX2 BUFX2_63 ( .A(_9_), .Y(_10__4_) );
BUFX2 BUFX2_64 ( .A(w_cout_5_), .Y(_12__0_) );
BUFX2 BUFX2_65 ( .A(_11_), .Y(_12__4_) );
BUFX2 BUFX2_66 ( .A(w_cout_6_), .Y(_14__0_) );
BUFX2 BUFX2_67 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_68 ( .A(w_cout_7_), .Y(_16__0_) );
BUFX2 BUFX2_69 ( .A(_15_), .Y(_16__4_) );
BUFX2 BUFX2_70 ( .A(w_cout_8_), .Y(_18__0_) );
BUFX2 BUFX2_71 ( .A(_17_), .Y(_18__4_) );
BUFX2 BUFX2_72 ( .A(w_cout_9_), .Y(_20__0_) );
BUFX2 BUFX2_73 ( .A(_19_), .Y(_20__4_) );
BUFX2 BUFX2_74 ( .A(w_cout_10_), .Y(_22__0_) );
BUFX2 BUFX2_75 ( .A(_21_), .Y(_22__4_) );
BUFX2 BUFX2_76 ( .A(w_cout_11_), .Y(_24__0_) );
BUFX2 BUFX2_77 ( .A(_23_), .Y(_24__4_) );
BUFX2 BUFX2_78 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_79 ( .A(cout0), .Y(rca_inst_w_CARRY_4_) );
BUFX2 BUFX2_80 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
