module CSkipA_53bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [52:0] i_add_term1;
input [52:0] i_add_term2;
output [52:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

OAI21X1 OAI21X1_1 ( .A(_307_), .B(_304_), .C(_309_), .Y(_8__1_) );
INVX1 INVX1_1 ( .A(_8__1_), .Y(_314_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_315_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_316_) );
NAND3X1 NAND3X1_1 ( .A(_314_), .B(_316_), .C(_315_), .Y(_317_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_311_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_312_) );
OAI21X1 OAI21X1_2 ( .A(_311_), .B(_312_), .C(_8__1_), .Y(_313_) );
NAND2X1 NAND2X1_2 ( .A(_313_), .B(_317_), .Y(_0__9_) );
OAI21X1 OAI21X1_3 ( .A(_314_), .B(_311_), .C(_316_), .Y(_8__2_) );
INVX1 INVX1_2 ( .A(_8__2_), .Y(_321_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_322_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_323_) );
NAND3X1 NAND3X1_2 ( .A(_321_), .B(_323_), .C(_322_), .Y(_324_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_318_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_319_) );
OAI21X1 OAI21X1_4 ( .A(_318_), .B(_319_), .C(_8__2_), .Y(_320_) );
NAND2X1 NAND2X1_4 ( .A(_320_), .B(_324_), .Y(_0__10_) );
OAI21X1 OAI21X1_5 ( .A(_321_), .B(_318_), .C(_323_), .Y(_8__3_) );
INVX1 INVX1_3 ( .A(_8__3_), .Y(_328_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_329_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_330_) );
NAND3X1 NAND3X1_3 ( .A(_328_), .B(_330_), .C(_329_), .Y(_331_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_325_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_326_) );
OAI21X1 OAI21X1_6 ( .A(_325_), .B(_326_), .C(_8__3_), .Y(_327_) );
NAND2X1 NAND2X1_6 ( .A(_327_), .B(_331_), .Y(_0__11_) );
OAI21X1 OAI21X1_7 ( .A(_328_), .B(_325_), .C(_330_), .Y(_7_) );
INVX1 INVX1_4 ( .A(w_cout_3_), .Y(_335_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_336_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_337_) );
NAND3X1 NAND3X1_4 ( .A(_335_), .B(_337_), .C(_336_), .Y(_338_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_332_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_333_) );
OAI21X1 OAI21X1_8 ( .A(_332_), .B(_333_), .C(w_cout_3_), .Y(_334_) );
NAND2X1 NAND2X1_8 ( .A(_334_), .B(_338_), .Y(_0__12_) );
OAI21X1 OAI21X1_9 ( .A(_335_), .B(_332_), .C(_337_), .Y(_11__1_) );
INVX1 INVX1_5 ( .A(_11__1_), .Y(_342_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_343_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_344_) );
NAND3X1 NAND3X1_5 ( .A(_342_), .B(_344_), .C(_343_), .Y(_345_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_339_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_340_) );
OAI21X1 OAI21X1_10 ( .A(_339_), .B(_340_), .C(_11__1_), .Y(_341_) );
NAND2X1 NAND2X1_10 ( .A(_341_), .B(_345_), .Y(_0__13_) );
OAI21X1 OAI21X1_11 ( .A(_342_), .B(_339_), .C(_344_), .Y(_11__2_) );
INVX1 INVX1_6 ( .A(_11__2_), .Y(_349_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_350_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_351_) );
NAND3X1 NAND3X1_6 ( .A(_349_), .B(_351_), .C(_350_), .Y(_352_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_346_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_347_) );
OAI21X1 OAI21X1_12 ( .A(_346_), .B(_347_), .C(_11__2_), .Y(_348_) );
NAND2X1 NAND2X1_12 ( .A(_348_), .B(_352_), .Y(_0__14_) );
OAI21X1 OAI21X1_13 ( .A(_349_), .B(_346_), .C(_351_), .Y(_11__3_) );
INVX1 INVX1_7 ( .A(_11__3_), .Y(_356_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_357_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_358_) );
NAND3X1 NAND3X1_7 ( .A(_356_), .B(_358_), .C(_357_), .Y(_359_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_353_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_354_) );
OAI21X1 OAI21X1_14 ( .A(_353_), .B(_354_), .C(_11__3_), .Y(_355_) );
NAND2X1 NAND2X1_14 ( .A(_355_), .B(_359_), .Y(_0__15_) );
OAI21X1 OAI21X1_15 ( .A(_356_), .B(_353_), .C(_358_), .Y(_10_) );
INVX1 INVX1_8 ( .A(w_cout_4_), .Y(_363_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_364_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_365_) );
NAND3X1 NAND3X1_8 ( .A(_363_), .B(_365_), .C(_364_), .Y(_366_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_360_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_361_) );
OAI21X1 OAI21X1_16 ( .A(_360_), .B(_361_), .C(w_cout_4_), .Y(_362_) );
NAND2X1 NAND2X1_16 ( .A(_362_), .B(_366_), .Y(_0__16_) );
OAI21X1 OAI21X1_17 ( .A(_363_), .B(_360_), .C(_365_), .Y(_14__1_) );
INVX1 INVX1_9 ( .A(_14__1_), .Y(_370_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_371_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_372_) );
NAND3X1 NAND3X1_9 ( .A(_370_), .B(_372_), .C(_371_), .Y(_373_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_367_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_368_) );
OAI21X1 OAI21X1_18 ( .A(_367_), .B(_368_), .C(_14__1_), .Y(_369_) );
NAND2X1 NAND2X1_18 ( .A(_369_), .B(_373_), .Y(_0__17_) );
OAI21X1 OAI21X1_19 ( .A(_370_), .B(_367_), .C(_372_), .Y(_14__2_) );
INVX1 INVX1_10 ( .A(_14__2_), .Y(_377_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_378_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_379_) );
NAND3X1 NAND3X1_10 ( .A(_377_), .B(_379_), .C(_378_), .Y(_380_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_374_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_375_) );
OAI21X1 OAI21X1_20 ( .A(_374_), .B(_375_), .C(_14__2_), .Y(_376_) );
NAND2X1 NAND2X1_20 ( .A(_376_), .B(_380_), .Y(_0__18_) );
OAI21X1 OAI21X1_21 ( .A(_377_), .B(_374_), .C(_379_), .Y(_14__3_) );
INVX1 INVX1_11 ( .A(_14__3_), .Y(_384_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_385_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_386_) );
NAND3X1 NAND3X1_11 ( .A(_384_), .B(_386_), .C(_385_), .Y(_387_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_381_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_382_) );
OAI21X1 OAI21X1_22 ( .A(_381_), .B(_382_), .C(_14__3_), .Y(_383_) );
NAND2X1 NAND2X1_22 ( .A(_383_), .B(_387_), .Y(_0__19_) );
OAI21X1 OAI21X1_23 ( .A(_384_), .B(_381_), .C(_386_), .Y(_13_) );
INVX1 INVX1_12 ( .A(w_cout_5_), .Y(_391_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_392_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_393_) );
NAND3X1 NAND3X1_12 ( .A(_391_), .B(_393_), .C(_392_), .Y(_394_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_388_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_389_) );
OAI21X1 OAI21X1_24 ( .A(_388_), .B(_389_), .C(w_cout_5_), .Y(_390_) );
NAND2X1 NAND2X1_24 ( .A(_390_), .B(_394_), .Y(_0__20_) );
OAI21X1 OAI21X1_25 ( .A(_391_), .B(_388_), .C(_393_), .Y(_17__1_) );
INVX1 INVX1_13 ( .A(_17__1_), .Y(_398_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_399_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_400_) );
NAND3X1 NAND3X1_13 ( .A(_398_), .B(_400_), .C(_399_), .Y(_401_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_395_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_396_) );
OAI21X1 OAI21X1_26 ( .A(_395_), .B(_396_), .C(_17__1_), .Y(_397_) );
NAND2X1 NAND2X1_26 ( .A(_397_), .B(_401_), .Y(_0__21_) );
OAI21X1 OAI21X1_27 ( .A(_398_), .B(_395_), .C(_400_), .Y(_17__2_) );
INVX1 INVX1_14 ( .A(_17__2_), .Y(_405_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_406_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_407_) );
NAND3X1 NAND3X1_14 ( .A(_405_), .B(_407_), .C(_406_), .Y(_408_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_402_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_403_) );
OAI21X1 OAI21X1_28 ( .A(_402_), .B(_403_), .C(_17__2_), .Y(_404_) );
NAND2X1 NAND2X1_28 ( .A(_404_), .B(_408_), .Y(_0__22_) );
OAI21X1 OAI21X1_29 ( .A(_405_), .B(_402_), .C(_407_), .Y(_17__3_) );
INVX1 INVX1_15 ( .A(_17__3_), .Y(_412_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_413_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_414_) );
NAND3X1 NAND3X1_15 ( .A(_412_), .B(_414_), .C(_413_), .Y(_415_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_409_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_410_) );
OAI21X1 OAI21X1_30 ( .A(_409_), .B(_410_), .C(_17__3_), .Y(_411_) );
NAND2X1 NAND2X1_30 ( .A(_411_), .B(_415_), .Y(_0__23_) );
OAI21X1 OAI21X1_31 ( .A(_412_), .B(_409_), .C(_414_), .Y(_16_) );
INVX1 INVX1_16 ( .A(w_cout_6_), .Y(_419_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_420_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_421_) );
NAND3X1 NAND3X1_16 ( .A(_419_), .B(_421_), .C(_420_), .Y(_422_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_416_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_417_) );
OAI21X1 OAI21X1_32 ( .A(_416_), .B(_417_), .C(w_cout_6_), .Y(_418_) );
NAND2X1 NAND2X1_32 ( .A(_418_), .B(_422_), .Y(_0__24_) );
OAI21X1 OAI21X1_33 ( .A(_419_), .B(_416_), .C(_421_), .Y(_20__1_) );
INVX1 INVX1_17 ( .A(_20__1_), .Y(_426_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_427_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_428_) );
NAND3X1 NAND3X1_17 ( .A(_426_), .B(_428_), .C(_427_), .Y(_429_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_423_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_424_) );
OAI21X1 OAI21X1_34 ( .A(_423_), .B(_424_), .C(_20__1_), .Y(_425_) );
NAND2X1 NAND2X1_34 ( .A(_425_), .B(_429_), .Y(_0__25_) );
OAI21X1 OAI21X1_35 ( .A(_426_), .B(_423_), .C(_428_), .Y(_20__2_) );
INVX1 INVX1_18 ( .A(_20__2_), .Y(_433_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_434_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_435_) );
NAND3X1 NAND3X1_18 ( .A(_433_), .B(_435_), .C(_434_), .Y(_436_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_430_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_431_) );
OAI21X1 OAI21X1_36 ( .A(_430_), .B(_431_), .C(_20__2_), .Y(_432_) );
NAND2X1 NAND2X1_36 ( .A(_432_), .B(_436_), .Y(_0__26_) );
OAI21X1 OAI21X1_37 ( .A(_433_), .B(_430_), .C(_435_), .Y(_20__3_) );
INVX1 INVX1_19 ( .A(_20__3_), .Y(_440_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_441_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_442_) );
NAND3X1 NAND3X1_19 ( .A(_440_), .B(_442_), .C(_441_), .Y(_443_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_437_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_438_) );
OAI21X1 OAI21X1_38 ( .A(_437_), .B(_438_), .C(_20__3_), .Y(_439_) );
NAND2X1 NAND2X1_38 ( .A(_439_), .B(_443_), .Y(_0__27_) );
OAI21X1 OAI21X1_39 ( .A(_440_), .B(_437_), .C(_442_), .Y(_19_) );
INVX1 INVX1_20 ( .A(w_cout_7_), .Y(_447_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_448_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_449_) );
NAND3X1 NAND3X1_20 ( .A(_447_), .B(_449_), .C(_448_), .Y(_450_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_444_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_445_) );
OAI21X1 OAI21X1_40 ( .A(_444_), .B(_445_), .C(w_cout_7_), .Y(_446_) );
NAND2X1 NAND2X1_40 ( .A(_446_), .B(_450_), .Y(_0__28_) );
OAI21X1 OAI21X1_41 ( .A(_447_), .B(_444_), .C(_449_), .Y(_23__1_) );
INVX1 INVX1_21 ( .A(_23__1_), .Y(_454_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_455_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_456_) );
NAND3X1 NAND3X1_21 ( .A(_454_), .B(_456_), .C(_455_), .Y(_457_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_451_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_452_) );
OAI21X1 OAI21X1_42 ( .A(_451_), .B(_452_), .C(_23__1_), .Y(_453_) );
NAND2X1 NAND2X1_42 ( .A(_453_), .B(_457_), .Y(_0__29_) );
OAI21X1 OAI21X1_43 ( .A(_454_), .B(_451_), .C(_456_), .Y(_23__2_) );
INVX1 INVX1_22 ( .A(_23__2_), .Y(_461_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_462_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_463_) );
NAND3X1 NAND3X1_22 ( .A(_461_), .B(_463_), .C(_462_), .Y(_464_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_458_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_459_) );
OAI21X1 OAI21X1_44 ( .A(_458_), .B(_459_), .C(_23__2_), .Y(_460_) );
NAND2X1 NAND2X1_44 ( .A(_460_), .B(_464_), .Y(_0__30_) );
OAI21X1 OAI21X1_45 ( .A(_461_), .B(_458_), .C(_463_), .Y(_23__3_) );
INVX1 INVX1_23 ( .A(_23__3_), .Y(_468_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_469_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_470_) );
NAND3X1 NAND3X1_23 ( .A(_468_), .B(_470_), .C(_469_), .Y(_471_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_465_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_466_) );
OAI21X1 OAI21X1_46 ( .A(_465_), .B(_466_), .C(_23__3_), .Y(_467_) );
NAND2X1 NAND2X1_46 ( .A(_467_), .B(_471_), .Y(_0__31_) );
OAI21X1 OAI21X1_47 ( .A(_468_), .B(_465_), .C(_470_), .Y(_22_) );
INVX1 INVX1_24 ( .A(w_cout_8_), .Y(_475_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_476_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_477_) );
NAND3X1 NAND3X1_24 ( .A(_475_), .B(_477_), .C(_476_), .Y(_478_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_472_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_473_) );
OAI21X1 OAI21X1_48 ( .A(_472_), .B(_473_), .C(w_cout_8_), .Y(_474_) );
NAND2X1 NAND2X1_48 ( .A(_474_), .B(_478_), .Y(_0__32_) );
OAI21X1 OAI21X1_49 ( .A(_475_), .B(_472_), .C(_477_), .Y(_26__1_) );
INVX1 INVX1_25 ( .A(_26__1_), .Y(_482_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_483_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_484_) );
NAND3X1 NAND3X1_25 ( .A(_482_), .B(_484_), .C(_483_), .Y(_485_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_479_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_480_) );
OAI21X1 OAI21X1_50 ( .A(_479_), .B(_480_), .C(_26__1_), .Y(_481_) );
NAND2X1 NAND2X1_50 ( .A(_481_), .B(_485_), .Y(_0__33_) );
OAI21X1 OAI21X1_51 ( .A(_482_), .B(_479_), .C(_484_), .Y(_26__2_) );
INVX1 INVX1_26 ( .A(_26__2_), .Y(_489_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_490_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_491_) );
NAND3X1 NAND3X1_26 ( .A(_489_), .B(_491_), .C(_490_), .Y(_492_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_486_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_487_) );
OAI21X1 OAI21X1_52 ( .A(_486_), .B(_487_), .C(_26__2_), .Y(_488_) );
NAND2X1 NAND2X1_52 ( .A(_488_), .B(_492_), .Y(_0__34_) );
OAI21X1 OAI21X1_53 ( .A(_489_), .B(_486_), .C(_491_), .Y(_26__3_) );
INVX1 INVX1_27 ( .A(_26__3_), .Y(_496_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_497_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_498_) );
NAND3X1 NAND3X1_27 ( .A(_496_), .B(_498_), .C(_497_), .Y(_499_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_493_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_494_) );
OAI21X1 OAI21X1_54 ( .A(_493_), .B(_494_), .C(_26__3_), .Y(_495_) );
NAND2X1 NAND2X1_54 ( .A(_495_), .B(_499_), .Y(_0__35_) );
OAI21X1 OAI21X1_55 ( .A(_496_), .B(_493_), .C(_498_), .Y(_25_) );
INVX1 INVX1_28 ( .A(w_cout_9_), .Y(_503_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_504_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_505_) );
NAND3X1 NAND3X1_28 ( .A(_503_), .B(_505_), .C(_504_), .Y(_506_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_500_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_501_) );
OAI21X1 OAI21X1_56 ( .A(_500_), .B(_501_), .C(w_cout_9_), .Y(_502_) );
NAND2X1 NAND2X1_56 ( .A(_502_), .B(_506_), .Y(_0__36_) );
OAI21X1 OAI21X1_57 ( .A(_503_), .B(_500_), .C(_505_), .Y(_29__1_) );
INVX1 INVX1_29 ( .A(_29__1_), .Y(_510_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_511_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_512_) );
NAND3X1 NAND3X1_29 ( .A(_510_), .B(_512_), .C(_511_), .Y(_513_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_507_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_508_) );
OAI21X1 OAI21X1_58 ( .A(_507_), .B(_508_), .C(_29__1_), .Y(_509_) );
NAND2X1 NAND2X1_58 ( .A(_509_), .B(_513_), .Y(_0__37_) );
OAI21X1 OAI21X1_59 ( .A(_510_), .B(_507_), .C(_512_), .Y(_29__2_) );
INVX1 INVX1_30 ( .A(_29__2_), .Y(_517_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_518_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_519_) );
NAND3X1 NAND3X1_30 ( .A(_517_), .B(_519_), .C(_518_), .Y(_520_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_514_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_515_) );
OAI21X1 OAI21X1_60 ( .A(_514_), .B(_515_), .C(_29__2_), .Y(_516_) );
NAND2X1 NAND2X1_60 ( .A(_516_), .B(_520_), .Y(_0__38_) );
OAI21X1 OAI21X1_61 ( .A(_517_), .B(_514_), .C(_519_), .Y(_29__3_) );
INVX1 INVX1_31 ( .A(_29__3_), .Y(_524_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_525_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_526_) );
NAND3X1 NAND3X1_31 ( .A(_524_), .B(_526_), .C(_525_), .Y(_527_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_521_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_522_) );
OAI21X1 OAI21X1_62 ( .A(_521_), .B(_522_), .C(_29__3_), .Y(_523_) );
NAND2X1 NAND2X1_62 ( .A(_523_), .B(_527_), .Y(_0__39_) );
OAI21X1 OAI21X1_63 ( .A(_524_), .B(_521_), .C(_526_), .Y(_28_) );
INVX1 INVX1_32 ( .A(w_cout_10_), .Y(_531_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_532_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_533_) );
NAND3X1 NAND3X1_32 ( .A(_531_), .B(_533_), .C(_532_), .Y(_534_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_528_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_529_) );
OAI21X1 OAI21X1_64 ( .A(_528_), .B(_529_), .C(w_cout_10_), .Y(_530_) );
NAND2X1 NAND2X1_64 ( .A(_530_), .B(_534_), .Y(_0__40_) );
OAI21X1 OAI21X1_65 ( .A(_531_), .B(_528_), .C(_533_), .Y(_32__1_) );
INVX1 INVX1_33 ( .A(_32__1_), .Y(_538_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_539_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_540_) );
NAND3X1 NAND3X1_33 ( .A(_538_), .B(_540_), .C(_539_), .Y(_541_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_535_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_536_) );
OAI21X1 OAI21X1_66 ( .A(_535_), .B(_536_), .C(_32__1_), .Y(_537_) );
NAND2X1 NAND2X1_66 ( .A(_537_), .B(_541_), .Y(_0__41_) );
OAI21X1 OAI21X1_67 ( .A(_538_), .B(_535_), .C(_540_), .Y(_32__2_) );
INVX1 INVX1_34 ( .A(_32__2_), .Y(_545_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_546_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_547_) );
NAND3X1 NAND3X1_34 ( .A(_545_), .B(_547_), .C(_546_), .Y(_548_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_542_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_543_) );
OAI21X1 OAI21X1_68 ( .A(_542_), .B(_543_), .C(_32__2_), .Y(_544_) );
NAND2X1 NAND2X1_68 ( .A(_544_), .B(_548_), .Y(_0__42_) );
OAI21X1 OAI21X1_69 ( .A(_545_), .B(_542_), .C(_547_), .Y(_32__3_) );
INVX1 INVX1_35 ( .A(_32__3_), .Y(_552_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_553_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_554_) );
NAND3X1 NAND3X1_35 ( .A(_552_), .B(_554_), .C(_553_), .Y(_555_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_549_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_550_) );
OAI21X1 OAI21X1_70 ( .A(_549_), .B(_550_), .C(_32__3_), .Y(_551_) );
NAND2X1 NAND2X1_70 ( .A(_551_), .B(_555_), .Y(_0__43_) );
OAI21X1 OAI21X1_71 ( .A(_552_), .B(_549_), .C(_554_), .Y(_31_) );
INVX1 INVX1_36 ( .A(w_cout_11_), .Y(_559_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_560_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_561_) );
NAND3X1 NAND3X1_36 ( .A(_559_), .B(_561_), .C(_560_), .Y(_562_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_556_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_557_) );
OAI21X1 OAI21X1_72 ( .A(_556_), .B(_557_), .C(w_cout_11_), .Y(_558_) );
NAND2X1 NAND2X1_72 ( .A(_558_), .B(_562_), .Y(_0__44_) );
OAI21X1 OAI21X1_73 ( .A(_559_), .B(_556_), .C(_561_), .Y(_35__1_) );
INVX1 INVX1_37 ( .A(_35__1_), .Y(_566_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_567_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_568_) );
NAND3X1 NAND3X1_37 ( .A(_566_), .B(_568_), .C(_567_), .Y(_569_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_563_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_564_) );
OAI21X1 OAI21X1_74 ( .A(_563_), .B(_564_), .C(_35__1_), .Y(_565_) );
NAND2X1 NAND2X1_74 ( .A(_565_), .B(_569_), .Y(_0__45_) );
OAI21X1 OAI21X1_75 ( .A(_566_), .B(_563_), .C(_568_), .Y(_35__2_) );
INVX1 INVX1_38 ( .A(_35__2_), .Y(_573_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_574_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_575_) );
NAND3X1 NAND3X1_38 ( .A(_573_), .B(_575_), .C(_574_), .Y(_576_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_570_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_571_) );
OAI21X1 OAI21X1_76 ( .A(_570_), .B(_571_), .C(_35__2_), .Y(_572_) );
NAND2X1 NAND2X1_76 ( .A(_572_), .B(_576_), .Y(_0__46_) );
OAI21X1 OAI21X1_77 ( .A(_573_), .B(_570_), .C(_575_), .Y(_35__3_) );
INVX1 INVX1_39 ( .A(_35__3_), .Y(_580_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_581_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_582_) );
NAND3X1 NAND3X1_39 ( .A(_580_), .B(_582_), .C(_581_), .Y(_583_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_577_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_578_) );
OAI21X1 OAI21X1_78 ( .A(_577_), .B(_578_), .C(_35__3_), .Y(_579_) );
NAND2X1 NAND2X1_78 ( .A(_579_), .B(_583_), .Y(_0__47_) );
OAI21X1 OAI21X1_79 ( .A(_580_), .B(_577_), .C(_582_), .Y(_34_) );
INVX1 INVX1_40 ( .A(w_cout_12_), .Y(_587_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_588_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_589_) );
NAND3X1 NAND3X1_40 ( .A(_587_), .B(_589_), .C(_588_), .Y(_590_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_584_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_585_) );
OAI21X1 OAI21X1_80 ( .A(_584_), .B(_585_), .C(w_cout_12_), .Y(_586_) );
NAND2X1 NAND2X1_80 ( .A(_586_), .B(_590_), .Y(_0__48_) );
OAI21X1 OAI21X1_81 ( .A(_587_), .B(_584_), .C(_589_), .Y(_38__1_) );
INVX1 INVX1_41 ( .A(_38__1_), .Y(_594_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_595_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_596_) );
NAND3X1 NAND3X1_41 ( .A(_594_), .B(_596_), .C(_595_), .Y(_597_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_591_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_592_) );
OAI21X1 OAI21X1_82 ( .A(_591_), .B(_592_), .C(_38__1_), .Y(_593_) );
NAND2X1 NAND2X1_82 ( .A(_593_), .B(_597_), .Y(_0__49_) );
OAI21X1 OAI21X1_83 ( .A(_594_), .B(_591_), .C(_596_), .Y(_38__2_) );
INVX1 INVX1_42 ( .A(_38__2_), .Y(_601_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_602_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_603_) );
NAND3X1 NAND3X1_42 ( .A(_601_), .B(_603_), .C(_602_), .Y(_604_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_598_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_599_) );
OAI21X1 OAI21X1_84 ( .A(_598_), .B(_599_), .C(_38__2_), .Y(_600_) );
NAND2X1 NAND2X1_84 ( .A(_600_), .B(_604_), .Y(_0__50_) );
OAI21X1 OAI21X1_85 ( .A(_601_), .B(_598_), .C(_603_), .Y(_38__3_) );
INVX1 INVX1_43 ( .A(_38__3_), .Y(_608_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_609_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_610_) );
NAND3X1 NAND3X1_43 ( .A(_608_), .B(_610_), .C(_609_), .Y(_611_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_605_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_606_) );
OAI21X1 OAI21X1_86 ( .A(_605_), .B(_606_), .C(_38__3_), .Y(_607_) );
NAND2X1 NAND2X1_86 ( .A(_607_), .B(_611_), .Y(_0__51_) );
OAI21X1 OAI21X1_87 ( .A(_608_), .B(_605_), .C(_610_), .Y(_37_) );
INVX1 INVX1_44 ( .A(cskip1_inst_cin), .Y(_615_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_616_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_617_) );
NAND3X1 NAND3X1_44 ( .A(_615_), .B(_617_), .C(_616_), .Y(_618_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_612_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_613_) );
OAI21X1 OAI21X1_88 ( .A(_612_), .B(_613_), .C(cskip1_inst_cin), .Y(_614_) );
NAND2X1 NAND2X1_88 ( .A(_614_), .B(_618_), .Y(cskip1_inst_sum) );
OAI21X1 OAI21X1_89 ( .A(_615_), .B(_612_), .C(_617_), .Y(cskip1_inst_rca0_w_CARRY_1_) );
INVX1 INVX1_45 ( .A(cskip1_inst_rca0_w_CARRY_1_), .Y(_620_) );
NAND2X1 NAND2X1_89 ( .A(gnd), .B(gnd), .Y(_621_) );
NOR2X1 NOR2X1_45 ( .A(gnd), .B(gnd), .Y(_619_) );
OAI21X1 OAI21X1_90 ( .A(_620_), .B(_619_), .C(_621_), .Y(cskip1_inst_rca0_w_CARRY_2_) );
INVX1 INVX1_46 ( .A(cskip1_inst_rca0_w_CARRY_2_), .Y(_623_) );
NAND2X1 NAND2X1_90 ( .A(gnd), .B(gnd), .Y(_624_) );
NOR2X1 NOR2X1_46 ( .A(gnd), .B(gnd), .Y(_622_) );
OAI21X1 OAI21X1_91 ( .A(_623_), .B(_622_), .C(_624_), .Y(cskip1_inst_rca0_w_CARRY_3_) );
INVX1 INVX1_47 ( .A(cskip1_inst_rca0_w_CARRY_3_), .Y(_626_) );
NAND2X1 NAND2X1_91 ( .A(gnd), .B(gnd), .Y(_627_) );
NOR2X1 NOR2X1_47 ( .A(gnd), .B(gnd), .Y(_625_) );
OAI21X1 OAI21X1_92 ( .A(_626_), .B(_625_), .C(_627_), .Y(cskip1_inst_cout0) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_628_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_629_) );
NOR2X1 NOR2X1_49 ( .A(_628_), .B(_629_), .Y(cskip1_inst_skip0_P) );
INVX1 INVX1_48 ( .A(cskip1_inst_cout0), .Y(_630_) );
NAND2X1 NAND2X1_92 ( .A(gnd), .B(cskip1_inst_skip0_P), .Y(_631_) );
OAI21X1 OAI21X1_93 ( .A(cskip1_inst_skip0_P), .B(_630_), .C(_631_), .Y(w_cout_14_) );
BUFX2 BUFX2_1 ( .A(w_cout_14_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .A(cskip1_inst_sum), .Y(sum[52]) );
INVX1 INVX1_49 ( .A(i_add_term1[0]), .Y(_40_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[0]), .B(_40_), .Y(_41_) );
INVX1 INVX1_50 ( .A(i_add_term2[0]), .Y(_42_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term1[0]), .B(_42_), .Y(_43_) );
INVX1 INVX1_51 ( .A(i_add_term1[1]), .Y(_44_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[1]), .B(_44_), .Y(_45_) );
INVX1 INVX1_52 ( .A(i_add_term2[1]), .Y(_46_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term1[1]), .B(_46_), .Y(_47_) );
OAI22X1 OAI22X1_1 ( .A(_41_), .B(_43_), .C(_45_), .D(_47_), .Y(_48_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_49_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_50_) );
NOR2X1 NOR2X1_55 ( .A(_49_), .B(_50_), .Y(_51_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_52_) );
NAND2X1 NAND2X1_93 ( .A(_51_), .B(_52_), .Y(_53_) );
NOR2X1 NOR2X1_56 ( .A(_48_), .B(_53_), .Y(_3_) );
INVX1 INVX1_53 ( .A(_1_), .Y(_54_) );
NAND2X1 NAND2X1_94 ( .A(gnd), .B(_3_), .Y(_55_) );
OAI21X1 OAI21X1_94 ( .A(_3_), .B(_54_), .C(_55_), .Y(w_cout_1_) );
INVX1 INVX1_54 ( .A(i_add_term1[4]), .Y(_56_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[4]), .B(_56_), .Y(_57_) );
INVX1 INVX1_55 ( .A(i_add_term2[4]), .Y(_58_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term1[4]), .B(_58_), .Y(_59_) );
INVX1 INVX1_56 ( .A(i_add_term1[5]), .Y(_60_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[5]), .B(_60_), .Y(_61_) );
INVX1 INVX1_57 ( .A(i_add_term2[5]), .Y(_62_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term1[5]), .B(_62_), .Y(_63_) );
OAI22X1 OAI22X1_2 ( .A(_57_), .B(_59_), .C(_61_), .D(_63_), .Y(_64_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_65_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_66_) );
NOR2X1 NOR2X1_62 ( .A(_65_), .B(_66_), .Y(_67_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_68_) );
NAND2X1 NAND2X1_95 ( .A(_67_), .B(_68_), .Y(_69_) );
NOR2X1 NOR2X1_63 ( .A(_64_), .B(_69_), .Y(_6_) );
INVX1 INVX1_58 ( .A(_4_), .Y(_70_) );
NAND2X1 NAND2X1_96 ( .A(gnd), .B(_6_), .Y(_71_) );
OAI21X1 OAI21X1_95 ( .A(_6_), .B(_70_), .C(_71_), .Y(w_cout_2_) );
INVX1 INVX1_59 ( .A(i_add_term1[8]), .Y(_72_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[8]), .B(_72_), .Y(_73_) );
INVX1 INVX1_60 ( .A(i_add_term2[8]), .Y(_74_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term1[8]), .B(_74_), .Y(_75_) );
INVX1 INVX1_61 ( .A(i_add_term1[9]), .Y(_76_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[9]), .B(_76_), .Y(_77_) );
INVX1 INVX1_62 ( .A(i_add_term2[9]), .Y(_78_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term1[9]), .B(_78_), .Y(_79_) );
OAI22X1 OAI22X1_3 ( .A(_73_), .B(_75_), .C(_77_), .D(_79_), .Y(_80_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_81_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_82_) );
NOR2X1 NOR2X1_69 ( .A(_81_), .B(_82_), .Y(_83_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_84_) );
NAND2X1 NAND2X1_97 ( .A(_83_), .B(_84_), .Y(_85_) );
NOR2X1 NOR2X1_70 ( .A(_80_), .B(_85_), .Y(_9_) );
INVX1 INVX1_63 ( .A(_7_), .Y(_86_) );
NAND2X1 NAND2X1_98 ( .A(gnd), .B(_9_), .Y(_87_) );
OAI21X1 OAI21X1_96 ( .A(_9_), .B(_86_), .C(_87_), .Y(w_cout_3_) );
INVX1 INVX1_64 ( .A(i_add_term1[12]), .Y(_88_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[12]), .B(_88_), .Y(_89_) );
INVX1 INVX1_65 ( .A(i_add_term2[12]), .Y(_90_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term1[12]), .B(_90_), .Y(_91_) );
INVX1 INVX1_66 ( .A(i_add_term1[13]), .Y(_92_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[13]), .B(_92_), .Y(_93_) );
INVX1 INVX1_67 ( .A(i_add_term2[13]), .Y(_94_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term1[13]), .B(_94_), .Y(_95_) );
OAI22X1 OAI22X1_4 ( .A(_89_), .B(_91_), .C(_93_), .D(_95_), .Y(_96_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_97_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_98_) );
NOR2X1 NOR2X1_76 ( .A(_97_), .B(_98_), .Y(_99_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_100_) );
NAND2X1 NAND2X1_99 ( .A(_99_), .B(_100_), .Y(_101_) );
NOR2X1 NOR2X1_77 ( .A(_96_), .B(_101_), .Y(_12_) );
INVX1 INVX1_68 ( .A(_10_), .Y(_102_) );
NAND2X1 NAND2X1_100 ( .A(gnd), .B(_12_), .Y(_103_) );
OAI21X1 OAI21X1_97 ( .A(_12_), .B(_102_), .C(_103_), .Y(w_cout_4_) );
INVX1 INVX1_69 ( .A(i_add_term1[16]), .Y(_104_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[16]), .B(_104_), .Y(_105_) );
INVX1 INVX1_70 ( .A(i_add_term2[16]), .Y(_106_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term1[16]), .B(_106_), .Y(_107_) );
INVX1 INVX1_71 ( .A(i_add_term1[17]), .Y(_108_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[17]), .B(_108_), .Y(_109_) );
INVX1 INVX1_72 ( .A(i_add_term2[17]), .Y(_110_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term1[17]), .B(_110_), .Y(_111_) );
OAI22X1 OAI22X1_5 ( .A(_105_), .B(_107_), .C(_109_), .D(_111_), .Y(_112_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_113_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_114_) );
NOR2X1 NOR2X1_83 ( .A(_113_), .B(_114_), .Y(_115_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_116_) );
NAND2X1 NAND2X1_101 ( .A(_115_), .B(_116_), .Y(_117_) );
NOR2X1 NOR2X1_84 ( .A(_112_), .B(_117_), .Y(_15_) );
INVX1 INVX1_73 ( .A(_13_), .Y(_118_) );
NAND2X1 NAND2X1_102 ( .A(gnd), .B(_15_), .Y(_119_) );
OAI21X1 OAI21X1_98 ( .A(_15_), .B(_118_), .C(_119_), .Y(w_cout_5_) );
INVX1 INVX1_74 ( .A(i_add_term1[20]), .Y(_120_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[20]), .B(_120_), .Y(_121_) );
INVX1 INVX1_75 ( .A(i_add_term2[20]), .Y(_122_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term1[20]), .B(_122_), .Y(_123_) );
INVX1 INVX1_76 ( .A(i_add_term1[21]), .Y(_124_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[21]), .B(_124_), .Y(_125_) );
INVX1 INVX1_77 ( .A(i_add_term2[21]), .Y(_126_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term1[21]), .B(_126_), .Y(_127_) );
OAI22X1 OAI22X1_6 ( .A(_121_), .B(_123_), .C(_125_), .D(_127_), .Y(_128_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_129_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_130_) );
NOR2X1 NOR2X1_90 ( .A(_129_), .B(_130_), .Y(_131_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_132_) );
NAND2X1 NAND2X1_103 ( .A(_131_), .B(_132_), .Y(_133_) );
NOR2X1 NOR2X1_91 ( .A(_128_), .B(_133_), .Y(_18_) );
INVX1 INVX1_78 ( .A(_16_), .Y(_134_) );
NAND2X1 NAND2X1_104 ( .A(gnd), .B(_18_), .Y(_135_) );
OAI21X1 OAI21X1_99 ( .A(_18_), .B(_134_), .C(_135_), .Y(w_cout_6_) );
INVX1 INVX1_79 ( .A(i_add_term1[24]), .Y(_136_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[24]), .B(_136_), .Y(_137_) );
INVX1 INVX1_80 ( .A(i_add_term2[24]), .Y(_138_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term1[24]), .B(_138_), .Y(_139_) );
INVX1 INVX1_81 ( .A(i_add_term1[25]), .Y(_140_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[25]), .B(_140_), .Y(_141_) );
INVX1 INVX1_82 ( .A(i_add_term2[25]), .Y(_142_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term1[25]), .B(_142_), .Y(_143_) );
OAI22X1 OAI22X1_7 ( .A(_137_), .B(_139_), .C(_141_), .D(_143_), .Y(_144_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_145_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_146_) );
NOR2X1 NOR2X1_97 ( .A(_145_), .B(_146_), .Y(_147_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_148_) );
NAND2X1 NAND2X1_105 ( .A(_147_), .B(_148_), .Y(_149_) );
NOR2X1 NOR2X1_98 ( .A(_144_), .B(_149_), .Y(_21_) );
INVX1 INVX1_83 ( .A(_19_), .Y(_150_) );
NAND2X1 NAND2X1_106 ( .A(gnd), .B(_21_), .Y(_151_) );
OAI21X1 OAI21X1_100 ( .A(_21_), .B(_150_), .C(_151_), .Y(w_cout_7_) );
INVX1 INVX1_84 ( .A(i_add_term1[28]), .Y(_152_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[28]), .B(_152_), .Y(_153_) );
INVX1 INVX1_85 ( .A(i_add_term2[28]), .Y(_154_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term1[28]), .B(_154_), .Y(_155_) );
INVX1 INVX1_86 ( .A(i_add_term1[29]), .Y(_156_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[29]), .B(_156_), .Y(_157_) );
INVX1 INVX1_87 ( .A(i_add_term2[29]), .Y(_158_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term1[29]), .B(_158_), .Y(_159_) );
OAI22X1 OAI22X1_8 ( .A(_153_), .B(_155_), .C(_157_), .D(_159_), .Y(_160_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_161_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_162_) );
NOR2X1 NOR2X1_104 ( .A(_161_), .B(_162_), .Y(_163_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_164_) );
NAND2X1 NAND2X1_107 ( .A(_163_), .B(_164_), .Y(_165_) );
NOR2X1 NOR2X1_105 ( .A(_160_), .B(_165_), .Y(_24_) );
INVX1 INVX1_88 ( .A(_22_), .Y(_166_) );
NAND2X1 NAND2X1_108 ( .A(gnd), .B(_24_), .Y(_167_) );
OAI21X1 OAI21X1_101 ( .A(_24_), .B(_166_), .C(_167_), .Y(w_cout_8_) );
INVX1 INVX1_89 ( .A(i_add_term1[32]), .Y(_168_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term2[32]), .B(_168_), .Y(_169_) );
INVX1 INVX1_90 ( .A(i_add_term2[32]), .Y(_170_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term1[32]), .B(_170_), .Y(_171_) );
INVX1 INVX1_91 ( .A(i_add_term1[33]), .Y(_172_) );
NOR2X1 NOR2X1_108 ( .A(i_add_term2[33]), .B(_172_), .Y(_173_) );
INVX1 INVX1_92 ( .A(i_add_term2[33]), .Y(_174_) );
NOR2X1 NOR2X1_109 ( .A(i_add_term1[33]), .B(_174_), .Y(_175_) );
OAI22X1 OAI22X1_9 ( .A(_169_), .B(_171_), .C(_173_), .D(_175_), .Y(_176_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_177_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_178_) );
NOR2X1 NOR2X1_111 ( .A(_177_), .B(_178_), .Y(_179_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_180_) );
NAND2X1 NAND2X1_109 ( .A(_179_), .B(_180_), .Y(_181_) );
NOR2X1 NOR2X1_112 ( .A(_176_), .B(_181_), .Y(_27_) );
INVX1 INVX1_93 ( .A(_25_), .Y(_182_) );
NAND2X1 NAND2X1_110 ( .A(gnd), .B(_27_), .Y(_183_) );
OAI21X1 OAI21X1_102 ( .A(_27_), .B(_182_), .C(_183_), .Y(w_cout_9_) );
INVX1 INVX1_94 ( .A(i_add_term1[36]), .Y(_184_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term2[36]), .B(_184_), .Y(_185_) );
INVX1 INVX1_95 ( .A(i_add_term2[36]), .Y(_186_) );
NOR2X1 NOR2X1_114 ( .A(i_add_term1[36]), .B(_186_), .Y(_187_) );
INVX1 INVX1_96 ( .A(i_add_term1[37]), .Y(_188_) );
NOR2X1 NOR2X1_115 ( .A(i_add_term2[37]), .B(_188_), .Y(_189_) );
INVX1 INVX1_97 ( .A(i_add_term2[37]), .Y(_190_) );
NOR2X1 NOR2X1_116 ( .A(i_add_term1[37]), .B(_190_), .Y(_191_) );
OAI22X1 OAI22X1_10 ( .A(_185_), .B(_187_), .C(_189_), .D(_191_), .Y(_192_) );
NOR2X1 NOR2X1_117 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_193_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_194_) );
NOR2X1 NOR2X1_118 ( .A(_193_), .B(_194_), .Y(_195_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_196_) );
NAND2X1 NAND2X1_111 ( .A(_195_), .B(_196_), .Y(_197_) );
NOR2X1 NOR2X1_119 ( .A(_192_), .B(_197_), .Y(_30_) );
INVX1 INVX1_98 ( .A(_28_), .Y(_198_) );
NAND2X1 NAND2X1_112 ( .A(gnd), .B(_30_), .Y(_199_) );
OAI21X1 OAI21X1_103 ( .A(_30_), .B(_198_), .C(_199_), .Y(w_cout_10_) );
INVX1 INVX1_99 ( .A(i_add_term1[40]), .Y(_200_) );
NOR2X1 NOR2X1_120 ( .A(i_add_term2[40]), .B(_200_), .Y(_201_) );
INVX1 INVX1_100 ( .A(i_add_term2[40]), .Y(_202_) );
NOR2X1 NOR2X1_121 ( .A(i_add_term1[40]), .B(_202_), .Y(_203_) );
INVX1 INVX1_101 ( .A(i_add_term1[41]), .Y(_204_) );
NOR2X1 NOR2X1_122 ( .A(i_add_term2[41]), .B(_204_), .Y(_205_) );
INVX1 INVX1_102 ( .A(i_add_term2[41]), .Y(_206_) );
NOR2X1 NOR2X1_123 ( .A(i_add_term1[41]), .B(_206_), .Y(_207_) );
OAI22X1 OAI22X1_11 ( .A(_201_), .B(_203_), .C(_205_), .D(_207_), .Y(_208_) );
NOR2X1 NOR2X1_124 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_209_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_210_) );
NOR2X1 NOR2X1_125 ( .A(_209_), .B(_210_), .Y(_211_) );
XOR2X1 XOR2X1_11 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_212_) );
NAND2X1 NAND2X1_113 ( .A(_211_), .B(_212_), .Y(_213_) );
NOR2X1 NOR2X1_126 ( .A(_208_), .B(_213_), .Y(_33_) );
INVX1 INVX1_103 ( .A(_31_), .Y(_214_) );
NAND2X1 NAND2X1_114 ( .A(gnd), .B(_33_), .Y(_215_) );
OAI21X1 OAI21X1_104 ( .A(_33_), .B(_214_), .C(_215_), .Y(w_cout_11_) );
INVX1 INVX1_104 ( .A(i_add_term1[44]), .Y(_216_) );
NOR2X1 NOR2X1_127 ( .A(i_add_term2[44]), .B(_216_), .Y(_217_) );
INVX1 INVX1_105 ( .A(i_add_term2[44]), .Y(_218_) );
NOR2X1 NOR2X1_128 ( .A(i_add_term1[44]), .B(_218_), .Y(_219_) );
INVX1 INVX1_106 ( .A(i_add_term1[45]), .Y(_220_) );
NOR2X1 NOR2X1_129 ( .A(i_add_term2[45]), .B(_220_), .Y(_221_) );
INVX1 INVX1_107 ( .A(i_add_term2[45]), .Y(_222_) );
NOR2X1 NOR2X1_130 ( .A(i_add_term1[45]), .B(_222_), .Y(_223_) );
OAI22X1 OAI22X1_12 ( .A(_217_), .B(_219_), .C(_221_), .D(_223_), .Y(_224_) );
NOR2X1 NOR2X1_131 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_225_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_226_) );
NOR2X1 NOR2X1_132 ( .A(_225_), .B(_226_), .Y(_227_) );
XOR2X1 XOR2X1_12 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_228_) );
NAND2X1 NAND2X1_115 ( .A(_227_), .B(_228_), .Y(_229_) );
NOR2X1 NOR2X1_133 ( .A(_224_), .B(_229_), .Y(_36_) );
INVX1 INVX1_108 ( .A(_34_), .Y(_230_) );
NAND2X1 NAND2X1_116 ( .A(gnd), .B(_36_), .Y(_231_) );
OAI21X1 OAI21X1_105 ( .A(_36_), .B(_230_), .C(_231_), .Y(w_cout_12_) );
INVX1 INVX1_109 ( .A(i_add_term1[48]), .Y(_232_) );
NOR2X1 NOR2X1_134 ( .A(i_add_term2[48]), .B(_232_), .Y(_233_) );
INVX1 INVX1_110 ( .A(i_add_term2[48]), .Y(_234_) );
NOR2X1 NOR2X1_135 ( .A(i_add_term1[48]), .B(_234_), .Y(_235_) );
INVX1 INVX1_111 ( .A(i_add_term1[49]), .Y(_236_) );
NOR2X1 NOR2X1_136 ( .A(i_add_term2[49]), .B(_236_), .Y(_237_) );
INVX1 INVX1_112 ( .A(i_add_term2[49]), .Y(_238_) );
NOR2X1 NOR2X1_137 ( .A(i_add_term1[49]), .B(_238_), .Y(_239_) );
OAI22X1 OAI22X1_13 ( .A(_233_), .B(_235_), .C(_237_), .D(_239_), .Y(_240_) );
NOR2X1 NOR2X1_138 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_241_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_242_) );
NOR2X1 NOR2X1_139 ( .A(_241_), .B(_242_), .Y(_243_) );
XOR2X1 XOR2X1_13 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_244_) );
NAND2X1 NAND2X1_117 ( .A(_243_), .B(_244_), .Y(_245_) );
NOR2X1 NOR2X1_140 ( .A(_240_), .B(_245_), .Y(_39_) );
INVX1 INVX1_113 ( .A(_37_), .Y(_246_) );
NAND2X1 NAND2X1_118 ( .A(gnd), .B(_39_), .Y(_247_) );
OAI21X1 OAI21X1_106 ( .A(_39_), .B(_246_), .C(_247_), .Y(cskip1_inst_cin) );
INVX1 INVX1_114 ( .A(gnd), .Y(_251_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_252_) );
NAND2X1 NAND2X1_119 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_253_) );
NAND3X1 NAND3X1_45 ( .A(_251_), .B(_253_), .C(_252_), .Y(_254_) );
NOR2X1 NOR2X1_141 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_248_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_249_) );
OAI21X1 OAI21X1_107 ( .A(_248_), .B(_249_), .C(gnd), .Y(_250_) );
NAND2X1 NAND2X1_120 ( .A(_250_), .B(_254_), .Y(_0__0_) );
OAI21X1 OAI21X1_108 ( .A(_251_), .B(_248_), .C(_253_), .Y(_2__1_) );
INVX1 INVX1_115 ( .A(_2__1_), .Y(_258_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_259_) );
NAND2X1 NAND2X1_121 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_260_) );
NAND3X1 NAND3X1_46 ( .A(_258_), .B(_260_), .C(_259_), .Y(_261_) );
NOR2X1 NOR2X1_142 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_255_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_256_) );
OAI21X1 OAI21X1_109 ( .A(_255_), .B(_256_), .C(_2__1_), .Y(_257_) );
NAND2X1 NAND2X1_122 ( .A(_257_), .B(_261_), .Y(_0__1_) );
OAI21X1 OAI21X1_110 ( .A(_258_), .B(_255_), .C(_260_), .Y(_2__2_) );
INVX1 INVX1_116 ( .A(_2__2_), .Y(_265_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_266_) );
NAND2X1 NAND2X1_123 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_267_) );
NAND3X1 NAND3X1_47 ( .A(_265_), .B(_267_), .C(_266_), .Y(_268_) );
NOR2X1 NOR2X1_143 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_262_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_263_) );
OAI21X1 OAI21X1_111 ( .A(_262_), .B(_263_), .C(_2__2_), .Y(_264_) );
NAND2X1 NAND2X1_124 ( .A(_264_), .B(_268_), .Y(_0__2_) );
OAI21X1 OAI21X1_112 ( .A(_265_), .B(_262_), .C(_267_), .Y(_2__3_) );
INVX1 INVX1_117 ( .A(_2__3_), .Y(_272_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_273_) );
NAND2X1 NAND2X1_125 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_274_) );
NAND3X1 NAND3X1_48 ( .A(_272_), .B(_274_), .C(_273_), .Y(_275_) );
NOR2X1 NOR2X1_144 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_269_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_270_) );
OAI21X1 OAI21X1_113 ( .A(_269_), .B(_270_), .C(_2__3_), .Y(_271_) );
NAND2X1 NAND2X1_126 ( .A(_271_), .B(_275_), .Y(_0__3_) );
OAI21X1 OAI21X1_114 ( .A(_272_), .B(_269_), .C(_274_), .Y(_1_) );
INVX1 INVX1_118 ( .A(w_cout_1_), .Y(_279_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_280_) );
NAND2X1 NAND2X1_127 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_281_) );
NAND3X1 NAND3X1_49 ( .A(_279_), .B(_281_), .C(_280_), .Y(_282_) );
NOR2X1 NOR2X1_145 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_276_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_277_) );
OAI21X1 OAI21X1_115 ( .A(_276_), .B(_277_), .C(w_cout_1_), .Y(_278_) );
NAND2X1 NAND2X1_128 ( .A(_278_), .B(_282_), .Y(_0__4_) );
OAI21X1 OAI21X1_116 ( .A(_279_), .B(_276_), .C(_281_), .Y(_5__1_) );
INVX1 INVX1_119 ( .A(_5__1_), .Y(_286_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_287_) );
NAND2X1 NAND2X1_129 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_288_) );
NAND3X1 NAND3X1_50 ( .A(_286_), .B(_288_), .C(_287_), .Y(_289_) );
NOR2X1 NOR2X1_146 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_283_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_284_) );
OAI21X1 OAI21X1_117 ( .A(_283_), .B(_284_), .C(_5__1_), .Y(_285_) );
NAND2X1 NAND2X1_130 ( .A(_285_), .B(_289_), .Y(_0__5_) );
OAI21X1 OAI21X1_118 ( .A(_286_), .B(_283_), .C(_288_), .Y(_5__2_) );
INVX1 INVX1_120 ( .A(_5__2_), .Y(_293_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_294_) );
NAND2X1 NAND2X1_131 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_295_) );
NAND3X1 NAND3X1_51 ( .A(_293_), .B(_295_), .C(_294_), .Y(_296_) );
NOR2X1 NOR2X1_147 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_290_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_291_) );
OAI21X1 OAI21X1_119 ( .A(_290_), .B(_291_), .C(_5__2_), .Y(_292_) );
NAND2X1 NAND2X1_132 ( .A(_292_), .B(_296_), .Y(_0__6_) );
OAI21X1 OAI21X1_120 ( .A(_293_), .B(_290_), .C(_295_), .Y(_5__3_) );
INVX1 INVX1_121 ( .A(_5__3_), .Y(_300_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_301_) );
NAND2X1 NAND2X1_133 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_302_) );
NAND3X1 NAND3X1_52 ( .A(_300_), .B(_302_), .C(_301_), .Y(_303_) );
NOR2X1 NOR2X1_148 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_297_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_298_) );
OAI21X1 OAI21X1_121 ( .A(_297_), .B(_298_), .C(_5__3_), .Y(_299_) );
NAND2X1 NAND2X1_134 ( .A(_299_), .B(_303_), .Y(_0__7_) );
OAI21X1 OAI21X1_122 ( .A(_300_), .B(_297_), .C(_302_), .Y(_4_) );
INVX1 INVX1_122 ( .A(w_cout_2_), .Y(_307_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_308_) );
NAND2X1 NAND2X1_135 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_309_) );
NAND3X1 NAND3X1_53 ( .A(_307_), .B(_309_), .C(_308_), .Y(_310_) );
NOR2X1 NOR2X1_149 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_304_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_305_) );
OAI21X1 OAI21X1_123 ( .A(_304_), .B(_305_), .C(w_cout_2_), .Y(_306_) );
NAND2X1 NAND2X1_136 ( .A(_306_), .B(_310_), .Y(_0__8_) );
BUFX2 BUFX2_55 ( .A(cskip1_inst_sum), .Y(_0__52_) );
BUFX2 BUFX2_56 ( .A(gnd), .Y(_2__0_) );
BUFX2 BUFX2_57 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_58 ( .A(w_cout_1_), .Y(_5__0_) );
BUFX2 BUFX2_59 ( .A(_4_), .Y(_5__4_) );
BUFX2 BUFX2_60 ( .A(w_cout_2_), .Y(_8__0_) );
BUFX2 BUFX2_61 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_62 ( .A(w_cout_3_), .Y(_11__0_) );
BUFX2 BUFX2_63 ( .A(_10_), .Y(_11__4_) );
BUFX2 BUFX2_64 ( .A(w_cout_4_), .Y(_14__0_) );
BUFX2 BUFX2_65 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_66 ( .A(w_cout_5_), .Y(_17__0_) );
BUFX2 BUFX2_67 ( .A(_16_), .Y(_17__4_) );
BUFX2 BUFX2_68 ( .A(w_cout_6_), .Y(_20__0_) );
BUFX2 BUFX2_69 ( .A(_19_), .Y(_20__4_) );
BUFX2 BUFX2_70 ( .A(w_cout_7_), .Y(_23__0_) );
BUFX2 BUFX2_71 ( .A(_22_), .Y(_23__4_) );
BUFX2 BUFX2_72 ( .A(w_cout_8_), .Y(_26__0_) );
BUFX2 BUFX2_73 ( .A(_25_), .Y(_26__4_) );
BUFX2 BUFX2_74 ( .A(w_cout_9_), .Y(_29__0_) );
BUFX2 BUFX2_75 ( .A(_28_), .Y(_29__4_) );
BUFX2 BUFX2_76 ( .A(w_cout_10_), .Y(_32__0_) );
BUFX2 BUFX2_77 ( .A(_31_), .Y(_32__4_) );
BUFX2 BUFX2_78 ( .A(w_cout_11_), .Y(_35__0_) );
BUFX2 BUFX2_79 ( .A(_34_), .Y(_35__4_) );
BUFX2 BUFX2_80 ( .A(w_cout_12_), .Y(_38__0_) );
BUFX2 BUFX2_81 ( .A(_37_), .Y(_38__4_) );
BUFX2 BUFX2_82 ( .A(cskip1_inst_cin), .Y(cskip1_inst_rca0_w_CARRY_0_) );
BUFX2 BUFX2_83 ( .A(cskip1_inst_cout0), .Y(cskip1_inst_rca0_w_CARRY_4_) );
BUFX2 BUFX2_84 ( .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_85 ( .A(cskip1_inst_cin), .Y(w_cout_13_) );
endmodule
