module cla_31bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [30:0] i_add1;
input [30:0] i_add2;
output [31:0] o_result;

NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_167_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_167_), .Y(w_C_1_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_168_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_168_), .Y(_169_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .C(_169_), .Y(_170_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_170_), .Y(w_C_2_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_0_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_2_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_2_), .C(_169_), .Y(_3_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_3_), .Y(w_C_3_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .Y(_4_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add1[3]), .Y(_5_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_5_), .Y(_6_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_7_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_7_), .C(_3_), .Y(_8_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_6_), .Y(w_C_4_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_9_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_10_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_10_), .C(_8_), .Y(_11_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_11_), .Y(w_C_5_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_12_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_12_), .C(_11_), .Y(_13_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .C(_13_), .Y(_14_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_14_), .Y(w_C_6_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .Y(_15_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add1[6]), .Y(_16_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_17_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_17_), .Y(_18_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_19_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_20_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_20_), .C(_13_), .Y(_21_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_16_), .C(_21_), .Y(w_C_7_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_16_), .Y(_22_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_23_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_24_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_24_), .Y(_25_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_25_), .C(_21_), .Y(_26_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .C(_26_), .Y(_27_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(w_C_8_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .Y(_28_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add1[8]), .Y(_29_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_30_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_31_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_32_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_32_), .Y(_33_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_33_), .C(_26_), .Y(_34_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_29_), .C(_34_), .Y(w_C_9_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_29_), .Y(_35_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_35_), .Y(_36_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_37_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_37_), .Y(_38_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_38_), .C(_34_), .Y(_39_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .C(_39_), .Y(_40_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_40_), .Y(w_C_10_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .Y(_41_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add1[10]), .Y(_42_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_43_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(_44_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_45_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_45_), .Y(_46_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_46_), .C(_39_), .Y(_47_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_42_), .C(_47_), .Y(w_C_11_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_42_), .Y(_48_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_48_), .Y(_49_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_50_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_50_), .Y(_51_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_51_), .C(_47_), .Y(_52_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .C(_52_), .Y(_53_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_53_), .Y(w_C_12_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .Y(_54_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add1[12]), .Y(_55_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_56_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_56_), .Y(_57_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_58_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_58_), .Y(_59_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_59_), .C(_52_), .Y(_60_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_55_), .C(_60_), .Y(w_C_13_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_55_), .Y(_61_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_61_), .Y(_62_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_63_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_63_), .Y(_64_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_64_), .C(_60_), .Y(_65_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .C(_65_), .Y(_66_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_66_), .Y(w_C_14_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .Y(_67_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add1[14]), .Y(_68_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_68_), .Y(_69_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(_70_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_71_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_71_), .Y(_72_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_73_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_73_), .Y(_74_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_74_), .C(_65_), .Y(_75_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_70_), .Y(_76_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_76_), .Y(w_C_15_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_77_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(_78_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_78_), .C(_75_), .Y(_79_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .C(_79_), .Y(_80_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_80_), .Y(w_C_16_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .Y(_81_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add1[16]), .Y(_82_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_82_), .Y(_83_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_83_), .Y(_84_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_85_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_85_), .Y(_86_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_87_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_87_), .Y(_88_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_88_), .C(_79_), .Y(_89_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_84_), .Y(_90_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_90_), .Y(w_C_17_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_91_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_91_), .Y(_92_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_92_), .C(_89_), .Y(_93_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .C(_93_), .Y(_94_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_94_), .Y(w_C_18_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .Y(_95_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add1[18]), .Y(_96_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_96_), .Y(_97_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_97_), .Y(_98_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_99_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_99_), .Y(_100_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_101_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_101_), .Y(_102_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_102_), .C(_93_), .Y(_103_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_98_), .Y(_104_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_104_), .Y(w_C_19_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_105_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_105_), .Y(_106_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_106_), .C(_103_), .Y(_107_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .C(_107_), .Y(_108_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_108_), .Y(w_C_20_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .Y(_109_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add1[20]), .Y(_110_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_110_), .Y(_111_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_111_), .Y(_112_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_113_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_113_), .Y(_114_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_115_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_115_), .Y(_116_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_116_), .C(_107_), .Y(_117_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_112_), .Y(_118_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_118_), .Y(w_C_21_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_119_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_119_), .Y(_120_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_120_), .C(_117_), .Y(_121_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .C(_121_), .Y(_122_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_122_), .Y(w_C_22_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .Y(_123_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add1[22]), .Y(_124_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_123_), .B(_124_), .Y(_125_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_125_), .Y(_126_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_127_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_127_), .Y(_128_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_129_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_129_), .Y(_130_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_130_), .C(_121_), .Y(_131_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_126_), .Y(_132_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(_132_), .Y(w_C_23_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_133_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_133_), .Y(_134_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_134_), .C(_131_), .Y(_135_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .C(_135_), .Y(_136_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(_136_), .Y(w_C_24_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_137_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_138_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_136_), .C(_137_), .Y(w_C_25_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_139_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_140_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_140_), .Y(_141_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_138_), .Y(_142_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_142_), .C(_135_), .Y(_143_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_144_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(_144_), .C(_143_), .Y(_145_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_139_), .Y(w_C_26_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .Y(_146_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add1[26]), .Y(_147_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_147_), .Y(_148_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_148_), .C(_145_), .Y(_149_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_147_), .C(_149_), .Y(w_C_27_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .Y(_150_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add1[27]), .Y(_151_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_151_), .Y(_152_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_153_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_154_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_154_), .C(_149_), .Y(_155_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_152_), .Y(w_C_28_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .Y(_156_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add1[28]), .Y(_157_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_157_), .Y(_158_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_158_), .C(_155_), .Y(_159_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_157_), .C(_159_), .Y(w_C_29_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_160_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_161_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_162_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_162_), .C(_159_), .Y(_163_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_160_), .Y(w_C_30_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_164_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_165_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_165_), .C(_163_), .Y(_166_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_166_), .Y(w_C_31_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_171__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_171__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_171__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_171__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_171__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_171__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_171__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_171__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_171__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_171__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_171__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_171__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_171__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_171__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_171__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_171__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_171__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_171__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_171__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_171__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_171__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_171__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_171__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_171__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_171__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_171__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_171__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_171__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_171__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_171__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_171__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(w_C_31_), .Y(o_result[31]) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_175_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_176_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_177_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_175_), .B(_177_), .C(_176_), .Y(_178_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_172_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_173_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_173_), .C(w_C_4_), .Y(_174_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_178_), .Y(_171__4_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_182_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_183_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_184_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_184_), .C(_183_), .Y(_185_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_179_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_180_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_180_), .C(w_C_5_), .Y(_181_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_185_), .Y(_171__5_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_189_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_190_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_191_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_191_), .C(_190_), .Y(_192_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_186_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_187_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_187_), .C(w_C_6_), .Y(_188_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_192_), .Y(_171__6_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_196_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_197_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_198_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_198_), .C(_197_), .Y(_199_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_193_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_194_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_194_), .C(w_C_7_), .Y(_195_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_199_), .Y(_171__7_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_203_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_204_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_205_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_205_), .C(_204_), .Y(_206_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_200_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_201_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_201_), .C(w_C_8_), .Y(_202_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_206_), .Y(_171__8_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_210_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_211_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_212_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_210_), .B(_212_), .C(_211_), .Y(_213_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_207_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_208_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_208_), .C(w_C_9_), .Y(_209_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_213_), .Y(_171__9_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_217_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_218_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_219_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_219_), .C(_218_), .Y(_220_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_214_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_215_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_215_), .C(w_C_10_), .Y(_216_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_220_), .Y(_171__10_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_224_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_225_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_226_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_226_), .C(_225_), .Y(_227_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_221_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_222_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_222_), .C(w_C_11_), .Y(_223_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_227_), .Y(_171__11_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(w_C_12_), .Y(_231_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_232_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_233_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_233_), .C(_232_), .Y(_234_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_228_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_229_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_229_), .C(w_C_12_), .Y(_230_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_234_), .Y(_171__12_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(w_C_13_), .Y(_238_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_239_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_240_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_238_), .B(_240_), .C(_239_), .Y(_241_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_235_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_236_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_236_), .C(w_C_13_), .Y(_237_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_241_), .Y(_171__13_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(w_C_14_), .Y(_245_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_246_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_247_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_247_), .C(_246_), .Y(_248_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_242_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_243_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_243_), .C(w_C_14_), .Y(_244_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_248_), .Y(_171__14_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(_252_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_253_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_254_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_254_), .C(_253_), .Y(_255_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_249_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_250_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_250_), .C(w_C_15_), .Y(_251_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_255_), .Y(_171__15_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(w_C_16_), .Y(_259_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_260_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_261_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_261_), .C(_260_), .Y(_262_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_256_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_257_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_257_), .C(w_C_16_), .Y(_258_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_262_), .Y(_171__16_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(w_C_17_), .Y(_266_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_267_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_268_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_268_), .C(_267_), .Y(_269_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_263_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_264_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_264_), .C(w_C_17_), .Y(_265_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_269_), .Y(_171__17_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(w_C_18_), .Y(_273_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_274_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_275_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_275_), .C(_274_), .Y(_276_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_270_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_271_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_271_), .C(w_C_18_), .Y(_272_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_276_), .Y(_171__18_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(w_C_19_), .Y(_280_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_281_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_282_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_282_), .C(_281_), .Y(_283_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_277_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_278_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_278_), .C(w_C_19_), .Y(_279_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_279_), .B(_283_), .Y(_171__19_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(w_C_20_), .Y(_287_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_288_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_289_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_287_), .B(_289_), .C(_288_), .Y(_290_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_284_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_285_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_285_), .C(w_C_20_), .Y(_286_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_290_), .Y(_171__20_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(w_C_21_), .Y(_294_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_295_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_296_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_296_), .C(_295_), .Y(_297_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_291_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_292_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_292_), .C(w_C_21_), .Y(_293_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_297_), .Y(_171__21_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(w_C_22_), .Y(_301_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_302_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_303_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_303_), .C(_302_), .Y(_304_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_298_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_299_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_299_), .C(w_C_22_), .Y(_300_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_304_), .Y(_171__22_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(w_C_23_), .Y(_308_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_309_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_310_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_310_), .C(_309_), .Y(_311_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_305_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_306_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_306_), .C(w_C_23_), .Y(_307_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_311_), .Y(_171__23_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(w_C_24_), .Y(_315_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_316_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_317_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_317_), .C(_316_), .Y(_318_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_312_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_313_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_313_), .C(w_C_24_), .Y(_314_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_318_), .Y(_171__24_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(w_C_25_), .Y(_322_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_323_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_324_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_324_), .C(_323_), .Y(_325_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_319_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_320_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_320_), .C(w_C_25_), .Y(_321_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_325_), .Y(_171__25_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(w_C_26_), .Y(_329_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_330_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_331_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_331_), .C(_330_), .Y(_332_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_326_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_327_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_327_), .C(w_C_26_), .Y(_328_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_332_), .Y(_171__26_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(w_C_27_), .Y(_336_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_337_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_338_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_338_), .C(_337_), .Y(_339_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_333_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_334_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_334_), .C(w_C_27_), .Y(_335_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_335_), .B(_339_), .Y(_171__27_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(w_C_28_), .Y(_343_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_344_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_345_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_345_), .C(_344_), .Y(_346_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_340_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_341_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_341_), .C(w_C_28_), .Y(_342_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_346_), .Y(_171__28_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(w_C_29_), .Y(_350_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_351_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_352_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_352_), .C(_351_), .Y(_353_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_347_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_348_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_348_), .C(w_C_29_), .Y(_349_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_353_), .Y(_171__29_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(w_C_30_), .Y(_357_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_358_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_359_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_359_), .C(_358_), .Y(_360_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_354_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_355_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_355_), .C(w_C_30_), .Y(_356_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_360_), .Y(_171__30_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_364_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_365_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_366_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_366_), .C(_365_), .Y(_367_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_361_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_362_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_362_), .C(gnd), .Y(_363_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_367_), .Y(_171__0_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_371_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_372_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_373_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_373_), .C(_372_), .Y(_374_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_368_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_369_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_369_), .C(w_C_1_), .Y(_370_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_374_), .Y(_171__1_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_378_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_379_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_380_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_380_), .C(_379_), .Y(_381_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_375_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_376_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_376_), .C(w_C_2_), .Y(_377_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_381_), .Y(_171__2_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_385_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_386_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_387_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_385_), .B(_387_), .C(_386_), .Y(_388_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_382_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_383_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_382_), .B(_383_), .C(w_C_3_), .Y(_384_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_388_), .Y(_171__3_) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(w_C_31_), .Y(_171__31_) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
