module CSkipA_11bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_2_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_5_) );
OAI21X1 OAI21X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .C(1'b0), .Y(_6_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_7_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_8_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_9_) );
NAND3X1 NAND3X1_1 ( .A(_7_), .B(_8_), .C(_9_), .Y(_10_) );
OAI21X1 OAI21X1_2 ( .A(_6_), .B(_10_), .C(_5_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3_), .Y(_11_) );
OAI21X1 OAI21X1_3 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .C(1'b0), .Y(_12_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_13_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_14_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_15_) );
NAND3X1 NAND3X1_2 ( .A(_13_), .B(_14_), .C(_15_), .Y(_16_) );
OAI21X1 OAI21X1_4 ( .A(_12_), .B(_16_), .C(_11_), .Y(w_cout_2_) );
INVX1 INVX1_3 ( .A(skip0_cin_next), .Y(_20_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_21_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_22_) );
NAND3X1 NAND3X1_3 ( .A(_20_), .B(_22_), .C(_21_), .Y(_23_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_17_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_18_) );
OAI21X1 OAI21X1_5 ( .A(_17_), .B(_18_), .C(skip0_cin_next), .Y(_19_) );
NAND2X1 NAND2X1_2 ( .A(_19_), .B(_23_), .Y(_0__4_) );
OAI21X1 OAI21X1_6 ( .A(_20_), .B(_17_), .C(_22_), .Y(_2__1_) );
INVX1 INVX1_4 ( .A(_2__1_), .Y(_27_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_28_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_29_) );
NAND3X1 NAND3X1_4 ( .A(_27_), .B(_29_), .C(_28_), .Y(_30_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_24_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_25_) );
OAI21X1 OAI21X1_7 ( .A(_24_), .B(_25_), .C(_2__1_), .Y(_26_) );
NAND2X1 NAND2X1_4 ( .A(_26_), .B(_30_), .Y(_0__5_) );
OAI21X1 OAI21X1_8 ( .A(_27_), .B(_24_), .C(_29_), .Y(_2__2_) );
INVX1 INVX1_5 ( .A(_2__2_), .Y(_34_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_35_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_36_) );
NAND3X1 NAND3X1_5 ( .A(_34_), .B(_36_), .C(_35_), .Y(_37_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_31_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_32_) );
OAI21X1 OAI21X1_9 ( .A(_31_), .B(_32_), .C(_2__2_), .Y(_33_) );
NAND2X1 NAND2X1_6 ( .A(_33_), .B(_37_), .Y(_0__6_) );
OAI21X1 OAI21X1_10 ( .A(_34_), .B(_31_), .C(_36_), .Y(_2__3_) );
INVX1 INVX1_6 ( .A(_2__3_), .Y(_41_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_42_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_43_) );
NAND3X1 NAND3X1_6 ( .A(_41_), .B(_43_), .C(_42_), .Y(_44_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_38_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_39_) );
OAI21X1 OAI21X1_11 ( .A(_38_), .B(_39_), .C(_2__3_), .Y(_40_) );
NAND2X1 NAND2X1_8 ( .A(_40_), .B(_44_), .Y(_0__7_) );
OAI21X1 OAI21X1_12 ( .A(_41_), .B(_38_), .C(_43_), .Y(_1_) );
INVX1 INVX1_7 ( .A(w_cout_1_), .Y(_48_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_49_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_50_) );
NAND3X1 NAND3X1_7 ( .A(_48_), .B(_50_), .C(_49_), .Y(_51_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_45_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_46_) );
OAI21X1 OAI21X1_13 ( .A(_45_), .B(_46_), .C(w_cout_1_), .Y(_47_) );
NAND2X1 NAND2X1_10 ( .A(_47_), .B(_51_), .Y(_0__8_) );
OAI21X1 OAI21X1_14 ( .A(_48_), .B(_45_), .C(_50_), .Y(_4__1_) );
INVX1 INVX1_8 ( .A(_4__1_), .Y(_55_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_56_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_57_) );
NAND3X1 NAND3X1_8 ( .A(_55_), .B(_57_), .C(_56_), .Y(_58_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_52_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_53_) );
OAI21X1 OAI21X1_15 ( .A(_52_), .B(_53_), .C(_4__1_), .Y(_54_) );
NAND2X1 NAND2X1_12 ( .A(_54_), .B(_58_), .Y(_0__9_) );
OAI21X1 OAI21X1_16 ( .A(_55_), .B(_52_), .C(_57_), .Y(_4__2_) );
INVX1 INVX1_9 ( .A(_4__2_), .Y(_62_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_63_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_64_) );
NAND3X1 NAND3X1_9 ( .A(_62_), .B(_64_), .C(_63_), .Y(_65_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_59_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_60_) );
OAI21X1 OAI21X1_17 ( .A(_59_), .B(_60_), .C(_4__2_), .Y(_61_) );
NAND2X1 NAND2X1_14 ( .A(_61_), .B(_65_), .Y(_0__10_) );
OAI21X1 OAI21X1_18 ( .A(_62_), .B(_59_), .C(_64_), .Y(_4__3_) );
INVX1 INVX1_10 ( .A(_4__3_), .Y(_69_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_70_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_71_) );
NAND3X1 NAND3X1_10 ( .A(_69_), .B(_71_), .C(_70_), .Y(_72_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_66_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_67_) );
OAI21X1 OAI21X1_19 ( .A(_66_), .B(_67_), .C(_4__3_), .Y(_68_) );
NAND2X1 NAND2X1_16 ( .A(_68_), .B(_72_), .Y(_0__11_) );
OAI21X1 OAI21X1_20 ( .A(_69_), .B(_66_), .C(_71_), .Y(_3_) );
INVX1 INVX1_11 ( .A(1'b0), .Y(_76_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_77_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_78_) );
NAND3X1 NAND3X1_11 ( .A(_76_), .B(_78_), .C(_77_), .Y(_79_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_73_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_74_) );
OAI21X1 OAI21X1_21 ( .A(_73_), .B(_74_), .C(1'b0), .Y(_75_) );
NAND2X1 NAND2X1_18 ( .A(_75_), .B(_79_), .Y(_0__0_) );
OAI21X1 OAI21X1_22 ( .A(_76_), .B(_73_), .C(_78_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_12 ( .A(rca_inst_w_CARRY_1_), .Y(_83_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_84_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_85_) );
NAND3X1 NAND3X1_12 ( .A(_83_), .B(_85_), .C(_84_), .Y(_86_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_80_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_81_) );
OAI21X1 OAI21X1_23 ( .A(_80_), .B(_81_), .C(rca_inst_w_CARRY_1_), .Y(_82_) );
NAND2X1 NAND2X1_20 ( .A(_82_), .B(_86_), .Y(_0__1_) );
OAI21X1 OAI21X1_24 ( .A(_83_), .B(_80_), .C(_85_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_13 ( .A(rca_inst_w_CARRY_2_), .Y(_90_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_91_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_92_) );
NAND3X1 NAND3X1_13 ( .A(_90_), .B(_92_), .C(_91_), .Y(_93_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_87_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_88_) );
OAI21X1 OAI21X1_25 ( .A(_87_), .B(_88_), .C(rca_inst_w_CARRY_2_), .Y(_89_) );
NAND2X1 NAND2X1_22 ( .A(_89_), .B(_93_), .Y(_0__2_) );
OAI21X1 OAI21X1_26 ( .A(_90_), .B(_87_), .C(_92_), .Y(rca_inst_w_CARRY_3_) );
INVX1 INVX1_14 ( .A(rca_inst_w_CARRY_3_), .Y(_97_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_98_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_99_) );
NAND3X1 NAND3X1_14 ( .A(_97_), .B(_99_), .C(_98_), .Y(_100_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_94_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_95_) );
OAI21X1 OAI21X1_27 ( .A(_94_), .B(_95_), .C(rca_inst_w_CARRY_3_), .Y(_96_) );
NAND2X1 NAND2X1_24 ( .A(_96_), .B(_100_), .Y(_0__3_) );
OAI21X1 OAI21X1_28 ( .A(_97_), .B(_94_), .C(_99_), .Y(cout0) );
INVX1 INVX1_15 ( .A(cout0), .Y(_101_) );
OAI21X1 OAI21X1_29 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .C(1'b0), .Y(_102_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_103_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_104_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_105_) );
NAND3X1 NAND3X1_15 ( .A(_103_), .B(_104_), .C(_105_), .Y(_106_) );
OAI21X1 OAI21X1_30 ( .A(_102_), .B(_106_), .C(_101_), .Y(skip0_cin_next) );
BUFX2 BUFX2_14 ( .A(skip0_cin_next), .Y(_2__0_) );
BUFX2 BUFX2_15 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_16 ( .A(w_cout_1_), .Y(_4__0_) );
BUFX2 BUFX2_17 ( .A(_3_), .Y(_4__4_) );
BUFX2 BUFX2_18 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_19 ( .A(cout0), .Y(rca_inst_w_CARRY_4_) );
BUFX2 BUFX2_20 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
