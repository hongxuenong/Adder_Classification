module cla_22bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [21:0] i_add1;
input [21:0] i_add2;
output [22:0] o_result;

NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_85_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_85_), .Y(w_C_1_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_86_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_87_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_87_), .Y(w_C_2_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .Y(_88_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add1[2]), .Y(_89_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_89_), .Y(_90_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_91_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_87_), .C(_91_), .Y(_92_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_90_), .Y(w_C_3_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_93_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_94_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_94_), .C(_92_), .Y(_95_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_93_), .Y(_96_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_96_), .Y(w_C_4_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_97_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_98_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_96_), .C(_97_), .Y(w_C_5_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_99_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_99_), .Y(_100_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_98_), .Y(_101_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_97_), .C(_95_), .Y(_102_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_103_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_103_), .Y(_104_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_104_), .C(_102_), .Y(_105_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_100_), .Y(_106_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_106_), .Y(w_C_6_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_107_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_107_), .Y(_108_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_109_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_106_), .C(_108_), .Y(w_C_7_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .Y(_110_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add1[7]), .Y(_0_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_109_), .Y(_1_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_108_), .C(_105_), .Y(_2_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_3_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_3_), .Y(_4_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_4_), .C(_2_), .Y(_5_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_0_), .C(_5_), .Y(w_C_8_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_0_), .Y(_6_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_6_), .Y(_7_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_8_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_8_), .Y(_9_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_9_), .C(_5_), .Y(_10_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .C(_10_), .Y(_11_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(w_C_9_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .Y(_12_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add1[9]), .Y(_13_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_14_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_14_), .Y(_15_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_16_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_17_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_17_), .C(_10_), .Y(_18_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_13_), .C(_18_), .Y(w_C_10_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_13_), .Y(_19_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_20_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_21_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_21_), .Y(_22_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_22_), .C(_18_), .Y(_23_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .C(_23_), .Y(_24_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_24_), .Y(w_C_11_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .Y(_25_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add1[11]), .Y(_26_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_27_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(_28_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_29_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_29_), .Y(_30_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_30_), .C(_23_), .Y(_31_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_26_), .C(_31_), .Y(w_C_12_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_26_), .Y(_32_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_32_), .Y(_33_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_34_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_34_), .Y(_35_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_35_), .C(_31_), .Y(_36_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .C(_36_), .Y(_37_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_37_), .Y(w_C_13_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .Y(_38_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add1[13]), .Y(_39_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_40_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_40_), .Y(_41_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_42_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_42_), .Y(_43_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_43_), .C(_36_), .Y(_44_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_39_), .C(_44_), .Y(w_C_14_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_39_), .Y(_45_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_45_), .Y(_46_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_47_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_47_), .Y(_48_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_48_), .C(_44_), .Y(_49_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .C(_49_), .Y(_50_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_50_), .Y(w_C_15_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .Y(_51_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add1[15]), .Y(_52_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_53_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_53_), .Y(_54_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_55_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_55_), .Y(_56_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_56_), .C(_49_), .Y(_57_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_52_), .C(_57_), .Y(w_C_16_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_58_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_58_), .Y(_59_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_52_), .Y(_60_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_60_), .Y(_61_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_62_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_62_), .C(_57_), .Y(_63_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_59_), .Y(w_C_17_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .Y(_64_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add1[17]), .Y(_65_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_65_), .Y(_66_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_66_), .C(_63_), .Y(_67_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_65_), .C(_67_), .Y(w_C_18_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .Y(_68_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add1[18]), .Y(_69_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_69_), .Y(_70_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_71_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_72_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_72_), .C(_67_), .Y(_73_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_70_), .Y(w_C_19_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .Y(_74_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add1[19]), .Y(_75_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_75_), .Y(_76_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_76_), .C(_73_), .Y(_77_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_75_), .C(_77_), .Y(w_C_20_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_78_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_79_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_80_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_80_), .C(_77_), .Y(_81_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_78_), .Y(w_C_21_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_82_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_83_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_83_), .C(_81_), .Y(_84_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_84_), .Y(w_C_22_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_111__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_111__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_111__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_111__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_111__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_111__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_111__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_111__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_111__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_111__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_111__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_111__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_111__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_111__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_111__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_111__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_111__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_111__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_111__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_111__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_111__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_111__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(w_C_22_), .Y(o_result[22]) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_115_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_116_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_117_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_117_), .C(_116_), .Y(_118_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_112_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_113_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_113_), .C(w_C_4_), .Y(_114_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_118_), .Y(_111__4_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_122_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_123_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_124_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_124_), .C(_123_), .Y(_125_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_119_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_120_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_120_), .C(w_C_5_), .Y(_121_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_125_), .Y(_111__5_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_129_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_130_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_131_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_129_), .B(_131_), .C(_130_), .Y(_132_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_126_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_127_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_127_), .C(w_C_6_), .Y(_128_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_132_), .Y(_111__6_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_136_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_137_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_138_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_138_), .C(_137_), .Y(_139_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_133_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_134_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_134_), .C(w_C_7_), .Y(_135_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_139_), .Y(_111__7_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_143_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_144_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_145_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_145_), .C(_144_), .Y(_146_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_140_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_141_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_141_), .C(w_C_8_), .Y(_142_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_146_), .Y(_111__8_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_150_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_151_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_152_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_152_), .C(_151_), .Y(_153_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_147_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_148_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_148_), .C(w_C_9_), .Y(_149_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_153_), .Y(_111__9_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_157_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_158_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_159_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_159_), .C(_158_), .Y(_160_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_154_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_155_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_155_), .C(w_C_10_), .Y(_156_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_160_), .Y(_111__10_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_164_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_165_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_166_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_166_), .C(_165_), .Y(_167_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_161_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_162_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_162_), .C(w_C_11_), .Y(_163_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_167_), .Y(_111__11_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(w_C_12_), .Y(_171_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_172_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_173_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_173_), .C(_172_), .Y(_174_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_168_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_169_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_169_), .C(w_C_12_), .Y(_170_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_174_), .Y(_111__12_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(w_C_13_), .Y(_178_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_179_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_180_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_180_), .C(_179_), .Y(_181_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_175_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_176_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_175_), .B(_176_), .C(w_C_13_), .Y(_177_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_181_), .Y(_111__13_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(w_C_14_), .Y(_185_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_186_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_187_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_187_), .C(_186_), .Y(_188_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_182_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_183_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_183_), .C(w_C_14_), .Y(_184_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_188_), .Y(_111__14_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(_192_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_193_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_194_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(_194_), .C(_193_), .Y(_195_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_189_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_190_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_190_), .C(w_C_15_), .Y(_191_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_195_), .Y(_111__15_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(w_C_16_), .Y(_199_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_200_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_201_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_201_), .C(_200_), .Y(_202_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_196_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_197_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_197_), .C(w_C_16_), .Y(_198_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_202_), .Y(_111__16_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(w_C_17_), .Y(_206_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_207_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_208_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_208_), .C(_207_), .Y(_209_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_203_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_204_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_204_), .C(w_C_17_), .Y(_205_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_209_), .Y(_111__17_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(w_C_18_), .Y(_213_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_214_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_215_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_215_), .C(_214_), .Y(_216_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_210_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_211_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_210_), .B(_211_), .C(w_C_18_), .Y(_212_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_216_), .Y(_111__18_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(w_C_19_), .Y(_220_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_221_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_222_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_222_), .C(_221_), .Y(_223_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_217_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_218_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_218_), .C(w_C_19_), .Y(_219_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_223_), .Y(_111__19_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(w_C_20_), .Y(_227_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_228_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_229_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_229_), .C(_228_), .Y(_230_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_224_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_225_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_225_), .C(w_C_20_), .Y(_226_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_230_), .Y(_111__20_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(w_C_21_), .Y(_234_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_235_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_236_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_236_), .C(_235_), .Y(_237_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_231_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_232_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_232_), .C(w_C_21_), .Y(_233_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_237_), .Y(_111__21_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_241_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_242_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_243_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_243_), .C(_242_), .Y(_244_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_238_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_239_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_238_), .B(_239_), .C(gnd), .Y(_240_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_244_), .Y(_111__0_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_248_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_249_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_250_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_250_), .C(_249_), .Y(_251_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_245_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_246_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_246_), .C(w_C_1_), .Y(_247_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_251_), .Y(_111__1_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_255_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_256_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_257_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_257_), .C(_256_), .Y(_258_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_252_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_253_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_253_), .C(w_C_2_), .Y(_254_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_258_), .Y(_111__2_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_262_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_263_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_264_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_264_), .C(_263_), .Y(_265_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_259_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_260_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_260_), .C(w_C_3_), .Y(_261_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_265_), .Y(_111__3_) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(w_C_22_), .Y(_111__22_) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
