module cla_37bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add1[19], i_add1[20], i_add1[21], i_add1[22], i_add1[23], i_add1[24], i_add1[25], i_add1[26], i_add1[27], i_add1[28], i_add1[29], i_add1[30], i_add1[31], i_add1[32], i_add1[33], i_add1[34], i_add1[35], i_add1[36], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], i_add2[19], i_add2[20], i_add2[21], i_add2[22], i_add2[23], i_add2[24], i_add2[25], i_add2[26], i_add2[27], i_add2[28], i_add2[29], i_add2[30], i_add2[31], i_add2[32], i_add2[33], i_add2[34], i_add2[35], i_add2[36], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21], o_result[22], o_result[23], o_result[24], o_result[25], o_result[26], o_result[27], o_result[28], o_result[29], o_result[30], o_result[31], o_result[32], o_result[33], o_result[34], o_result[35], o_result[36], o_result[37]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add1[19];
input i_add1[20];
input i_add1[21];
input i_add1[22];
input i_add1[23];
input i_add1[24];
input i_add1[25];
input i_add1[26];
input i_add1[27];
input i_add1[28];
input i_add1[29];
input i_add1[30];
input i_add1[31];
input i_add1[32];
input i_add1[33];
input i_add1[34];
input i_add1[35];
input i_add1[36];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
input i_add2[19];
input i_add2[20];
input i_add2[21];
input i_add2[22];
input i_add2[23];
input i_add2[24];
input i_add2[25];
input i_add2[26];
input i_add2[27];
input i_add2[28];
input i_add2[29];
input i_add2[30];
input i_add2[31];
input i_add2[32];
input i_add2[33];
input i_add2[34];
input i_add2[35];
input i_add2[36];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];
output o_result[22];
output o_result[23];
output o_result[24];
output o_result[25];
output o_result[26];
output o_result[27];
output o_result[28];
output o_result[29];
output o_result[30];
output o_result[31];
output o_result[32];
output o_result[33];
output o_result[34];
output o_result[35];
output o_result[36];
output o_result[37];

OR2X2 OR2X2_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_436_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_437_) );
NAND3X1 NAND3X1_1 ( .A(_435_), .B(_437_), .C(_436_), .Y(_438_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_432_) );
AND2X2 AND2X2_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_433_) );
OAI21X1 OAI21X1_1 ( .A(_432_), .B(_433_), .C(1'b0), .Y(_434_) );
NAND2X1 NAND2X1_2 ( .A(_434_), .B(_438_), .Y(_200__0_) );
INVX1 INVX1_1 ( .A(w_C_1_), .Y(_442_) );
OR2X2 OR2X2_2 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_443_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_444_) );
NAND3X1 NAND3X1_2 ( .A(_442_), .B(_444_), .C(_443_), .Y(_445_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_439_) );
AND2X2 AND2X2_2 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_440_) );
OAI21X1 OAI21X1_2 ( .A(_439_), .B(_440_), .C(w_C_1_), .Y(_441_) );
NAND2X1 NAND2X1_4 ( .A(_441_), .B(_445_), .Y(_200__1_) );
INVX1 INVX1_2 ( .A(w_C_2_), .Y(_449_) );
OR2X2 OR2X2_3 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_450_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_451_) );
NAND3X1 NAND3X1_3 ( .A(_449_), .B(_451_), .C(_450_), .Y(_452_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_446_) );
AND2X2 AND2X2_3 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_447_) );
OAI21X1 OAI21X1_3 ( .A(_446_), .B(_447_), .C(w_C_2_), .Y(_448_) );
NAND2X1 NAND2X1_6 ( .A(_448_), .B(_452_), .Y(_200__2_) );
INVX1 INVX1_3 ( .A(w_C_3_), .Y(_456_) );
OR2X2 OR2X2_4 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_457_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_458_) );
NAND3X1 NAND3X1_4 ( .A(_456_), .B(_458_), .C(_457_), .Y(_459_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_453_) );
AND2X2 AND2X2_4 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_454_) );
OAI21X1 OAI21X1_4 ( .A(_453_), .B(_454_), .C(w_C_3_), .Y(_455_) );
NAND2X1 NAND2X1_8 ( .A(_455_), .B(_459_), .Y(_200__3_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_4 ( .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_11 ( .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_5 ( .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_5 ( .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_5 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_6 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_5 ( .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_13 ( .A(_4_), .B(_7_), .Y(w_C_3_) );
OR2X2 OR2X2_7 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_6 ( .A(_4_), .B(_9_), .C(_7_), .Y(_10_) );
AND2X2 AND2X2_5 ( .A(_10_), .B(_8_), .Y(w_C_4_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
OR2X2 OR2X2_8 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_12_) );
NAND3X1 NAND3X1_7 ( .A(_8_), .B(_12_), .C(_10_), .Y(_13_) );
NAND2X1 NAND2X1_16 ( .A(_11_), .B(_13_), .Y(w_C_5_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_14_) );
INVX1 INVX1_6 ( .A(_14_), .Y(_15_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_16_) );
NAND3X1 NAND3X1_8 ( .A(_11_), .B(_16_), .C(_13_), .Y(_17_) );
AND2X2 AND2X2_6 ( .A(_17_), .B(_15_), .Y(w_C_6_) );
AND2X2 AND2X2_7 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_18_) );
INVX1 INVX1_7 ( .A(_18_), .Y(_19_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_20_) );
INVX1 INVX1_8 ( .A(_20_), .Y(_21_) );
NAND3X1 NAND3X1_9 ( .A(_15_), .B(_21_), .C(_17_), .Y(_22_) );
AND2X2 AND2X2_8 ( .A(_22_), .B(_19_), .Y(_23_) );
INVX1 INVX1_9 ( .A(_23_), .Y(w_C_7_) );
AND2X2 AND2X2_9 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_24_) );
INVX1 INVX1_10 ( .A(_24_), .Y(_25_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_26_) );
OAI21X1 OAI21X1_6 ( .A(_26_), .B(_23_), .C(_25_), .Y(w_C_8_) );
AND2X2 AND2X2_10 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_27_) );
INVX1 INVX1_11 ( .A(_27_), .Y(_28_) );
INVX1 INVX1_12 ( .A(_26_), .Y(_29_) );
NAND3X1 NAND3X1_10 ( .A(_19_), .B(_25_), .C(_22_), .Y(_30_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_31_) );
INVX1 INVX1_13 ( .A(_31_), .Y(_32_) );
NAND3X1 NAND3X1_11 ( .A(_29_), .B(_32_), .C(_30_), .Y(_33_) );
AND2X2 AND2X2_11 ( .A(_33_), .B(_28_), .Y(_34_) );
INVX1 INVX1_14 ( .A(_34_), .Y(w_C_9_) );
AND2X2 AND2X2_12 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_35_) );
INVX1 INVX1_15 ( .A(_35_), .Y(_36_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_37_) );
OAI21X1 OAI21X1_7 ( .A(_37_), .B(_34_), .C(_36_), .Y(w_C_10_) );
INVX1 INVX1_16 ( .A(i_add2[10]), .Y(_38_) );
INVX1 INVX1_17 ( .A(i_add1[10]), .Y(_39_) );
INVX1 INVX1_18 ( .A(_37_), .Y(_40_) );
NAND3X1 NAND3X1_12 ( .A(_28_), .B(_36_), .C(_33_), .Y(_41_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_42_) );
INVX1 INVX1_19 ( .A(_42_), .Y(_43_) );
NAND3X1 NAND3X1_13 ( .A(_40_), .B(_43_), .C(_41_), .Y(_44_) );
OAI21X1 OAI21X1_8 ( .A(_38_), .B(_39_), .C(_44_), .Y(w_C_11_) );
NOR2X1 NOR2X1_11 ( .A(_38_), .B(_39_), .Y(_45_) );
INVX1 INVX1_20 ( .A(_45_), .Y(_46_) );
AND2X2 AND2X2_13 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_47_) );
INVX1 INVX1_21 ( .A(_47_), .Y(_48_) );
NAND3X1 NAND3X1_14 ( .A(_46_), .B(_48_), .C(_44_), .Y(_49_) );
OAI21X1 OAI21X1_9 ( .A(i_add2[11]), .B(i_add1[11]), .C(_49_), .Y(_50_) );
INVX1 INVX1_22 ( .A(_50_), .Y(w_C_12_) );
INVX1 INVX1_23 ( .A(i_add2[12]), .Y(_51_) );
INVX1 INVX1_24 ( .A(i_add1[12]), .Y(_52_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_53_) );
INVX1 INVX1_25 ( .A(_53_), .Y(_54_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_55_) );
INVX1 INVX1_26 ( .A(_55_), .Y(_56_) );
NAND3X1 NAND3X1_15 ( .A(_54_), .B(_56_), .C(_49_), .Y(_57_) );
OAI21X1 OAI21X1_10 ( .A(_51_), .B(_52_), .C(_57_), .Y(w_C_13_) );
NOR2X1 NOR2X1_14 ( .A(_51_), .B(_52_), .Y(_58_) );
INVX1 INVX1_27 ( .A(_58_), .Y(_59_) );
AND2X2 AND2X2_14 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_60_) );
INVX1 INVX1_28 ( .A(_60_), .Y(_61_) );
NAND3X1 NAND3X1_16 ( .A(_59_), .B(_61_), .C(_57_), .Y(_62_) );
OAI21X1 OAI21X1_11 ( .A(i_add2[13]), .B(i_add1[13]), .C(_62_), .Y(_63_) );
INVX1 INVX1_29 ( .A(_63_), .Y(w_C_14_) );
INVX1 INVX1_30 ( .A(i_add2[14]), .Y(_64_) );
INVX1 INVX1_31 ( .A(i_add1[14]), .Y(_65_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_66_) );
INVX1 INVX1_32 ( .A(_66_), .Y(_67_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_68_) );
INVX1 INVX1_33 ( .A(_68_), .Y(_69_) );
NAND3X1 NAND3X1_17 ( .A(_67_), .B(_69_), .C(_62_), .Y(_70_) );
OAI21X1 OAI21X1_12 ( .A(_64_), .B(_65_), .C(_70_), .Y(w_C_15_) );
NOR2X1 NOR2X1_17 ( .A(_64_), .B(_65_), .Y(_71_) );
INVX1 INVX1_34 ( .A(_71_), .Y(_72_) );
AND2X2 AND2X2_15 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_73_) );
INVX1 INVX1_35 ( .A(_73_), .Y(_74_) );
NAND3X1 NAND3X1_18 ( .A(_72_), .B(_74_), .C(_70_), .Y(_75_) );
OAI21X1 OAI21X1_13 ( .A(i_add2[15]), .B(i_add1[15]), .C(_75_), .Y(_76_) );
INVX1 INVX1_36 ( .A(_76_), .Y(w_C_16_) );
INVX1 INVX1_37 ( .A(i_add2[16]), .Y(_77_) );
INVX1 INVX1_38 ( .A(i_add1[16]), .Y(_78_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_79_) );
INVX1 INVX1_39 ( .A(_79_), .Y(_80_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_81_) );
INVX1 INVX1_40 ( .A(_81_), .Y(_82_) );
NAND3X1 NAND3X1_19 ( .A(_80_), .B(_82_), .C(_75_), .Y(_83_) );
OAI21X1 OAI21X1_14 ( .A(_77_), .B(_78_), .C(_83_), .Y(w_C_17_) );
NOR2X1 NOR2X1_20 ( .A(_77_), .B(_78_), .Y(_84_) );
INVX1 INVX1_41 ( .A(_84_), .Y(_85_) );
AND2X2 AND2X2_16 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_86_) );
INVX1 INVX1_42 ( .A(_86_), .Y(_87_) );
NAND3X1 NAND3X1_20 ( .A(_85_), .B(_87_), .C(_83_), .Y(_88_) );
OAI21X1 OAI21X1_15 ( .A(i_add2[17]), .B(i_add1[17]), .C(_88_), .Y(_89_) );
INVX1 INVX1_43 ( .A(_89_), .Y(w_C_18_) );
INVX1 INVX1_44 ( .A(i_add2[18]), .Y(_90_) );
INVX1 INVX1_45 ( .A(i_add1[18]), .Y(_91_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_92_) );
INVX1 INVX1_46 ( .A(_92_), .Y(_93_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_94_) );
INVX1 INVX1_47 ( .A(_94_), .Y(_95_) );
NAND3X1 NAND3X1_21 ( .A(_93_), .B(_95_), .C(_88_), .Y(_96_) );
OAI21X1 OAI21X1_16 ( .A(_90_), .B(_91_), .C(_96_), .Y(w_C_19_) );
NOR2X1 NOR2X1_23 ( .A(_90_), .B(_91_), .Y(_97_) );
INVX1 INVX1_48 ( .A(_97_), .Y(_98_) );
AND2X2 AND2X2_17 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_99_) );
INVX1 INVX1_49 ( .A(_99_), .Y(_100_) );
NAND3X1 NAND3X1_22 ( .A(_98_), .B(_100_), .C(_96_), .Y(_101_) );
OAI21X1 OAI21X1_17 ( .A(i_add2[19]), .B(i_add1[19]), .C(_101_), .Y(_102_) );
INVX1 INVX1_50 ( .A(_102_), .Y(w_C_20_) );
INVX1 INVX1_51 ( .A(i_add2[20]), .Y(_103_) );
INVX1 INVX1_52 ( .A(i_add1[20]), .Y(_104_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_105_) );
INVX1 INVX1_53 ( .A(_105_), .Y(_106_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_107_) );
INVX1 INVX1_54 ( .A(_107_), .Y(_108_) );
NAND3X1 NAND3X1_23 ( .A(_106_), .B(_108_), .C(_101_), .Y(_109_) );
OAI21X1 OAI21X1_18 ( .A(_103_), .B(_104_), .C(_109_), .Y(w_C_21_) );
NOR2X1 NOR2X1_26 ( .A(_103_), .B(_104_), .Y(_110_) );
INVX1 INVX1_55 ( .A(_110_), .Y(_111_) );
AND2X2 AND2X2_18 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_112_) );
INVX1 INVX1_56 ( .A(_112_), .Y(_113_) );
NAND3X1 NAND3X1_24 ( .A(_111_), .B(_113_), .C(_109_), .Y(_114_) );
OAI21X1 OAI21X1_19 ( .A(i_add2[21]), .B(i_add1[21]), .C(_114_), .Y(_115_) );
INVX1 INVX1_57 ( .A(_115_), .Y(w_C_22_) );
INVX1 INVX1_58 ( .A(i_add2[22]), .Y(_116_) );
INVX1 INVX1_59 ( .A(i_add1[22]), .Y(_117_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_118_) );
INVX1 INVX1_60 ( .A(_118_), .Y(_119_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_120_) );
INVX1 INVX1_61 ( .A(_120_), .Y(_121_) );
NAND3X1 NAND3X1_25 ( .A(_119_), .B(_121_), .C(_114_), .Y(_122_) );
OAI21X1 OAI21X1_20 ( .A(_116_), .B(_117_), .C(_122_), .Y(w_C_23_) );
NOR2X1 NOR2X1_29 ( .A(_116_), .B(_117_), .Y(_123_) );
INVX1 INVX1_62 ( .A(_123_), .Y(_124_) );
AND2X2 AND2X2_19 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_125_) );
INVX1 INVX1_63 ( .A(_125_), .Y(_126_) );
NAND3X1 NAND3X1_26 ( .A(_124_), .B(_126_), .C(_122_), .Y(_127_) );
OAI21X1 OAI21X1_21 ( .A(i_add2[23]), .B(i_add1[23]), .C(_127_), .Y(_128_) );
INVX1 INVX1_64 ( .A(_128_), .Y(w_C_24_) );
INVX1 INVX1_65 ( .A(i_add2[24]), .Y(_129_) );
INVX1 INVX1_66 ( .A(i_add1[24]), .Y(_130_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_131_) );
INVX1 INVX1_67 ( .A(_131_), .Y(_132_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_133_) );
INVX1 INVX1_68 ( .A(_133_), .Y(_134_) );
NAND3X1 NAND3X1_27 ( .A(_132_), .B(_134_), .C(_127_), .Y(_135_) );
OAI21X1 OAI21X1_22 ( .A(_129_), .B(_130_), .C(_135_), .Y(w_C_25_) );
NOR2X1 NOR2X1_32 ( .A(_129_), .B(_130_), .Y(_136_) );
INVX1 INVX1_69 ( .A(_136_), .Y(_137_) );
AND2X2 AND2X2_20 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_138_) );
INVX1 INVX1_70 ( .A(_138_), .Y(_139_) );
NAND3X1 NAND3X1_28 ( .A(_137_), .B(_139_), .C(_135_), .Y(_140_) );
OAI21X1 OAI21X1_23 ( .A(i_add2[25]), .B(i_add1[25]), .C(_140_), .Y(_141_) );
INVX1 INVX1_71 ( .A(_141_), .Y(w_C_26_) );
INVX1 INVX1_72 ( .A(i_add2[26]), .Y(_142_) );
INVX1 INVX1_73 ( .A(i_add1[26]), .Y(_143_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_144_) );
INVX1 INVX1_74 ( .A(_144_), .Y(_145_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_146_) );
INVX1 INVX1_75 ( .A(_146_), .Y(_147_) );
NAND3X1 NAND3X1_29 ( .A(_145_), .B(_147_), .C(_140_), .Y(_148_) );
OAI21X1 OAI21X1_24 ( .A(_142_), .B(_143_), .C(_148_), .Y(w_C_27_) );
NOR2X1 NOR2X1_35 ( .A(_142_), .B(_143_), .Y(_149_) );
INVX1 INVX1_76 ( .A(_149_), .Y(_150_) );
AND2X2 AND2X2_21 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_151_) );
INVX1 INVX1_77 ( .A(_151_), .Y(_152_) );
NAND3X1 NAND3X1_30 ( .A(_150_), .B(_152_), .C(_148_), .Y(_153_) );
OAI21X1 OAI21X1_25 ( .A(i_add2[27]), .B(i_add1[27]), .C(_153_), .Y(_154_) );
INVX1 INVX1_78 ( .A(_154_), .Y(w_C_28_) );
INVX1 INVX1_79 ( .A(i_add2[28]), .Y(_155_) );
INVX1 INVX1_80 ( .A(i_add1[28]), .Y(_156_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_157_) );
INVX1 INVX1_81 ( .A(_157_), .Y(_158_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_159_) );
INVX1 INVX1_82 ( .A(_159_), .Y(_160_) );
NAND3X1 NAND3X1_31 ( .A(_158_), .B(_160_), .C(_153_), .Y(_161_) );
OAI21X1 OAI21X1_26 ( .A(_155_), .B(_156_), .C(_161_), .Y(w_C_29_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_162_) );
INVX1 INVX1_83 ( .A(_162_), .Y(_163_) );
NOR2X1 NOR2X1_39 ( .A(_155_), .B(_156_), .Y(_164_) );
INVX1 INVX1_84 ( .A(_164_), .Y(_165_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_166_) );
NAND3X1 NAND3X1_32 ( .A(_165_), .B(_166_), .C(_161_), .Y(_167_) );
AND2X2 AND2X2_22 ( .A(_167_), .B(_163_), .Y(w_C_30_) );
INVX1 INVX1_85 ( .A(i_add2[30]), .Y(_168_) );
INVX1 INVX1_86 ( .A(i_add1[30]), .Y(_169_) );
NAND2X1 NAND2X1_19 ( .A(_168_), .B(_169_), .Y(_170_) );
NAND3X1 NAND3X1_33 ( .A(_163_), .B(_170_), .C(_167_), .Y(_171_) );
OAI21X1 OAI21X1_27 ( .A(_168_), .B(_169_), .C(_171_), .Y(w_C_31_) );
INVX1 INVX1_87 ( .A(i_add2[31]), .Y(_172_) );
INVX1 INVX1_88 ( .A(i_add1[31]), .Y(_173_) );
NAND2X1 NAND2X1_20 ( .A(_172_), .B(_173_), .Y(_174_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_175_) );
NAND2X1 NAND2X1_22 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_176_) );
NAND3X1 NAND3X1_34 ( .A(_175_), .B(_176_), .C(_171_), .Y(_177_) );
AND2X2 AND2X2_23 ( .A(_177_), .B(_174_), .Y(w_C_32_) );
INVX1 INVX1_89 ( .A(i_add2[32]), .Y(_178_) );
INVX1 INVX1_90 ( .A(i_add1[32]), .Y(_179_) );
NAND2X1 NAND2X1_23 ( .A(_178_), .B(_179_), .Y(_180_) );
NAND3X1 NAND3X1_35 ( .A(_174_), .B(_180_), .C(_177_), .Y(_181_) );
OAI21X1 OAI21X1_28 ( .A(_178_), .B(_179_), .C(_181_), .Y(w_C_33_) );
NOR2X1 NOR2X1_40 ( .A(_178_), .B(_179_), .Y(_182_) );
INVX1 INVX1_91 ( .A(_182_), .Y(_183_) );
AND2X2 AND2X2_24 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_184_) );
INVX1 INVX1_92 ( .A(_184_), .Y(_185_) );
NAND3X1 NAND3X1_36 ( .A(_183_), .B(_185_), .C(_181_), .Y(_186_) );
OAI21X1 OAI21X1_29 ( .A(i_add2[33]), .B(i_add1[33]), .C(_186_), .Y(_187_) );
INVX1 INVX1_93 ( .A(_187_), .Y(w_C_34_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_188_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_189_) );
OAI21X1 OAI21X1_30 ( .A(_189_), .B(_187_), .C(_188_), .Y(w_C_35_) );
OR2X2 OR2X2_9 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_190_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_191_) );
INVX1 INVX1_94 ( .A(_191_), .Y(_192_) );
INVX1 INVX1_95 ( .A(_189_), .Y(_193_) );
NAND3X1 NAND3X1_37 ( .A(_192_), .B(_193_), .C(_186_), .Y(_194_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_195_) );
NAND3X1 NAND3X1_38 ( .A(_188_), .B(_195_), .C(_194_), .Y(_196_) );
AND2X2 AND2X2_25 ( .A(_196_), .B(_190_), .Y(w_C_36_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_197_) );
OR2X2 OR2X2_10 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_198_) );
NAND3X1 NAND3X1_39 ( .A(_190_), .B(_198_), .C(_196_), .Y(_199_) );
NAND2X1 NAND2X1_27 ( .A(_197_), .B(_199_), .Y(w_C_37_) );
BUFX2 BUFX2_1 ( .A(_200__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_200__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_200__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_200__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_200__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_200__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_200__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_200__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_200__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_200__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_200__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_200__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_200__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_200__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_200__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_200__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_200__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_200__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_200__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_200__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_200__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_200__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_200__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_200__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_200__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_200__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_200__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_200__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_200__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_200__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_200__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_200__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_200__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_200__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_200__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_200__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_200__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(w_C_37_), .Y(o_result[37]) );
INVX1 INVX1_96 ( .A(w_C_4_), .Y(_204_) );
OR2X2 OR2X2_11 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_205_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_206_) );
NAND3X1 NAND3X1_40 ( .A(_204_), .B(_206_), .C(_205_), .Y(_207_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_201_) );
AND2X2 AND2X2_26 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_202_) );
OAI21X1 OAI21X1_31 ( .A(_201_), .B(_202_), .C(w_C_4_), .Y(_203_) );
NAND2X1 NAND2X1_29 ( .A(_203_), .B(_207_), .Y(_200__4_) );
INVX1 INVX1_97 ( .A(w_C_5_), .Y(_211_) );
OR2X2 OR2X2_12 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_212_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_213_) );
NAND3X1 NAND3X1_41 ( .A(_211_), .B(_213_), .C(_212_), .Y(_214_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_208_) );
AND2X2 AND2X2_27 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_209_) );
OAI21X1 OAI21X1_32 ( .A(_208_), .B(_209_), .C(w_C_5_), .Y(_210_) );
NAND2X1 NAND2X1_31 ( .A(_210_), .B(_214_), .Y(_200__5_) );
INVX1 INVX1_98 ( .A(w_C_6_), .Y(_218_) );
OR2X2 OR2X2_13 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_219_) );
NAND2X1 NAND2X1_32 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_220_) );
NAND3X1 NAND3X1_42 ( .A(_218_), .B(_220_), .C(_219_), .Y(_221_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_215_) );
AND2X2 AND2X2_28 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_216_) );
OAI21X1 OAI21X1_33 ( .A(_215_), .B(_216_), .C(w_C_6_), .Y(_217_) );
NAND2X1 NAND2X1_33 ( .A(_217_), .B(_221_), .Y(_200__6_) );
INVX1 INVX1_99 ( .A(w_C_7_), .Y(_225_) );
OR2X2 OR2X2_14 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_226_) );
NAND2X1 NAND2X1_34 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_227_) );
NAND3X1 NAND3X1_43 ( .A(_225_), .B(_227_), .C(_226_), .Y(_228_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_222_) );
AND2X2 AND2X2_29 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_223_) );
OAI21X1 OAI21X1_34 ( .A(_222_), .B(_223_), .C(w_C_7_), .Y(_224_) );
NAND2X1 NAND2X1_35 ( .A(_224_), .B(_228_), .Y(_200__7_) );
INVX1 INVX1_100 ( .A(w_C_8_), .Y(_232_) );
OR2X2 OR2X2_15 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_233_) );
NAND2X1 NAND2X1_36 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_234_) );
NAND3X1 NAND3X1_44 ( .A(_232_), .B(_234_), .C(_233_), .Y(_235_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_229_) );
AND2X2 AND2X2_30 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_230_) );
OAI21X1 OAI21X1_35 ( .A(_229_), .B(_230_), .C(w_C_8_), .Y(_231_) );
NAND2X1 NAND2X1_37 ( .A(_231_), .B(_235_), .Y(_200__8_) );
INVX1 INVX1_101 ( .A(w_C_9_), .Y(_239_) );
OR2X2 OR2X2_16 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_240_) );
NAND2X1 NAND2X1_38 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_241_) );
NAND3X1 NAND3X1_45 ( .A(_239_), .B(_241_), .C(_240_), .Y(_242_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_236_) );
AND2X2 AND2X2_31 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_237_) );
OAI21X1 OAI21X1_36 ( .A(_236_), .B(_237_), .C(w_C_9_), .Y(_238_) );
NAND2X1 NAND2X1_39 ( .A(_238_), .B(_242_), .Y(_200__9_) );
INVX1 INVX1_102 ( .A(w_C_10_), .Y(_246_) );
OR2X2 OR2X2_17 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_247_) );
NAND2X1 NAND2X1_40 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_248_) );
NAND3X1 NAND3X1_46 ( .A(_246_), .B(_248_), .C(_247_), .Y(_249_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_243_) );
AND2X2 AND2X2_32 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_244_) );
OAI21X1 OAI21X1_37 ( .A(_243_), .B(_244_), .C(w_C_10_), .Y(_245_) );
NAND2X1 NAND2X1_41 ( .A(_245_), .B(_249_), .Y(_200__10_) );
INVX1 INVX1_103 ( .A(w_C_11_), .Y(_253_) );
OR2X2 OR2X2_18 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_254_) );
NAND2X1 NAND2X1_42 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_255_) );
NAND3X1 NAND3X1_47 ( .A(_253_), .B(_255_), .C(_254_), .Y(_256_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_250_) );
AND2X2 AND2X2_33 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_251_) );
OAI21X1 OAI21X1_38 ( .A(_250_), .B(_251_), .C(w_C_11_), .Y(_252_) );
NAND2X1 NAND2X1_43 ( .A(_252_), .B(_256_), .Y(_200__11_) );
INVX1 INVX1_104 ( .A(w_C_12_), .Y(_260_) );
OR2X2 OR2X2_19 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_261_) );
NAND2X1 NAND2X1_44 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_262_) );
NAND3X1 NAND3X1_48 ( .A(_260_), .B(_262_), .C(_261_), .Y(_263_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_257_) );
AND2X2 AND2X2_34 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_258_) );
OAI21X1 OAI21X1_39 ( .A(_257_), .B(_258_), .C(w_C_12_), .Y(_259_) );
NAND2X1 NAND2X1_45 ( .A(_259_), .B(_263_), .Y(_200__12_) );
INVX1 INVX1_105 ( .A(w_C_13_), .Y(_267_) );
OR2X2 OR2X2_20 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_268_) );
NAND2X1 NAND2X1_46 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_269_) );
NAND3X1 NAND3X1_49 ( .A(_267_), .B(_269_), .C(_268_), .Y(_270_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_264_) );
AND2X2 AND2X2_35 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_265_) );
OAI21X1 OAI21X1_40 ( .A(_264_), .B(_265_), .C(w_C_13_), .Y(_266_) );
NAND2X1 NAND2X1_47 ( .A(_266_), .B(_270_), .Y(_200__13_) );
INVX1 INVX1_106 ( .A(w_C_14_), .Y(_274_) );
OR2X2 OR2X2_21 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_275_) );
NAND2X1 NAND2X1_48 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_276_) );
NAND3X1 NAND3X1_50 ( .A(_274_), .B(_276_), .C(_275_), .Y(_277_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_271_) );
AND2X2 AND2X2_36 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_272_) );
OAI21X1 OAI21X1_41 ( .A(_271_), .B(_272_), .C(w_C_14_), .Y(_273_) );
NAND2X1 NAND2X1_49 ( .A(_273_), .B(_277_), .Y(_200__14_) );
INVX1 INVX1_107 ( .A(w_C_15_), .Y(_281_) );
OR2X2 OR2X2_22 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_282_) );
NAND2X1 NAND2X1_50 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_283_) );
NAND3X1 NAND3X1_51 ( .A(_281_), .B(_283_), .C(_282_), .Y(_284_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_278_) );
AND2X2 AND2X2_37 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_279_) );
OAI21X1 OAI21X1_42 ( .A(_278_), .B(_279_), .C(w_C_15_), .Y(_280_) );
NAND2X1 NAND2X1_51 ( .A(_280_), .B(_284_), .Y(_200__15_) );
INVX1 INVX1_108 ( .A(w_C_16_), .Y(_288_) );
OR2X2 OR2X2_23 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_289_) );
NAND2X1 NAND2X1_52 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_290_) );
NAND3X1 NAND3X1_52 ( .A(_288_), .B(_290_), .C(_289_), .Y(_291_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_285_) );
AND2X2 AND2X2_38 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_286_) );
OAI21X1 OAI21X1_43 ( .A(_285_), .B(_286_), .C(w_C_16_), .Y(_287_) );
NAND2X1 NAND2X1_53 ( .A(_287_), .B(_291_), .Y(_200__16_) );
INVX1 INVX1_109 ( .A(w_C_17_), .Y(_295_) );
OR2X2 OR2X2_24 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_296_) );
NAND2X1 NAND2X1_54 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_297_) );
NAND3X1 NAND3X1_53 ( .A(_295_), .B(_297_), .C(_296_), .Y(_298_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_292_) );
AND2X2 AND2X2_39 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_293_) );
OAI21X1 OAI21X1_44 ( .A(_292_), .B(_293_), .C(w_C_17_), .Y(_294_) );
NAND2X1 NAND2X1_55 ( .A(_294_), .B(_298_), .Y(_200__17_) );
INVX1 INVX1_110 ( .A(w_C_18_), .Y(_302_) );
OR2X2 OR2X2_25 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_303_) );
NAND2X1 NAND2X1_56 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_304_) );
NAND3X1 NAND3X1_54 ( .A(_302_), .B(_304_), .C(_303_), .Y(_305_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_299_) );
AND2X2 AND2X2_40 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_300_) );
OAI21X1 OAI21X1_45 ( .A(_299_), .B(_300_), .C(w_C_18_), .Y(_301_) );
NAND2X1 NAND2X1_57 ( .A(_301_), .B(_305_), .Y(_200__18_) );
INVX1 INVX1_111 ( .A(w_C_19_), .Y(_309_) );
OR2X2 OR2X2_26 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_310_) );
NAND2X1 NAND2X1_58 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_311_) );
NAND3X1 NAND3X1_55 ( .A(_309_), .B(_311_), .C(_310_), .Y(_312_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_306_) );
AND2X2 AND2X2_41 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_307_) );
OAI21X1 OAI21X1_46 ( .A(_306_), .B(_307_), .C(w_C_19_), .Y(_308_) );
NAND2X1 NAND2X1_59 ( .A(_308_), .B(_312_), .Y(_200__19_) );
INVX1 INVX1_112 ( .A(w_C_20_), .Y(_316_) );
OR2X2 OR2X2_27 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_317_) );
NAND2X1 NAND2X1_60 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_318_) );
NAND3X1 NAND3X1_56 ( .A(_316_), .B(_318_), .C(_317_), .Y(_319_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_313_) );
AND2X2 AND2X2_42 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_314_) );
OAI21X1 OAI21X1_47 ( .A(_313_), .B(_314_), .C(w_C_20_), .Y(_315_) );
NAND2X1 NAND2X1_61 ( .A(_315_), .B(_319_), .Y(_200__20_) );
INVX1 INVX1_113 ( .A(w_C_21_), .Y(_323_) );
OR2X2 OR2X2_28 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_324_) );
NAND2X1 NAND2X1_62 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_325_) );
NAND3X1 NAND3X1_57 ( .A(_323_), .B(_325_), .C(_324_), .Y(_326_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_320_) );
AND2X2 AND2X2_43 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_321_) );
OAI21X1 OAI21X1_48 ( .A(_320_), .B(_321_), .C(w_C_21_), .Y(_322_) );
NAND2X1 NAND2X1_63 ( .A(_322_), .B(_326_), .Y(_200__21_) );
INVX1 INVX1_114 ( .A(w_C_22_), .Y(_330_) );
OR2X2 OR2X2_29 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_331_) );
NAND2X1 NAND2X1_64 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_332_) );
NAND3X1 NAND3X1_58 ( .A(_330_), .B(_332_), .C(_331_), .Y(_333_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_327_) );
AND2X2 AND2X2_44 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_328_) );
OAI21X1 OAI21X1_49 ( .A(_327_), .B(_328_), .C(w_C_22_), .Y(_329_) );
NAND2X1 NAND2X1_65 ( .A(_329_), .B(_333_), .Y(_200__22_) );
INVX1 INVX1_115 ( .A(w_C_23_), .Y(_337_) );
OR2X2 OR2X2_30 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_338_) );
NAND2X1 NAND2X1_66 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_339_) );
NAND3X1 NAND3X1_59 ( .A(_337_), .B(_339_), .C(_338_), .Y(_340_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_334_) );
AND2X2 AND2X2_45 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_335_) );
OAI21X1 OAI21X1_50 ( .A(_334_), .B(_335_), .C(w_C_23_), .Y(_336_) );
NAND2X1 NAND2X1_67 ( .A(_336_), .B(_340_), .Y(_200__23_) );
INVX1 INVX1_116 ( .A(w_C_24_), .Y(_344_) );
OR2X2 OR2X2_31 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_345_) );
NAND2X1 NAND2X1_68 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_346_) );
NAND3X1 NAND3X1_60 ( .A(_344_), .B(_346_), .C(_345_), .Y(_347_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_341_) );
AND2X2 AND2X2_46 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_342_) );
OAI21X1 OAI21X1_51 ( .A(_341_), .B(_342_), .C(w_C_24_), .Y(_343_) );
NAND2X1 NAND2X1_69 ( .A(_343_), .B(_347_), .Y(_200__24_) );
INVX1 INVX1_117 ( .A(w_C_25_), .Y(_351_) );
OR2X2 OR2X2_32 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_352_) );
NAND2X1 NAND2X1_70 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_353_) );
NAND3X1 NAND3X1_61 ( .A(_351_), .B(_353_), .C(_352_), .Y(_354_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_348_) );
AND2X2 AND2X2_47 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_349_) );
OAI21X1 OAI21X1_52 ( .A(_348_), .B(_349_), .C(w_C_25_), .Y(_350_) );
NAND2X1 NAND2X1_71 ( .A(_350_), .B(_354_), .Y(_200__25_) );
INVX1 INVX1_118 ( .A(w_C_26_), .Y(_358_) );
OR2X2 OR2X2_33 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_359_) );
NAND2X1 NAND2X1_72 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_360_) );
NAND3X1 NAND3X1_62 ( .A(_358_), .B(_360_), .C(_359_), .Y(_361_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_355_) );
AND2X2 AND2X2_48 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_356_) );
OAI21X1 OAI21X1_53 ( .A(_355_), .B(_356_), .C(w_C_26_), .Y(_357_) );
NAND2X1 NAND2X1_73 ( .A(_357_), .B(_361_), .Y(_200__26_) );
INVX1 INVX1_119 ( .A(w_C_27_), .Y(_365_) );
OR2X2 OR2X2_34 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_366_) );
NAND2X1 NAND2X1_74 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_367_) );
NAND3X1 NAND3X1_63 ( .A(_365_), .B(_367_), .C(_366_), .Y(_368_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_362_) );
AND2X2 AND2X2_49 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_363_) );
OAI21X1 OAI21X1_54 ( .A(_362_), .B(_363_), .C(w_C_27_), .Y(_364_) );
NAND2X1 NAND2X1_75 ( .A(_364_), .B(_368_), .Y(_200__27_) );
INVX1 INVX1_120 ( .A(w_C_28_), .Y(_372_) );
OR2X2 OR2X2_35 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_373_) );
NAND2X1 NAND2X1_76 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_374_) );
NAND3X1 NAND3X1_64 ( .A(_372_), .B(_374_), .C(_373_), .Y(_375_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_369_) );
AND2X2 AND2X2_50 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_370_) );
OAI21X1 OAI21X1_55 ( .A(_369_), .B(_370_), .C(w_C_28_), .Y(_371_) );
NAND2X1 NAND2X1_77 ( .A(_371_), .B(_375_), .Y(_200__28_) );
INVX1 INVX1_121 ( .A(w_C_29_), .Y(_379_) );
OR2X2 OR2X2_36 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_380_) );
NAND2X1 NAND2X1_78 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_381_) );
NAND3X1 NAND3X1_65 ( .A(_379_), .B(_381_), .C(_380_), .Y(_382_) );
NOR2X1 NOR2X1_68 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_376_) );
AND2X2 AND2X2_51 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_377_) );
OAI21X1 OAI21X1_56 ( .A(_376_), .B(_377_), .C(w_C_29_), .Y(_378_) );
NAND2X1 NAND2X1_79 ( .A(_378_), .B(_382_), .Y(_200__29_) );
INVX1 INVX1_122 ( .A(w_C_30_), .Y(_386_) );
OR2X2 OR2X2_37 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_387_) );
NAND2X1 NAND2X1_80 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_388_) );
NAND3X1 NAND3X1_66 ( .A(_386_), .B(_388_), .C(_387_), .Y(_389_) );
NOR2X1 NOR2X1_69 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_383_) );
AND2X2 AND2X2_52 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_384_) );
OAI21X1 OAI21X1_57 ( .A(_383_), .B(_384_), .C(w_C_30_), .Y(_385_) );
NAND2X1 NAND2X1_81 ( .A(_385_), .B(_389_), .Y(_200__30_) );
INVX1 INVX1_123 ( .A(w_C_31_), .Y(_393_) );
OR2X2 OR2X2_38 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_394_) );
NAND2X1 NAND2X1_82 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_395_) );
NAND3X1 NAND3X1_67 ( .A(_393_), .B(_395_), .C(_394_), .Y(_396_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_390_) );
AND2X2 AND2X2_53 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_391_) );
OAI21X1 OAI21X1_58 ( .A(_390_), .B(_391_), .C(w_C_31_), .Y(_392_) );
NAND2X1 NAND2X1_83 ( .A(_392_), .B(_396_), .Y(_200__31_) );
INVX1 INVX1_124 ( .A(w_C_32_), .Y(_400_) );
OR2X2 OR2X2_39 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_401_) );
NAND2X1 NAND2X1_84 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_402_) );
NAND3X1 NAND3X1_68 ( .A(_400_), .B(_402_), .C(_401_), .Y(_403_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_397_) );
AND2X2 AND2X2_54 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_398_) );
OAI21X1 OAI21X1_59 ( .A(_397_), .B(_398_), .C(w_C_32_), .Y(_399_) );
NAND2X1 NAND2X1_85 ( .A(_399_), .B(_403_), .Y(_200__32_) );
INVX1 INVX1_125 ( .A(w_C_33_), .Y(_407_) );
OR2X2 OR2X2_40 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_408_) );
NAND2X1 NAND2X1_86 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_409_) );
NAND3X1 NAND3X1_69 ( .A(_407_), .B(_409_), .C(_408_), .Y(_410_) );
NOR2X1 NOR2X1_72 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_404_) );
AND2X2 AND2X2_55 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_405_) );
OAI21X1 OAI21X1_60 ( .A(_404_), .B(_405_), .C(w_C_33_), .Y(_406_) );
NAND2X1 NAND2X1_87 ( .A(_406_), .B(_410_), .Y(_200__33_) );
INVX1 INVX1_126 ( .A(w_C_34_), .Y(_414_) );
OR2X2 OR2X2_41 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_415_) );
NAND2X1 NAND2X1_88 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_416_) );
NAND3X1 NAND3X1_70 ( .A(_414_), .B(_416_), .C(_415_), .Y(_417_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_411_) );
AND2X2 AND2X2_56 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_412_) );
OAI21X1 OAI21X1_61 ( .A(_411_), .B(_412_), .C(w_C_34_), .Y(_413_) );
NAND2X1 NAND2X1_89 ( .A(_413_), .B(_417_), .Y(_200__34_) );
INVX1 INVX1_127 ( .A(w_C_35_), .Y(_421_) );
OR2X2 OR2X2_42 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_422_) );
NAND2X1 NAND2X1_90 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_423_) );
NAND3X1 NAND3X1_71 ( .A(_421_), .B(_423_), .C(_422_), .Y(_424_) );
NOR2X1 NOR2X1_74 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_418_) );
AND2X2 AND2X2_57 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_419_) );
OAI21X1 OAI21X1_62 ( .A(_418_), .B(_419_), .C(w_C_35_), .Y(_420_) );
NAND2X1 NAND2X1_91 ( .A(_420_), .B(_424_), .Y(_200__35_) );
INVX1 INVX1_128 ( .A(w_C_36_), .Y(_428_) );
OR2X2 OR2X2_43 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_429_) );
NAND2X1 NAND2X1_92 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_430_) );
NAND3X1 NAND3X1_72 ( .A(_428_), .B(_430_), .C(_429_), .Y(_431_) );
NOR2X1 NOR2X1_75 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_425_) );
AND2X2 AND2X2_58 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_426_) );
OAI21X1 OAI21X1_63 ( .A(_425_), .B(_426_), .C(w_C_36_), .Y(_427_) );
NAND2X1 NAND2X1_93 ( .A(_427_), .B(_431_), .Y(_200__36_) );
INVX1 INVX1_129 ( .A(1'b0), .Y(_435_) );
BUFX2 BUFX2_39 ( .A(w_C_37_), .Y(_200__37_) );
BUFX2 BUFX2_40 ( .A(1'b0), .Y(w_C_0_) );
endmodule
