module cla_60bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [59:0] i_add1;
input [59:0] i_add2;
output [60:0] o_result;

NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_261_), .C(_254_), .Y(_262_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_257_), .C(_262_), .Y(w_C_44_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_257_), .Y(_263_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_263_), .Y(_264_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_265_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_265_), .Y(_266_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_266_), .C(_262_), .Y(_267_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .C(_267_), .Y(_268_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_268_), .Y(w_C_45_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .Y(_269_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add1[45]), .Y(_270_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_271_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_271_), .Y(_272_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_273_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_273_), .Y(_274_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_274_), .C(_267_), .Y(_275_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_270_), .C(_275_), .Y(w_C_46_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_270_), .Y(_276_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_276_), .Y(_277_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_278_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_278_), .Y(_279_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_279_), .C(_275_), .Y(_280_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .C(_280_), .Y(_281_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_281_), .Y(w_C_47_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .Y(_282_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add1[47]), .Y(_283_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_284_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_284_), .Y(_285_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_286_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_286_), .Y(_287_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_287_), .C(_280_), .Y(_288_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_283_), .C(_288_), .Y(w_C_48_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_289_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_289_), .Y(_290_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_283_), .Y(_291_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_291_), .Y(_292_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_293_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_292_), .B(_293_), .C(_288_), .Y(_294_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_290_), .Y(w_C_49_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .Y(_295_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add1[49]), .Y(_296_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_296_), .Y(_297_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_297_), .C(_294_), .Y(_298_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_296_), .C(_298_), .Y(w_C_50_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .Y(_299_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add1[50]), .Y(_300_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .C(w_C_50_), .Y(_301_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_300_), .C(_301_), .Y(w_C_51_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .Y(_302_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add1[51]), .Y(_303_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_303_), .Y(_304_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(w_C_51_), .B(_304_), .Y(_305_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .C(_305_), .Y(_306_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_306_), .Y(w_C_52_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_307_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_308_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_306_), .C(_307_), .Y(w_C_53_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .Y(_309_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add1[53]), .Y(_310_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_308_), .Y(_311_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_304_), .Y(_312_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_300_), .Y(_313_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_314_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_315_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_315_), .C(_298_), .Y(_316_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_303_), .Y(_317_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_317_), .C(_316_), .Y(_318_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_307_), .C(_318_), .Y(_319_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_310_), .Y(_320_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_320_), .C(_319_), .Y(_321_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_310_), .C(_321_), .Y(w_C_54_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .Y(_322_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add1[54]), .Y(_323_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .C(w_C_54_), .Y(_324_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_323_), .C(_324_), .Y(w_C_55_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_323_), .Y(_325_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_325_), .Y(_326_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_327_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_327_), .Y(_328_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_328_), .C(_324_), .Y(_329_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .C(_329_), .Y(_330_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_330_), .Y(w_C_56_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_331_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_332_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_330_), .C(_331_), .Y(w_C_57_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_333_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_332_), .Y(_334_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_335_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_335_), .Y(_336_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_310_), .Y(_337_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_337_), .Y(_338_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_326_), .C(_321_), .Y(_339_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_340_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_340_), .Y(_341_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_341_), .C(_339_), .Y(_342_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_331_), .C(_342_), .Y(_343_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_344_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_344_), .C(_343_), .Y(_345_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_345_), .Y(w_C_58_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_346_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_347_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_347_), .C(_345_), .Y(_348_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_346_), .Y(w_C_59_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_349_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_350_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_350_), .C(_348_), .Y(_351_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_351_), .Y(w_C_60_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_2_), .Y(w_C_2_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .Y(_3_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add1[2]), .Y(_4_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_2_), .C(_6_), .Y(_7_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_9_), .C(_7_), .Y(_10_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_10_), .Y(w_C_4_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(_12_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_13_), .C(_10_), .Y(_14_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_12_), .Y(w_C_5_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .Y(_15_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add1[5]), .Y(_16_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_17_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_17_), .Y(_18_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_18_), .C(_14_), .Y(_19_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_16_), .C(_19_), .Y(w_C_6_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_20_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_20_), .Y(_21_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_16_), .Y(_22_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_23_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_24_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_24_), .Y(_25_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_25_), .C(_19_), .Y(_26_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_21_), .Y(w_C_7_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_27_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(_28_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_29_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_29_), .Y(_30_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_30_), .C(_26_), .Y(_31_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_28_), .Y(_32_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_32_), .Y(w_C_8_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_33_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_33_), .Y(_34_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_35_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_32_), .C(_34_), .Y(w_C_9_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_36_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_36_), .Y(_37_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_35_), .Y(_38_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_34_), .C(_31_), .Y(_39_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_40_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_40_), .Y(_41_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_41_), .C(_39_), .Y(_42_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_37_), .Y(_43_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(w_C_10_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_44_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_44_), .Y(_45_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_45_), .C(_42_), .Y(_46_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .C(_46_), .Y(_47_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_47_), .Y(w_C_11_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .Y(_48_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add1[11]), .Y(_49_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_50_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_50_), .Y(_51_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_52_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_52_), .Y(_53_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_53_), .C(_46_), .Y(_54_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_49_), .C(_54_), .Y(w_C_12_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_49_), .Y(_55_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_55_), .Y(_56_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_57_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_57_), .Y(_58_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_58_), .C(_54_), .Y(_59_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .C(_59_), .Y(_60_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_60_), .Y(w_C_13_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .Y(_61_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add1[13]), .Y(_62_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_63_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_63_), .Y(_64_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_352__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_352__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_352__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_352__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_352__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_352__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_352__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_352__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_352__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_352__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_352__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_352__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_352__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_352__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_352__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_352__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_352__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_352__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_352__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_352__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_352__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_352__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_352__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_352__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_352__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_352__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_352__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_352__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_352__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_352__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_352__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_352__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_352__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_352__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_352__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_352__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_352__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_352__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_352__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_352__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_352__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_352__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_352__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_352__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_352__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_352__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_352__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_352__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_352__48_), .Y(o_result[48]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_352__49_), .Y(o_result[49]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_352__50_), .Y(o_result[50]) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_352__51_), .Y(o_result[51]) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(_352__52_), .Y(o_result[52]) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(_352__53_), .Y(o_result[53]) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(_352__54_), .Y(o_result[54]) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_352__55_), .Y(o_result[55]) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_352__56_), .Y(o_result[56]) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_352__57_), .Y(o_result[57]) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_352__58_), .Y(o_result[58]) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(_352__59_), .Y(o_result[59]) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(w_C_60_), .Y(o_result[60]) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_356_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_357_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_358_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_358_), .C(_357_), .Y(_359_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_353_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_354_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_354_), .C(w_C_4_), .Y(_355_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_359_), .Y(_352__4_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_363_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_364_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_365_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_365_), .C(_364_), .Y(_366_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_360_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_361_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_361_), .C(w_C_5_), .Y(_362_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_366_), .Y(_352__5_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_370_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_371_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_372_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_372_), .C(_371_), .Y(_373_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_367_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_368_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_368_), .C(w_C_6_), .Y(_369_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_373_), .Y(_352__6_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_377_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_378_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_379_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_379_), .C(_378_), .Y(_380_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_374_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_375_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_375_), .C(w_C_7_), .Y(_376_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_380_), .Y(_352__7_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_384_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_385_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_386_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_386_), .C(_385_), .Y(_387_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_381_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_382_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_382_), .C(w_C_8_), .Y(_383_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_387_), .Y(_352__8_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_391_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_392_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_393_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_393_), .C(_392_), .Y(_394_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_388_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_389_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(_389_), .C(w_C_9_), .Y(_390_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_394_), .Y(_352__9_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_398_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_399_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_400_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_400_), .C(_399_), .Y(_401_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_395_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_396_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_396_), .C(w_C_10_), .Y(_397_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_401_), .Y(_352__10_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_405_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_406_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_407_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_407_), .C(_406_), .Y(_408_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_402_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_403_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_403_), .C(w_C_11_), .Y(_404_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_408_), .Y(_352__11_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(w_C_12_), .Y(_412_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_413_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_414_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_414_), .C(_413_), .Y(_415_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_409_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_410_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_410_), .C(w_C_12_), .Y(_411_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_415_), .Y(_352__12_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(w_C_13_), .Y(_419_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_420_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_421_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_421_), .C(_420_), .Y(_422_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_416_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_417_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_417_), .C(w_C_13_), .Y(_418_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_422_), .Y(_352__13_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(w_C_14_), .Y(_426_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_427_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_428_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_428_), .C(_427_), .Y(_429_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_423_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_424_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_424_), .C(w_C_14_), .Y(_425_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(_429_), .Y(_352__14_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(_433_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_434_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_435_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_435_), .C(_434_), .Y(_436_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_430_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_431_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_431_), .C(w_C_15_), .Y(_432_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_432_), .B(_436_), .Y(_352__15_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(w_C_16_), .Y(_440_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_441_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_442_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_442_), .C(_441_), .Y(_443_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_437_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_438_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_438_), .C(w_C_16_), .Y(_439_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_443_), .Y(_352__16_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(w_C_17_), .Y(_447_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_448_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_449_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_449_), .C(_448_), .Y(_450_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_444_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_445_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_445_), .C(w_C_17_), .Y(_446_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(_450_), .Y(_352__17_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(w_C_18_), .Y(_454_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_455_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_456_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_454_), .B(_456_), .C(_455_), .Y(_457_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_451_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_452_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_452_), .C(w_C_18_), .Y(_453_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(_457_), .Y(_352__18_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(w_C_19_), .Y(_461_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_462_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_463_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_463_), .C(_462_), .Y(_464_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_458_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_459_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_459_), .C(w_C_19_), .Y(_460_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_464_), .Y(_352__19_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(w_C_20_), .Y(_468_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_469_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_470_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_468_), .B(_470_), .C(_469_), .Y(_471_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_465_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_466_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_466_), .C(w_C_20_), .Y(_467_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_467_), .B(_471_), .Y(_352__20_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(w_C_21_), .Y(_475_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_476_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_477_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_477_), .C(_476_), .Y(_478_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_472_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_473_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_473_), .C(w_C_21_), .Y(_474_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_474_), .B(_478_), .Y(_352__21_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(w_C_22_), .Y(_482_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_483_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_484_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_482_), .B(_484_), .C(_483_), .Y(_485_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_479_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_480_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_480_), .C(w_C_22_), .Y(_481_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_485_), .Y(_352__22_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(w_C_23_), .Y(_489_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_490_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_491_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_491_), .C(_490_), .Y(_492_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_486_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_487_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_487_), .C(w_C_23_), .Y(_488_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_492_), .Y(_352__23_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(w_C_24_), .Y(_496_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_497_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_498_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_498_), .C(_497_), .Y(_499_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_493_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_494_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_494_), .C(w_C_24_), .Y(_495_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_495_), .B(_499_), .Y(_352__24_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(w_C_25_), .Y(_503_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_504_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_505_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_505_), .C(_504_), .Y(_506_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_500_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_501_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_501_), .C(w_C_25_), .Y(_502_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_502_), .B(_506_), .Y(_352__25_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(w_C_26_), .Y(_510_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_511_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_512_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_512_), .C(_511_), .Y(_513_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_507_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_508_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_508_), .C(w_C_26_), .Y(_509_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_513_), .Y(_352__26_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(w_C_27_), .Y(_517_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_518_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_519_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_517_), .B(_519_), .C(_518_), .Y(_520_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_514_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_515_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_515_), .C(w_C_27_), .Y(_516_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_520_), .Y(_352__27_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(w_C_28_), .Y(_524_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_525_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_526_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_526_), .C(_525_), .Y(_527_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_521_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_522_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_522_), .C(w_C_28_), .Y(_523_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_527_), .Y(_352__28_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(w_C_29_), .Y(_531_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_532_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_533_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_533_), .C(_532_), .Y(_534_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_528_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_529_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_529_), .C(w_C_29_), .Y(_530_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_534_), .Y(_352__29_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(w_C_30_), .Y(_538_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_539_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_540_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_540_), .C(_539_), .Y(_541_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_535_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_536_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_536_), .C(w_C_30_), .Y(_537_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_541_), .Y(_352__30_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(w_C_31_), .Y(_545_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_546_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_547_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_547_), .C(_546_), .Y(_548_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_542_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_543_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_542_), .B(_543_), .C(w_C_31_), .Y(_544_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_548_), .Y(_352__31_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(w_C_32_), .Y(_552_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_553_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_554_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_552_), .B(_554_), .C(_553_), .Y(_555_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_549_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_550_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(_550_), .C(w_C_32_), .Y(_551_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_551_), .B(_555_), .Y(_352__32_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(w_C_33_), .Y(_559_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_560_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_561_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_561_), .C(_560_), .Y(_562_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_556_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_557_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_556_), .B(_557_), .C(w_C_33_), .Y(_558_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_562_), .Y(_352__33_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(w_C_34_), .Y(_566_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_567_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_568_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_568_), .C(_567_), .Y(_569_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_563_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_564_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(_564_), .C(w_C_34_), .Y(_565_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_569_), .Y(_352__34_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(w_C_35_), .Y(_573_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_574_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_575_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_575_), .C(_574_), .Y(_576_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_570_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_571_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_571_), .C(w_C_35_), .Y(_572_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_576_), .Y(_352__35_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(w_C_36_), .Y(_580_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_581_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_582_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(_582_), .C(_581_), .Y(_583_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_577_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_578_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_578_), .C(w_C_36_), .Y(_579_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_583_), .Y(_352__36_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(w_C_37_), .Y(_587_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_588_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_589_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(_589_), .C(_588_), .Y(_590_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_584_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_585_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_585_), .C(w_C_37_), .Y(_586_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_586_), .B(_590_), .Y(_352__37_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(w_C_38_), .Y(_594_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_595_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_596_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_594_), .B(_596_), .C(_595_), .Y(_597_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_591_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_592_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_592_), .C(w_C_38_), .Y(_593_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_597_), .Y(_352__38_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(w_C_39_), .Y(_601_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_602_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_603_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_601_), .B(_603_), .C(_602_), .Y(_604_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_598_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_599_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_598_), .B(_599_), .C(w_C_39_), .Y(_600_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_604_), .Y(_352__39_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(w_C_40_), .Y(_608_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_609_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_610_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_608_), .B(_610_), .C(_609_), .Y(_611_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_605_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_606_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_606_), .C(w_C_40_), .Y(_607_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_611_), .Y(_352__40_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(w_C_41_), .Y(_615_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_616_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_617_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(_617_), .C(_616_), .Y(_618_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_612_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_613_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_612_), .B(_613_), .C(w_C_41_), .Y(_614_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_618_), .Y(_352__41_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(w_C_42_), .Y(_622_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_623_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_624_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_622_), .B(_624_), .C(_623_), .Y(_625_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_619_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_620_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_620_), .C(w_C_42_), .Y(_621_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_625_), .Y(_352__42_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(w_C_43_), .Y(_629_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_630_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_631_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_629_), .B(_631_), .C(_630_), .Y(_632_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_626_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_627_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_627_), .C(w_C_43_), .Y(_628_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_632_), .Y(_352__43_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(w_C_44_), .Y(_636_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_637_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_638_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_636_), .B(_638_), .C(_637_), .Y(_639_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_633_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_634_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_634_), .C(w_C_44_), .Y(_635_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_639_), .Y(_352__44_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(w_C_45_), .Y(_643_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_644_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_645_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_645_), .C(_644_), .Y(_646_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_640_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_641_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(_641_), .C(w_C_45_), .Y(_642_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_642_), .B(_646_), .Y(_352__45_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(w_C_46_), .Y(_650_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_651_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_652_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(_652_), .C(_651_), .Y(_653_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_647_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_648_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_647_), .B(_648_), .C(w_C_46_), .Y(_649_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_653_), .Y(_352__46_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(w_C_47_), .Y(_657_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_658_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_659_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_657_), .B(_659_), .C(_658_), .Y(_660_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_654_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_655_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_655_), .C(w_C_47_), .Y(_656_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_656_), .B(_660_), .Y(_352__47_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(w_C_48_), .Y(_664_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_665_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_666_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_666_), .C(_665_), .Y(_667_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_661_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_662_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_661_), .B(_662_), .C(w_C_48_), .Y(_663_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(_667_), .Y(_352__48_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(w_C_49_), .Y(_671_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_672_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_673_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_671_), .B(_673_), .C(_672_), .Y(_674_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_668_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_669_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_669_), .C(w_C_49_), .Y(_670_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(_674_), .Y(_352__49_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(w_C_50_), .Y(_678_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_679_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_680_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_680_), .C(_679_), .Y(_681_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_675_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_676_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_676_), .C(w_C_50_), .Y(_677_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_681_), .Y(_352__50_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(w_C_51_), .Y(_685_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_686_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_687_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_687_), .C(_686_), .Y(_688_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_682_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_683_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_682_), .B(_683_), .C(w_C_51_), .Y(_684_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_684_), .B(_688_), .Y(_352__51_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(w_C_52_), .Y(_692_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_693_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_694_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_692_), .B(_694_), .C(_693_), .Y(_695_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_689_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_690_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_690_), .C(w_C_52_), .Y(_691_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_691_), .B(_695_), .Y(_352__52_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(w_C_53_), .Y(_699_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_700_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_701_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_701_), .C(_700_), .Y(_702_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_696_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_697_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_697_), .C(w_C_53_), .Y(_698_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_702_), .Y(_352__53_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(w_C_54_), .Y(_706_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_707_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_708_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_708_), .C(_707_), .Y(_709_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_703_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_704_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_704_), .C(w_C_54_), .Y(_705_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_705_), .B(_709_), .Y(_352__54_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(w_C_55_), .Y(_713_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_714_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_715_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_715_), .C(_714_), .Y(_716_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_710_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_711_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_710_), .B(_711_), .C(w_C_55_), .Y(_712_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_712_), .B(_716_), .Y(_352__55_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(w_C_56_), .Y(_720_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_721_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_722_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_720_), .B(_722_), .C(_721_), .Y(_723_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_717_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_718_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_717_), .B(_718_), .C(w_C_56_), .Y(_719_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(_723_), .Y(_352__56_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(w_C_57_), .Y(_727_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_728_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_729_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_727_), .B(_729_), .C(_728_), .Y(_730_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_724_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_725_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_724_), .B(_725_), .C(w_C_57_), .Y(_726_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_726_), .B(_730_), .Y(_352__57_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(w_C_58_), .Y(_734_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_735_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_736_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_734_), .B(_736_), .C(_735_), .Y(_737_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_731_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_732_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_731_), .B(_732_), .C(w_C_58_), .Y(_733_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_733_), .B(_737_), .Y(_352__58_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(w_C_59_), .Y(_741_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_742_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_743_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_741_), .B(_743_), .C(_742_), .Y(_744_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_738_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_739_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_738_), .B(_739_), .C(w_C_59_), .Y(_740_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_740_), .B(_744_), .Y(_352__59_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_748_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_749_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_750_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_748_), .B(_750_), .C(_749_), .Y(_751_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_745_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_746_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_745_), .B(_746_), .C(gnd), .Y(_747_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_747_), .B(_751_), .Y(_352__0_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_755_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_756_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_757_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_757_), .C(_756_), .Y(_758_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_752_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_753_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(_753_), .C(w_C_1_), .Y(_754_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_754_), .B(_758_), .Y(_352__1_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_762_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_763_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_764_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_762_), .B(_764_), .C(_763_), .Y(_765_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_759_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_760_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_759_), .B(_760_), .C(w_C_2_), .Y(_761_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_761_), .B(_765_), .Y(_352__2_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_769_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_770_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_771_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_769_), .B(_771_), .C(_770_), .Y(_772_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_766_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_767_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_766_), .B(_767_), .C(w_C_3_), .Y(_768_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_768_), .B(_772_), .Y(_352__3_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_65_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(_65_), .Y(_66_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_66_), .C(_59_), .Y(_67_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_62_), .C(_67_), .Y(w_C_14_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_62_), .Y(_68_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(_68_), .Y(_69_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_70_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(_70_), .Y(_71_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_71_), .C(_67_), .Y(_72_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .C(_72_), .Y(_73_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(_73_), .Y(w_C_15_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .Y(_74_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(i_add1[15]), .Y(_75_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_76_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(_76_), .Y(_77_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_78_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(_78_), .Y(_79_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_79_), .C(_72_), .Y(_80_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_75_), .C(_80_), .Y(w_C_16_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_75_), .Y(_81_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(_81_), .Y(_82_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_83_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(_83_), .Y(_84_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_84_), .C(_80_), .Y(_85_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .C(_85_), .Y(_86_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(_86_), .Y(w_C_17_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .Y(_87_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(i_add1[17]), .Y(_88_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_89_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(_89_), .Y(_90_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_91_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(_91_), .Y(_92_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_92_), .C(_85_), .Y(_93_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_88_), .C(_93_), .Y(w_C_18_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_88_), .Y(_94_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(_94_), .Y(_95_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_96_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(_96_), .Y(_97_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_97_), .C(_93_), .Y(_98_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .C(_98_), .Y(_99_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(_99_), .Y(w_C_19_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .Y(_100_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(i_add1[19]), .Y(_101_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_102_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(_102_), .Y(_103_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_104_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(_104_), .Y(_105_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_105_), .C(_98_), .Y(_106_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_101_), .C(_106_), .Y(w_C_20_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_101_), .Y(_107_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(_107_), .Y(_108_) );
AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_109_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(_109_), .Y(_110_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_110_), .C(_106_), .Y(_111_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .C(_111_), .Y(_112_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(_112_), .Y(w_C_21_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .Y(_113_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(i_add1[21]), .Y(_114_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_115_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(_115_), .Y(_116_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_117_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(_117_), .Y(_118_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_118_), .C(_111_), .Y(_119_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_114_), .C(_119_), .Y(w_C_22_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_114_), .Y(_120_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(_120_), .Y(_121_) );
AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_122_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(_122_), .Y(_123_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_123_), .C(_119_), .Y(_124_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .C(_124_), .Y(_125_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(_125_), .Y(w_C_23_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .Y(_126_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(i_add1[23]), .Y(_127_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_128_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(_128_), .Y(_129_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_130_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(_130_), .Y(_131_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_129_), .B(_131_), .C(_124_), .Y(_132_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_127_), .C(_132_), .Y(w_C_24_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_127_), .Y(_133_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(_133_), .Y(_134_) );
AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_135_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(_135_), .Y(_136_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_136_), .C(_132_), .Y(_137_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .C(_137_), .Y(_138_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(_138_), .Y(w_C_25_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .Y(_139_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(i_add1[25]), .Y(_140_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_141_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(_141_), .Y(_142_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_143_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(_143_), .Y(_144_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_144_), .C(_137_), .Y(_145_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_140_), .C(_145_), .Y(w_C_26_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_140_), .Y(_146_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(_146_), .Y(_147_) );
AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_148_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(_148_), .Y(_149_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_149_), .C(_145_), .Y(_150_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .C(_150_), .Y(_151_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(_151_), .Y(w_C_27_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .Y(_152_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(i_add1[27]), .Y(_153_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_154_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(_154_), .Y(_155_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_156_) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_157_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_157_), .C(_150_), .Y(_158_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_153_), .C(_158_), .Y(w_C_28_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_153_), .Y(_159_) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(_159_), .Y(_160_) );
AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_161_) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(_161_), .Y(_162_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_162_), .C(_158_), .Y(_163_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .C(_163_), .Y(_164_) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(_164_), .Y(w_C_29_) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .Y(_165_) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(i_add1[29]), .Y(_166_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_167_) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(_167_), .Y(_168_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_169_) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(_169_), .Y(_170_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_170_), .C(_163_), .Y(_171_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_166_), .C(_171_), .Y(w_C_30_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_166_), .Y(_172_) );
INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(_172_), .Y(_173_) );
AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_174_) );
INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(_174_), .Y(_175_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(_175_), .C(_171_), .Y(_176_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .C(_176_), .Y(_177_) );
INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(_177_), .Y(w_C_31_) );
INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .Y(_178_) );
INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(i_add1[31]), .Y(_179_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_180_) );
INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(_180_), .Y(_181_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_182_) );
INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(_182_), .Y(_183_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_183_), .C(_176_), .Y(_184_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_179_), .C(_184_), .Y(w_C_32_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_179_), .Y(_185_) );
INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(_185_), .Y(_186_) );
AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_187_) );
INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(_187_), .Y(_188_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_188_), .C(_184_), .Y(_189_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .C(_189_), .Y(_190_) );
INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(_190_), .Y(w_C_33_) );
INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .Y(_191_) );
INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(i_add1[33]), .Y(_192_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_193_) );
INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(_193_), .Y(_194_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_195_) );
INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(_195_), .Y(_196_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_196_), .C(_189_), .Y(_197_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_192_), .C(_197_), .Y(w_C_34_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_192_), .Y(_198_) );
INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(_198_), .Y(_199_) );
AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_200_) );
INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(_200_), .Y(_201_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_201_), .C(_197_), .Y(_202_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .C(_202_), .Y(_203_) );
INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(_203_), .Y(w_C_35_) );
INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .Y(_204_) );
INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(i_add1[35]), .Y(_205_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_206_) );
INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(_206_), .Y(_207_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_208_) );
INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(_208_), .Y(_209_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_209_), .C(_202_), .Y(_210_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_205_), .C(_210_), .Y(w_C_36_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_205_), .Y(_211_) );
INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(_211_), .Y(_212_) );
AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_213_) );
INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(_213_), .Y(_214_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_214_), .C(_210_), .Y(_215_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .C(_215_), .Y(_216_) );
INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(_216_), .Y(w_C_37_) );
INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .Y(_217_) );
INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(i_add1[37]), .Y(_218_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_219_) );
INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(_219_), .Y(_220_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_221_) );
INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(_221_), .Y(_222_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_222_), .C(_215_), .Y(_223_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_218_), .C(_223_), .Y(w_C_38_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_218_), .Y(_224_) );
INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(_224_), .Y(_225_) );
AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_226_) );
INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(_226_), .Y(_227_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_227_), .C(_223_), .Y(_228_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .C(_228_), .Y(_229_) );
INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(_229_), .Y(w_C_39_) );
INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .Y(_230_) );
INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(i_add1[39]), .Y(_231_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_232_) );
INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(_232_), .Y(_233_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_234_) );
INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(_234_), .Y(_235_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_235_), .C(_228_), .Y(_236_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_231_), .C(_236_), .Y(w_C_40_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_231_), .Y(_237_) );
INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(_237_), .Y(_238_) );
AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_239_) );
INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(_239_), .Y(_240_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_238_), .B(_240_), .C(_236_), .Y(_241_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .C(_241_), .Y(_242_) );
INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(_242_), .Y(w_C_41_) );
INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .Y(_243_) );
INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(i_add1[41]), .Y(_244_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_245_) );
INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(_245_), .Y(_246_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_247_) );
INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(_247_), .Y(_248_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_248_), .C(_241_), .Y(_249_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_244_), .C(_249_), .Y(w_C_42_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_244_), .Y(_250_) );
INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(_250_), .Y(_251_) );
AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_252_) );
INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(_252_), .Y(_253_) );
NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_253_), .C(_249_), .Y(_254_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .C(_254_), .Y(_255_) );
INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(_255_), .Y(w_C_43_) );
INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .Y(_256_) );
INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(i_add1[43]), .Y(_257_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_258_) );
INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(_258_), .Y(_259_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_260_) );
INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(_260_), .Y(_261_) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(w_C_60_), .Y(_352__60_) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
