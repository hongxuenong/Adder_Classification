module CSkipA_35bit ( gnd, vdd, i_add_term1, i_add_term2, sum, cout);

input gnd, vdd;
output cout;
input [34:0] i_add_term1;
input [34:0] i_add_term2;
output [34:0] sum;

BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .Y(cout) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_0__34_), .Y(sum[34]) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .Y(_25_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(_25_), .Y(_26_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .Y(_27_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .B(_27_), .Y(_28_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .Y(_29_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(_29_), .Y(_30_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .Y(_31_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .B(_31_), .Y(_32_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_28_), .C(_30_), .D(_32_), .Y(_33_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_34_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_35_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_35_), .Y(_36_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_37_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_37_), .Y(_38_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_38_), .Y(_3_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_39_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_3_), .Y(_40_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_39_), .C(_40_), .Y(w_cout_1_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[4]), .Y(_41_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(_41_), .Y(_42_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .Y(_43_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[4]), .B(_43_), .Y(_44_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[5]), .Y(_45_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(_45_), .Y(_46_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .Y(_47_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[5]), .B(_47_), .Y(_48_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_44_), .C(_46_), .D(_48_), .Y(_49_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_50_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_51_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_51_), .Y(_52_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_53_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_53_), .Y(_54_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_54_), .Y(_6_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(_55_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_6_), .Y(_56_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_55_), .C(_56_), .Y(w_cout_2_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[8]), .Y(_57_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(_57_), .Y(_58_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .Y(_59_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[8]), .B(_59_), .Y(_60_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[9]), .Y(_61_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(_61_), .Y(_62_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .Y(_63_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[9]), .B(_63_), .Y(_64_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_60_), .C(_62_), .D(_64_), .Y(_65_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_66_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_67_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_67_), .Y(_68_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_69_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_69_), .Y(_70_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_70_), .Y(_9_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_71_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_9_), .Y(_72_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_71_), .C(_72_), .Y(w_cout_3_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[12]), .Y(_73_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(_73_), .Y(_74_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .Y(_75_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[12]), .B(_75_), .Y(_76_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[13]), .Y(_77_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(_77_), .Y(_78_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .Y(_79_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[13]), .B(_79_), .Y(_80_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_76_), .C(_78_), .D(_80_), .Y(_81_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_82_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_83_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_83_), .Y(_84_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_85_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_85_), .Y(_86_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_86_), .Y(_12_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(_87_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_12_), .Y(_88_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_87_), .C(_88_), .Y(w_cout_4_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[16]), .Y(_89_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(_89_), .Y(_90_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .Y(_91_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[16]), .B(_91_), .Y(_92_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[17]), .Y(_93_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(_93_), .Y(_94_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .Y(_95_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[17]), .B(_95_), .Y(_96_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_92_), .C(_94_), .D(_96_), .Y(_97_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_98_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_99_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_99_), .Y(_100_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_101_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_101_), .Y(_102_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_102_), .Y(_15_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_103_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_15_), .Y(_104_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_103_), .C(_104_), .Y(w_cout_5_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[20]), .Y(_105_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(_105_), .Y(_106_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .Y(_107_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[20]), .B(_107_), .Y(_108_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[21]), .Y(_109_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(_109_), .Y(_110_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .Y(_111_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[21]), .B(_111_), .Y(_112_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_106_), .B(_108_), .C(_110_), .D(_112_), .Y(_113_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_114_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_115_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_115_), .Y(_116_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_117_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_117_), .Y(_118_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_118_), .Y(_18_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_119_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_18_), .Y(_120_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_119_), .C(_120_), .Y(w_cout_6_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[24]), .Y(_121_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(_121_), .Y(_122_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .Y(_123_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[24]), .B(_123_), .Y(_124_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[25]), .Y(_125_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(_125_), .Y(_126_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .Y(_127_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[25]), .B(_127_), .Y(_128_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_124_), .C(_126_), .D(_128_), .Y(_129_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_130_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_131_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_131_), .Y(_132_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_133_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_133_), .Y(_134_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_129_), .B(_134_), .Y(_21_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_135_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_21_), .Y(_136_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_135_), .C(_136_), .Y(w_cout_7_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[28]), .Y(_137_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(_137_), .Y(_138_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .Y(_139_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[28]), .B(_139_), .Y(_140_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[29]), .Y(_141_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(_141_), .Y(_142_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .Y(_143_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[29]), .B(_143_), .Y(_144_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_140_), .C(_142_), .D(_144_), .Y(_145_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_146_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_147_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_147_), .Y(_148_) );
XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_149_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_149_), .Y(_150_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_150_), .Y(_24_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_151_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_24_), .Y(_152_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_151_), .C(_152_), .Y(cskip3_inst_cin) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_156_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_157_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_158_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_158_), .C(_157_), .Y(_159_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_153_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_154_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_154_), .C(gnd), .Y(_155_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_159_), .Y(_0__0_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_153_), .C(_158_), .Y(_2__1_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_2__1_), .Y(_163_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_164_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_165_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_165_), .C(_164_), .Y(_166_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_160_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_161_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_161_), .C(_2__1_), .Y(_162_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_166_), .Y(_0__1_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_160_), .C(_165_), .Y(_2__2_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_2__2_), .Y(_170_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_171_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_172_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_172_), .C(_171_), .Y(_173_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_167_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_168_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_168_), .C(_2__2_), .Y(_169_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_173_), .Y(_0__2_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_167_), .C(_172_), .Y(_2__3_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_2__3_), .Y(_177_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_178_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_179_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_179_), .C(_178_), .Y(_180_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_174_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_175_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_175_), .C(_2__3_), .Y(_176_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_180_), .Y(_0__3_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_174_), .C(_179_), .Y(_1_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .Y(_184_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_185_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_186_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_186_), .C(_185_), .Y(_187_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_181_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_182_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_182_), .C(w_cout_1_), .Y(_183_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_187_), .Y(_0__4_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_181_), .C(_186_), .Y(_5__1_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_5__1_), .Y(_191_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_192_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_193_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_193_), .C(_192_), .Y(_194_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_188_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_189_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_189_), .C(_5__1_), .Y(_190_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_194_), .Y(_0__5_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_188_), .C(_193_), .Y(_5__2_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_5__2_), .Y(_198_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_199_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_200_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_200_), .C(_199_), .Y(_201_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_195_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_196_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_196_), .C(_5__2_), .Y(_197_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_201_), .Y(_0__6_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_195_), .C(_200_), .Y(_5__3_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_5__3_), .Y(_205_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_206_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_207_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_207_), .C(_206_), .Y(_208_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_202_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_203_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_203_), .C(_5__3_), .Y(_204_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_208_), .Y(_0__7_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_202_), .C(_207_), .Y(_4_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .Y(_212_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_213_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_214_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_214_), .C(_213_), .Y(_215_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_209_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_210_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_210_), .C(w_cout_2_), .Y(_211_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_215_), .Y(_0__8_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_209_), .C(_214_), .Y(_8__1_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_8__1_), .Y(_219_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_220_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_221_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_221_), .C(_220_), .Y(_222_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_216_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_217_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_217_), .C(_8__1_), .Y(_218_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(_222_), .Y(_0__9_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_216_), .C(_221_), .Y(_8__2_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_8__2_), .Y(_226_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_227_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_228_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_228_), .C(_227_), .Y(_229_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_223_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_224_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_224_), .C(_8__2_), .Y(_225_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_229_), .Y(_0__10_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_223_), .C(_228_), .Y(_8__3_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_8__3_), .Y(_233_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_234_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_235_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_235_), .C(_234_), .Y(_236_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_230_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_231_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_231_), .C(_8__3_), .Y(_232_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_236_), .Y(_0__11_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_230_), .C(_235_), .Y(_7_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .Y(_240_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_241_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_242_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_242_), .C(_241_), .Y(_243_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_237_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_238_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_238_), .C(w_cout_3_), .Y(_239_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_243_), .Y(_0__12_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_237_), .C(_242_), .Y(_11__1_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_11__1_), .Y(_247_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_248_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_249_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_249_), .C(_248_), .Y(_250_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_244_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_245_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_245_), .C(_11__1_), .Y(_246_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_250_), .Y(_0__13_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_244_), .C(_249_), .Y(_11__2_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_11__2_), .Y(_254_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_255_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_256_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_256_), .C(_255_), .Y(_257_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_251_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_252_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_252_), .C(_11__2_), .Y(_253_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_253_), .B(_257_), .Y(_0__14_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_251_), .C(_256_), .Y(_11__3_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_11__3_), .Y(_261_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_262_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_263_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_263_), .C(_262_), .Y(_264_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_258_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_259_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_259_), .C(_11__3_), .Y(_260_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_264_), .Y(_0__15_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_258_), .C(_263_), .Y(_10_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .Y(_268_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_269_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_270_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_270_), .C(_269_), .Y(_271_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_265_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_266_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_266_), .C(w_cout_4_), .Y(_267_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_271_), .Y(_0__16_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_265_), .C(_270_), .Y(_14__1_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_14__1_), .Y(_275_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_276_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_277_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_277_), .C(_276_), .Y(_278_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_272_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_273_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_273_), .C(_14__1_), .Y(_274_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_278_), .Y(_0__17_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_272_), .C(_277_), .Y(_14__2_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_14__2_), .Y(_282_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_283_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_284_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_284_), .C(_283_), .Y(_285_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_279_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_280_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_279_), .B(_280_), .C(_14__2_), .Y(_281_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_285_), .Y(_0__18_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_279_), .C(_284_), .Y(_14__3_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_14__3_), .Y(_289_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_290_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_291_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_291_), .C(_290_), .Y(_292_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_286_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_287_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_287_), .C(_14__3_), .Y(_288_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_292_), .Y(_0__19_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_286_), .C(_291_), .Y(_13_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .Y(_296_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_297_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_298_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_298_), .C(_297_), .Y(_299_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_293_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_294_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_294_), .C(w_cout_5_), .Y(_295_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_299_), .Y(_0__20_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_293_), .C(_298_), .Y(_17__1_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_17__1_), .Y(_303_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_304_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_305_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_305_), .C(_304_), .Y(_306_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_300_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_301_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_301_), .C(_17__1_), .Y(_302_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_306_), .Y(_0__21_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_300_), .C(_305_), .Y(_17__2_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_17__2_), .Y(_310_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_311_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_312_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_312_), .C(_311_), .Y(_313_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_307_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_308_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_308_), .C(_17__2_), .Y(_309_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_313_), .Y(_0__22_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_307_), .C(_312_), .Y(_17__3_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_17__3_), .Y(_317_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_318_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_319_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_319_), .C(_318_), .Y(_320_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_314_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_315_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_315_), .C(_17__3_), .Y(_316_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_316_), .B(_320_), .Y(_0__23_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_314_), .C(_319_), .Y(_16_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .Y(_324_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_325_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_326_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_326_), .C(_325_), .Y(_327_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_321_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_322_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_322_), .C(w_cout_6_), .Y(_323_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_327_), .Y(_0__24_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_321_), .C(_326_), .Y(_20__1_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_20__1_), .Y(_331_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_332_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_333_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_333_), .C(_332_), .Y(_334_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_328_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_329_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_329_), .C(_20__1_), .Y(_330_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_334_), .Y(_0__25_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_328_), .C(_333_), .Y(_20__2_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_20__2_), .Y(_338_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_339_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_340_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_340_), .C(_339_), .Y(_341_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_335_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_336_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_335_), .B(_336_), .C(_20__2_), .Y(_337_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_341_), .Y(_0__26_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_335_), .C(_340_), .Y(_20__3_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_20__3_), .Y(_345_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_346_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_347_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_347_), .C(_346_), .Y(_348_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_342_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_343_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_343_), .C(_20__3_), .Y(_344_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_348_), .Y(_0__27_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_342_), .C(_347_), .Y(_19_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .Y(_352_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_353_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_354_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_354_), .C(_353_), .Y(_355_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_349_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_350_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_350_), .C(w_cout_7_), .Y(_351_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_355_), .Y(_0__28_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_349_), .C(_354_), .Y(_23__1_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_23__1_), .Y(_359_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_360_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_361_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_361_), .C(_360_), .Y(_362_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_356_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_357_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_357_), .C(_23__1_), .Y(_358_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_358_), .B(_362_), .Y(_0__29_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_356_), .C(_361_), .Y(_23__2_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(_23__2_), .Y(_366_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_367_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_368_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_368_), .C(_367_), .Y(_369_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_363_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_364_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_364_), .C(_23__2_), .Y(_365_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_365_), .B(_369_), .Y(_0__30_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_363_), .C(_368_), .Y(_23__3_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_23__3_), .Y(_373_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_374_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_375_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_373_), .B(_375_), .C(_374_), .Y(_376_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_370_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_371_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_371_), .C(_23__3_), .Y(_372_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_376_), .Y(_0__31_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_373_), .B(_370_), .C(_375_), .Y(_22_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_cin), .Y(_380_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_381_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_382_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_382_), .C(_381_), .Y(_383_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_377_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_378_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_378_), .C(cskip3_inst_cin), .Y(_379_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_383_), .Y(_0__32_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_377_), .C(_382_), .Y(cskip3_inst_rca0_w_CARRY_1_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_rca0_w_CARRY_1_), .Y(_387_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_388_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_389_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_389_), .C(_388_), .Y(_390_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_384_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_385_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_385_), .C(cskip3_inst_rca0_w_CARRY_1_), .Y(_386_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_390_), .Y(_0__33_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_384_), .C(_389_), .Y(cskip3_inst_rca0_w_CARRY_2_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_rca0_w_CARRY_2_), .Y(_394_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_395_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_396_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_396_), .C(_395_), .Y(_397_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_391_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_392_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_392_), .C(cskip3_inst_rca0_w_CARRY_2_), .Y(_393_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_397_), .Y(_0__34_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_391_), .C(_396_), .Y(cskip3_inst_rca0_w_CARRY_3_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_rca0_w_CARRY_3_), .Y(_399_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_400_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_398_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_398_), .C(_400_), .Y(cskip3_inst_cout0) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_404_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_405_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_404_), .Y(_401_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_402_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_403_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_402_), .C(_403_), .Y(cskip3_inst_skip0_P) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_cout0), .Y(_406_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(cskip3_inst_skip0_P), .Y(_407_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_skip0_P), .B(_406_), .C(_407_), .Y(w_cout_9_) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_2__0_) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .Y(_5__0_) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(_5__4_) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .Y(_8__0_) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .Y(_11__0_) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(_11__4_) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .Y(_14__0_) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .Y(_17__0_) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_17__4_) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .Y(_20__0_) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_20__4_) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .Y(_23__0_) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_23__4_) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_cin), .Y(cskip3_inst_rca0_w_CARRY_0_) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_cout0), .Y(cskip3_inst_rca0_w_CARRY_4_) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_cin), .Y(w_cout_8_) );
endmodule
