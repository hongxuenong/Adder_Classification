module cla_47bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add1[19], i_add1[20], i_add1[21], i_add1[22], i_add1[23], i_add1[24], i_add1[25], i_add1[26], i_add1[27], i_add1[28], i_add1[29], i_add1[30], i_add1[31], i_add1[32], i_add1[33], i_add1[34], i_add1[35], i_add1[36], i_add1[37], i_add1[38], i_add1[39], i_add1[40], i_add1[41], i_add1[42], i_add1[43], i_add1[44], i_add1[45], i_add1[46], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], i_add2[19], i_add2[20], i_add2[21], i_add2[22], i_add2[23], i_add2[24], i_add2[25], i_add2[26], i_add2[27], i_add2[28], i_add2[29], i_add2[30], i_add2[31], i_add2[32], i_add2[33], i_add2[34], i_add2[35], i_add2[36], i_add2[37], i_add2[38], i_add2[39], i_add2[40], i_add2[41], i_add2[42], i_add2[43], i_add2[44], i_add2[45], i_add2[46], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21], o_result[22], o_result[23], o_result[24], o_result[25], o_result[26], o_result[27], o_result[28], o_result[29], o_result[30], o_result[31], o_result[32], o_result[33], o_result[34], o_result[35], o_result[36], o_result[37], o_result[38], o_result[39], o_result[40], o_result[41], o_result[42], o_result[43], o_result[44], o_result[45], o_result[46], o_result[47]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add1[19];
input i_add1[20];
input i_add1[21];
input i_add1[22];
input i_add1[23];
input i_add1[24];
input i_add1[25];
input i_add1[26];
input i_add1[27];
input i_add1[28];
input i_add1[29];
input i_add1[30];
input i_add1[31];
input i_add1[32];
input i_add1[33];
input i_add1[34];
input i_add1[35];
input i_add1[36];
input i_add1[37];
input i_add1[38];
input i_add1[39];
input i_add1[40];
input i_add1[41];
input i_add1[42];
input i_add1[43];
input i_add1[44];
input i_add1[45];
input i_add1[46];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
input i_add2[19];
input i_add2[20];
input i_add2[21];
input i_add2[22];
input i_add2[23];
input i_add2[24];
input i_add2[25];
input i_add2[26];
input i_add2[27];
input i_add2[28];
input i_add2[29];
input i_add2[30];
input i_add2[31];
input i_add2[32];
input i_add2[33];
input i_add2[34];
input i_add2[35];
input i_add2[36];
input i_add2[37];
input i_add2[38];
input i_add2[39];
input i_add2[40];
input i_add2[41];
input i_add2[42];
input i_add2[43];
input i_add2[44];
input i_add2[45];
input i_add2[46];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];
output o_result[22];
output o_result[23];
output o_result[24];
output o_result[25];
output o_result[26];
output o_result[27];
output o_result[28];
output o_result[29];
output o_result[30];
output o_result[31];
output o_result[32];
output o_result[33];
output o_result[34];
output o_result[35];
output o_result[36];
output o_result[37];
output o_result[38];
output o_result[39];
output o_result[40];
output o_result[41];
output o_result[42];
output o_result[43];
output o_result[44];
output o_result[45];
output o_result[46];
output o_result[47];

NAND3X1 NAND3X1_1 ( .A(_296_), .B(_298_), .C(_297_), .Y(_299_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_293_) );
AND2X2 AND2X2_1 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_294_) );
OAI21X1 OAI21X1_1 ( .A(_293_), .B(_294_), .C(w_C_6_), .Y(_295_) );
NAND2X1 NAND2X1_1 ( .A(_295_), .B(_299_), .Y(_278__6_) );
INVX1 INVX1_1 ( .A(w_C_7_), .Y(_303_) );
OR2X2 OR2X2_1 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_304_) );
NAND2X1 NAND2X1_2 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_305_) );
NAND3X1 NAND3X1_2 ( .A(_303_), .B(_305_), .C(_304_), .Y(_306_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_300_) );
AND2X2 AND2X2_2 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_301_) );
OAI21X1 OAI21X1_2 ( .A(_300_), .B(_301_), .C(w_C_7_), .Y(_302_) );
NAND2X1 NAND2X1_3 ( .A(_302_), .B(_306_), .Y(_278__7_) );
INVX1 INVX1_2 ( .A(w_C_8_), .Y(_310_) );
OR2X2 OR2X2_2 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_311_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_312_) );
NAND3X1 NAND3X1_3 ( .A(_310_), .B(_312_), .C(_311_), .Y(_313_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_307_) );
AND2X2 AND2X2_3 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_308_) );
OAI21X1 OAI21X1_3 ( .A(_307_), .B(_308_), .C(w_C_8_), .Y(_309_) );
NAND2X1 NAND2X1_5 ( .A(_309_), .B(_313_), .Y(_278__8_) );
INVX1 INVX1_3 ( .A(w_C_9_), .Y(_317_) );
OR2X2 OR2X2_3 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_318_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_319_) );
NAND3X1 NAND3X1_4 ( .A(_317_), .B(_319_), .C(_318_), .Y(_320_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_314_) );
AND2X2 AND2X2_4 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_315_) );
OAI21X1 OAI21X1_4 ( .A(_314_), .B(_315_), .C(w_C_9_), .Y(_316_) );
NAND2X1 NAND2X1_7 ( .A(_316_), .B(_320_), .Y(_278__9_) );
INVX1 INVX1_4 ( .A(w_C_10_), .Y(_324_) );
OR2X2 OR2X2_4 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_325_) );
NAND2X1 NAND2X1_8 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_326_) );
NAND3X1 NAND3X1_5 ( .A(_324_), .B(_326_), .C(_325_), .Y(_327_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_321_) );
AND2X2 AND2X2_5 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_322_) );
OAI21X1 OAI21X1_5 ( .A(_321_), .B(_322_), .C(w_C_10_), .Y(_323_) );
NAND2X1 NAND2X1_9 ( .A(_323_), .B(_327_), .Y(_278__10_) );
INVX1 INVX1_5 ( .A(w_C_11_), .Y(_331_) );
OR2X2 OR2X2_5 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_332_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_333_) );
NAND3X1 NAND3X1_6 ( .A(_331_), .B(_333_), .C(_332_), .Y(_334_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_328_) );
AND2X2 AND2X2_6 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_329_) );
OAI21X1 OAI21X1_6 ( .A(_328_), .B(_329_), .C(w_C_11_), .Y(_330_) );
NAND2X1 NAND2X1_11 ( .A(_330_), .B(_334_), .Y(_278__11_) );
INVX1 INVX1_6 ( .A(w_C_12_), .Y(_338_) );
OR2X2 OR2X2_6 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_339_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_340_) );
NAND3X1 NAND3X1_7 ( .A(_338_), .B(_340_), .C(_339_), .Y(_341_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_335_) );
AND2X2 AND2X2_7 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_336_) );
OAI21X1 OAI21X1_7 ( .A(_335_), .B(_336_), .C(w_C_12_), .Y(_337_) );
NAND2X1 NAND2X1_13 ( .A(_337_), .B(_341_), .Y(_278__12_) );
INVX1 INVX1_7 ( .A(w_C_13_), .Y(_345_) );
OR2X2 OR2X2_7 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_346_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_347_) );
NAND3X1 NAND3X1_8 ( .A(_345_), .B(_347_), .C(_346_), .Y(_348_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_342_) );
AND2X2 AND2X2_8 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_343_) );
OAI21X1 OAI21X1_8 ( .A(_342_), .B(_343_), .C(w_C_13_), .Y(_344_) );
NAND2X1 NAND2X1_15 ( .A(_344_), .B(_348_), .Y(_278__13_) );
INVX1 INVX1_8 ( .A(w_C_14_), .Y(_352_) );
OR2X2 OR2X2_8 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_353_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_354_) );
NAND3X1 NAND3X1_9 ( .A(_352_), .B(_354_), .C(_353_), .Y(_355_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_349_) );
AND2X2 AND2X2_9 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_350_) );
OAI21X1 OAI21X1_9 ( .A(_349_), .B(_350_), .C(w_C_14_), .Y(_351_) );
NAND2X1 NAND2X1_17 ( .A(_351_), .B(_355_), .Y(_278__14_) );
INVX1 INVX1_9 ( .A(w_C_15_), .Y(_359_) );
OR2X2 OR2X2_9 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_360_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_361_) );
NAND3X1 NAND3X1_10 ( .A(_359_), .B(_361_), .C(_360_), .Y(_362_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_356_) );
AND2X2 AND2X2_10 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_357_) );
OAI21X1 OAI21X1_10 ( .A(_356_), .B(_357_), .C(w_C_15_), .Y(_358_) );
NAND2X1 NAND2X1_19 ( .A(_358_), .B(_362_), .Y(_278__15_) );
INVX1 INVX1_10 ( .A(w_C_16_), .Y(_366_) );
OR2X2 OR2X2_10 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_367_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_368_) );
NAND3X1 NAND3X1_11 ( .A(_366_), .B(_368_), .C(_367_), .Y(_369_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_363_) );
AND2X2 AND2X2_11 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_364_) );
OAI21X1 OAI21X1_11 ( .A(_363_), .B(_364_), .C(w_C_16_), .Y(_365_) );
NAND2X1 NAND2X1_21 ( .A(_365_), .B(_369_), .Y(_278__16_) );
INVX1 INVX1_11 ( .A(w_C_17_), .Y(_373_) );
OR2X2 OR2X2_11 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_374_) );
NAND2X1 NAND2X1_22 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_375_) );
NAND3X1 NAND3X1_12 ( .A(_373_), .B(_375_), .C(_374_), .Y(_376_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_370_) );
AND2X2 AND2X2_12 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_371_) );
OAI21X1 OAI21X1_12 ( .A(_370_), .B(_371_), .C(w_C_17_), .Y(_372_) );
NAND2X1 NAND2X1_23 ( .A(_372_), .B(_376_), .Y(_278__17_) );
INVX1 INVX1_12 ( .A(w_C_18_), .Y(_380_) );
OR2X2 OR2X2_12 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_381_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_382_) );
NAND3X1 NAND3X1_13 ( .A(_380_), .B(_382_), .C(_381_), .Y(_383_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_377_) );
AND2X2 AND2X2_13 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_378_) );
OAI21X1 OAI21X1_13 ( .A(_377_), .B(_378_), .C(w_C_18_), .Y(_379_) );
NAND2X1 NAND2X1_25 ( .A(_379_), .B(_383_), .Y(_278__18_) );
INVX1 INVX1_13 ( .A(w_C_19_), .Y(_387_) );
OR2X2 OR2X2_13 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_388_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_389_) );
NAND3X1 NAND3X1_14 ( .A(_387_), .B(_389_), .C(_388_), .Y(_390_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_384_) );
AND2X2 AND2X2_14 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_385_) );
OAI21X1 OAI21X1_14 ( .A(_384_), .B(_385_), .C(w_C_19_), .Y(_386_) );
NAND2X1 NAND2X1_27 ( .A(_386_), .B(_390_), .Y(_278__19_) );
INVX1 INVX1_14 ( .A(w_C_20_), .Y(_394_) );
OR2X2 OR2X2_14 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_395_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_396_) );
NAND3X1 NAND3X1_15 ( .A(_394_), .B(_396_), .C(_395_), .Y(_397_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_391_) );
AND2X2 AND2X2_15 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_392_) );
OAI21X1 OAI21X1_15 ( .A(_391_), .B(_392_), .C(w_C_20_), .Y(_393_) );
NAND2X1 NAND2X1_29 ( .A(_393_), .B(_397_), .Y(_278__20_) );
INVX1 INVX1_15 ( .A(w_C_21_), .Y(_401_) );
OR2X2 OR2X2_15 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_402_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_403_) );
NAND3X1 NAND3X1_16 ( .A(_401_), .B(_403_), .C(_402_), .Y(_404_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_398_) );
AND2X2 AND2X2_16 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_399_) );
OAI21X1 OAI21X1_16 ( .A(_398_), .B(_399_), .C(w_C_21_), .Y(_400_) );
NAND2X1 NAND2X1_31 ( .A(_400_), .B(_404_), .Y(_278__21_) );
INVX1 INVX1_16 ( .A(w_C_22_), .Y(_408_) );
OR2X2 OR2X2_16 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_409_) );
NAND2X1 NAND2X1_32 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_410_) );
NAND3X1 NAND3X1_17 ( .A(_408_), .B(_410_), .C(_409_), .Y(_411_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_405_) );
AND2X2 AND2X2_17 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_406_) );
OAI21X1 OAI21X1_17 ( .A(_405_), .B(_406_), .C(w_C_22_), .Y(_407_) );
NAND2X1 NAND2X1_33 ( .A(_407_), .B(_411_), .Y(_278__22_) );
INVX1 INVX1_17 ( .A(w_C_23_), .Y(_415_) );
OR2X2 OR2X2_17 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_416_) );
NAND2X1 NAND2X1_34 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_417_) );
NAND3X1 NAND3X1_18 ( .A(_415_), .B(_417_), .C(_416_), .Y(_418_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_412_) );
AND2X2 AND2X2_18 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_413_) );
OAI21X1 OAI21X1_18 ( .A(_412_), .B(_413_), .C(w_C_23_), .Y(_414_) );
NAND2X1 NAND2X1_35 ( .A(_414_), .B(_418_), .Y(_278__23_) );
INVX1 INVX1_18 ( .A(w_C_24_), .Y(_422_) );
OR2X2 OR2X2_18 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_423_) );
NAND2X1 NAND2X1_36 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_424_) );
NAND3X1 NAND3X1_19 ( .A(_422_), .B(_424_), .C(_423_), .Y(_425_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_419_) );
AND2X2 AND2X2_19 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_420_) );
OAI21X1 OAI21X1_19 ( .A(_419_), .B(_420_), .C(w_C_24_), .Y(_421_) );
NAND2X1 NAND2X1_37 ( .A(_421_), .B(_425_), .Y(_278__24_) );
INVX1 INVX1_19 ( .A(w_C_25_), .Y(_429_) );
OR2X2 OR2X2_19 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_430_) );
NAND2X1 NAND2X1_38 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_431_) );
NAND3X1 NAND3X1_20 ( .A(_429_), .B(_431_), .C(_430_), .Y(_432_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_426_) );
AND2X2 AND2X2_20 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_427_) );
OAI21X1 OAI21X1_20 ( .A(_426_), .B(_427_), .C(w_C_25_), .Y(_428_) );
NAND2X1 NAND2X1_39 ( .A(_428_), .B(_432_), .Y(_278__25_) );
INVX1 INVX1_20 ( .A(w_C_26_), .Y(_436_) );
OR2X2 OR2X2_20 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_437_) );
NAND2X1 NAND2X1_40 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_438_) );
NAND3X1 NAND3X1_21 ( .A(_436_), .B(_438_), .C(_437_), .Y(_439_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_433_) );
AND2X2 AND2X2_21 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_434_) );
OAI21X1 OAI21X1_21 ( .A(_433_), .B(_434_), .C(w_C_26_), .Y(_435_) );
NAND2X1 NAND2X1_41 ( .A(_435_), .B(_439_), .Y(_278__26_) );
INVX1 INVX1_21 ( .A(w_C_27_), .Y(_443_) );
OR2X2 OR2X2_21 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_444_) );
NAND2X1 NAND2X1_42 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_445_) );
NAND3X1 NAND3X1_22 ( .A(_443_), .B(_445_), .C(_444_), .Y(_446_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_440_) );
AND2X2 AND2X2_22 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_441_) );
OAI21X1 OAI21X1_22 ( .A(_440_), .B(_441_), .C(w_C_27_), .Y(_442_) );
NAND2X1 NAND2X1_43 ( .A(_442_), .B(_446_), .Y(_278__27_) );
INVX1 INVX1_22 ( .A(w_C_28_), .Y(_450_) );
OR2X2 OR2X2_22 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_451_) );
NAND2X1 NAND2X1_44 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_452_) );
NAND3X1 NAND3X1_23 ( .A(_450_), .B(_452_), .C(_451_), .Y(_453_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_447_) );
AND2X2 AND2X2_23 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_448_) );
OAI21X1 OAI21X1_23 ( .A(_447_), .B(_448_), .C(w_C_28_), .Y(_449_) );
NAND2X1 NAND2X1_45 ( .A(_449_), .B(_453_), .Y(_278__28_) );
INVX1 INVX1_23 ( .A(w_C_29_), .Y(_457_) );
OR2X2 OR2X2_23 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_458_) );
NAND2X1 NAND2X1_46 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_459_) );
NAND3X1 NAND3X1_24 ( .A(_457_), .B(_459_), .C(_458_), .Y(_460_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_454_) );
AND2X2 AND2X2_24 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_455_) );
OAI21X1 OAI21X1_24 ( .A(_454_), .B(_455_), .C(w_C_29_), .Y(_456_) );
NAND2X1 NAND2X1_47 ( .A(_456_), .B(_460_), .Y(_278__29_) );
INVX1 INVX1_24 ( .A(w_C_30_), .Y(_464_) );
OR2X2 OR2X2_24 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_465_) );
NAND2X1 NAND2X1_48 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_466_) );
NAND3X1 NAND3X1_25 ( .A(_464_), .B(_466_), .C(_465_), .Y(_467_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_461_) );
AND2X2 AND2X2_25 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_462_) );
OAI21X1 OAI21X1_25 ( .A(_461_), .B(_462_), .C(w_C_30_), .Y(_463_) );
NAND2X1 NAND2X1_49 ( .A(_463_), .B(_467_), .Y(_278__30_) );
INVX1 INVX1_25 ( .A(w_C_31_), .Y(_471_) );
OR2X2 OR2X2_25 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_472_) );
NAND2X1 NAND2X1_50 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_473_) );
NAND3X1 NAND3X1_26 ( .A(_471_), .B(_473_), .C(_472_), .Y(_474_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_468_) );
AND2X2 AND2X2_26 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_469_) );
OAI21X1 OAI21X1_26 ( .A(_468_), .B(_469_), .C(w_C_31_), .Y(_470_) );
NAND2X1 NAND2X1_51 ( .A(_470_), .B(_474_), .Y(_278__31_) );
INVX1 INVX1_26 ( .A(w_C_32_), .Y(_478_) );
OR2X2 OR2X2_26 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_479_) );
NAND2X1 NAND2X1_52 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_480_) );
NAND3X1 NAND3X1_27 ( .A(_478_), .B(_480_), .C(_479_), .Y(_481_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_475_) );
AND2X2 AND2X2_27 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_476_) );
OAI21X1 OAI21X1_27 ( .A(_475_), .B(_476_), .C(w_C_32_), .Y(_477_) );
NAND2X1 NAND2X1_53 ( .A(_477_), .B(_481_), .Y(_278__32_) );
INVX1 INVX1_27 ( .A(w_C_33_), .Y(_485_) );
OR2X2 OR2X2_27 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_486_) );
NAND2X1 NAND2X1_54 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_487_) );
NAND3X1 NAND3X1_28 ( .A(_485_), .B(_487_), .C(_486_), .Y(_488_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_482_) );
AND2X2 AND2X2_28 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_483_) );
OAI21X1 OAI21X1_28 ( .A(_482_), .B(_483_), .C(w_C_33_), .Y(_484_) );
NAND2X1 NAND2X1_55 ( .A(_484_), .B(_488_), .Y(_278__33_) );
INVX1 INVX1_28 ( .A(w_C_34_), .Y(_492_) );
OR2X2 OR2X2_28 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_493_) );
NAND2X1 NAND2X1_56 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_494_) );
NAND3X1 NAND3X1_29 ( .A(_492_), .B(_494_), .C(_493_), .Y(_495_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_489_) );
AND2X2 AND2X2_29 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_490_) );
OAI21X1 OAI21X1_29 ( .A(_489_), .B(_490_), .C(w_C_34_), .Y(_491_) );
NAND2X1 NAND2X1_57 ( .A(_491_), .B(_495_), .Y(_278__34_) );
INVX1 INVX1_29 ( .A(w_C_35_), .Y(_499_) );
OR2X2 OR2X2_29 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_500_) );
NAND2X1 NAND2X1_58 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_501_) );
NAND3X1 NAND3X1_30 ( .A(_499_), .B(_501_), .C(_500_), .Y(_502_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_496_) );
AND2X2 AND2X2_30 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_497_) );
OAI21X1 OAI21X1_30 ( .A(_496_), .B(_497_), .C(w_C_35_), .Y(_498_) );
NAND2X1 NAND2X1_59 ( .A(_498_), .B(_502_), .Y(_278__35_) );
INVX1 INVX1_30 ( .A(w_C_36_), .Y(_506_) );
OR2X2 OR2X2_30 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_507_) );
NAND2X1 NAND2X1_60 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_508_) );
NAND3X1 NAND3X1_31 ( .A(_506_), .B(_508_), .C(_507_), .Y(_509_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_503_) );
AND2X2 AND2X2_31 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_504_) );
OAI21X1 OAI21X1_31 ( .A(_503_), .B(_504_), .C(w_C_36_), .Y(_505_) );
NAND2X1 NAND2X1_61 ( .A(_505_), .B(_509_), .Y(_278__36_) );
INVX1 INVX1_31 ( .A(w_C_37_), .Y(_513_) );
OR2X2 OR2X2_31 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_514_) );
NAND2X1 NAND2X1_62 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_515_) );
NAND3X1 NAND3X1_32 ( .A(_513_), .B(_515_), .C(_514_), .Y(_516_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_510_) );
AND2X2 AND2X2_32 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_511_) );
OAI21X1 OAI21X1_32 ( .A(_510_), .B(_511_), .C(w_C_37_), .Y(_512_) );
NAND2X1 NAND2X1_63 ( .A(_512_), .B(_516_), .Y(_278__37_) );
INVX1 INVX1_32 ( .A(w_C_38_), .Y(_520_) );
OR2X2 OR2X2_32 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_521_) );
NAND2X1 NAND2X1_64 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_522_) );
NAND3X1 NAND3X1_33 ( .A(_520_), .B(_522_), .C(_521_), .Y(_523_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_517_) );
AND2X2 AND2X2_33 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_518_) );
OAI21X1 OAI21X1_33 ( .A(_517_), .B(_518_), .C(w_C_38_), .Y(_519_) );
NAND2X1 NAND2X1_65 ( .A(_519_), .B(_523_), .Y(_278__38_) );
INVX1 INVX1_33 ( .A(w_C_39_), .Y(_527_) );
OR2X2 OR2X2_33 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_528_) );
NAND2X1 NAND2X1_66 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_529_) );
NAND3X1 NAND3X1_34 ( .A(_527_), .B(_529_), .C(_528_), .Y(_530_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_524_) );
AND2X2 AND2X2_34 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_525_) );
OAI21X1 OAI21X1_34 ( .A(_524_), .B(_525_), .C(w_C_39_), .Y(_526_) );
NAND2X1 NAND2X1_67 ( .A(_526_), .B(_530_), .Y(_278__39_) );
INVX1 INVX1_34 ( .A(w_C_40_), .Y(_534_) );
OR2X2 OR2X2_34 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_535_) );
NAND2X1 NAND2X1_68 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_536_) );
NAND3X1 NAND3X1_35 ( .A(_534_), .B(_536_), .C(_535_), .Y(_537_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_531_) );
AND2X2 AND2X2_35 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_532_) );
OAI21X1 OAI21X1_35 ( .A(_531_), .B(_532_), .C(w_C_40_), .Y(_533_) );
NAND2X1 NAND2X1_69 ( .A(_533_), .B(_537_), .Y(_278__40_) );
INVX1 INVX1_35 ( .A(w_C_41_), .Y(_541_) );
OR2X2 OR2X2_35 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_542_) );
NAND2X1 NAND2X1_70 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_543_) );
NAND3X1 NAND3X1_36 ( .A(_541_), .B(_543_), .C(_542_), .Y(_544_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_538_) );
AND2X2 AND2X2_36 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_539_) );
OAI21X1 OAI21X1_36 ( .A(_538_), .B(_539_), .C(w_C_41_), .Y(_540_) );
NAND2X1 NAND2X1_71 ( .A(_540_), .B(_544_), .Y(_278__41_) );
INVX1 INVX1_36 ( .A(w_C_42_), .Y(_548_) );
OR2X2 OR2X2_36 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_549_) );
NAND2X1 NAND2X1_72 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_550_) );
NAND3X1 NAND3X1_37 ( .A(_548_), .B(_550_), .C(_549_), .Y(_551_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_545_) );
AND2X2 AND2X2_37 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_546_) );
OAI21X1 OAI21X1_37 ( .A(_545_), .B(_546_), .C(w_C_42_), .Y(_547_) );
NAND2X1 NAND2X1_73 ( .A(_547_), .B(_551_), .Y(_278__42_) );
INVX1 INVX1_37 ( .A(w_C_43_), .Y(_555_) );
OR2X2 OR2X2_37 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_556_) );
NAND2X1 NAND2X1_74 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_557_) );
NAND3X1 NAND3X1_38 ( .A(_555_), .B(_557_), .C(_556_), .Y(_558_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_552_) );
AND2X2 AND2X2_38 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_553_) );
OAI21X1 OAI21X1_38 ( .A(_552_), .B(_553_), .C(w_C_43_), .Y(_554_) );
NAND2X1 NAND2X1_75 ( .A(_554_), .B(_558_), .Y(_278__43_) );
INVX1 INVX1_38 ( .A(w_C_44_), .Y(_562_) );
OR2X2 OR2X2_38 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_563_) );
NAND2X1 NAND2X1_76 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_564_) );
NAND3X1 NAND3X1_39 ( .A(_562_), .B(_564_), .C(_563_), .Y(_565_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_559_) );
AND2X2 AND2X2_39 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_560_) );
OAI21X1 OAI21X1_39 ( .A(_559_), .B(_560_), .C(w_C_44_), .Y(_561_) );
NAND2X1 NAND2X1_77 ( .A(_561_), .B(_565_), .Y(_278__44_) );
INVX1 INVX1_39 ( .A(w_C_45_), .Y(_569_) );
OR2X2 OR2X2_39 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_570_) );
NAND2X1 NAND2X1_78 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_571_) );
NAND3X1 NAND3X1_40 ( .A(_569_), .B(_571_), .C(_570_), .Y(_572_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_566_) );
AND2X2 AND2X2_40 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_567_) );
OAI21X1 OAI21X1_40 ( .A(_566_), .B(_567_), .C(w_C_45_), .Y(_568_) );
NAND2X1 NAND2X1_79 ( .A(_568_), .B(_572_), .Y(_278__45_) );
INVX1 INVX1_40 ( .A(w_C_46_), .Y(_576_) );
OR2X2 OR2X2_40 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_577_) );
NAND2X1 NAND2X1_80 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_578_) );
NAND3X1 NAND3X1_41 ( .A(_576_), .B(_578_), .C(_577_), .Y(_579_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_573_) );
AND2X2 AND2X2_41 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_574_) );
OAI21X1 OAI21X1_41 ( .A(_573_), .B(_574_), .C(w_C_46_), .Y(_575_) );
NAND2X1 NAND2X1_81 ( .A(_575_), .B(_579_), .Y(_278__46_) );
INVX1 INVX1_41 ( .A(1'b0), .Y(_583_) );
OR2X2 OR2X2_41 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_584_) );
NAND2X1 NAND2X1_82 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_585_) );
NAND3X1 NAND3X1_42 ( .A(_583_), .B(_585_), .C(_584_), .Y(_586_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_580_) );
AND2X2 AND2X2_42 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_581_) );
OAI21X1 OAI21X1_42 ( .A(_580_), .B(_581_), .C(1'b0), .Y(_582_) );
NAND2X1 NAND2X1_83 ( .A(_582_), .B(_586_), .Y(_278__0_) );
INVX1 INVX1_42 ( .A(w_C_1_), .Y(_590_) );
OR2X2 OR2X2_42 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_591_) );
NAND2X1 NAND2X1_84 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_592_) );
NAND3X1 NAND3X1_43 ( .A(_590_), .B(_592_), .C(_591_), .Y(_593_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_587_) );
AND2X2 AND2X2_43 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_588_) );
OAI21X1 OAI21X1_43 ( .A(_587_), .B(_588_), .C(w_C_1_), .Y(_589_) );
NAND2X1 NAND2X1_85 ( .A(_589_), .B(_593_), .Y(_278__1_) );
INVX1 INVX1_43 ( .A(w_C_2_), .Y(_597_) );
OR2X2 OR2X2_43 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_598_) );
NAND2X1 NAND2X1_86 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_599_) );
NAND3X1 NAND3X1_44 ( .A(_597_), .B(_599_), .C(_598_), .Y(_600_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_594_) );
AND2X2 AND2X2_44 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_595_) );
OAI21X1 OAI21X1_44 ( .A(_594_), .B(_595_), .C(w_C_2_), .Y(_596_) );
NAND2X1 NAND2X1_87 ( .A(_596_), .B(_600_), .Y(_278__2_) );
INVX1 INVX1_44 ( .A(w_C_3_), .Y(_604_) );
OR2X2 OR2X2_44 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_605_) );
NAND2X1 NAND2X1_88 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_606_) );
NAND3X1 NAND3X1_45 ( .A(_604_), .B(_606_), .C(_605_), .Y(_607_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_601_) );
AND2X2 AND2X2_45 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_602_) );
OAI21X1 OAI21X1_45 ( .A(_601_), .B(_602_), .C(w_C_3_), .Y(_603_) );
NAND2X1 NAND2X1_89 ( .A(_603_), .B(_607_), .Y(_278__3_) );
NAND3X1 NAND3X1_46 ( .A(_228_), .B(_230_), .C(_221_), .Y(_231_) );
AND2X2 AND2X2_46 ( .A(_231_), .B(_226_), .Y(_232_) );
INVX1 INVX1_45 ( .A(_232_), .Y(w_C_37_) );
AND2X2 AND2X2_47 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_233_) );
INVX1 INVX1_46 ( .A(_233_), .Y(_234_) );
NAND3X1 NAND3X1_47 ( .A(_226_), .B(_234_), .C(_231_), .Y(_235_) );
OAI21X1 OAI21X1_46 ( .A(i_add2[37]), .B(i_add1[37]), .C(_235_), .Y(_236_) );
INVX1 INVX1_47 ( .A(_236_), .Y(w_C_38_) );
NAND2X1 NAND2X1_90 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_237_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_238_) );
OAI21X1 OAI21X1_47 ( .A(_238_), .B(_236_), .C(_237_), .Y(w_C_39_) );
OR2X2 OR2X2_45 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_239_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_240_) );
INVX1 INVX1_48 ( .A(_240_), .Y(_241_) );
INVX1 INVX1_49 ( .A(_238_), .Y(_242_) );
NAND3X1 NAND3X1_48 ( .A(_241_), .B(_242_), .C(_235_), .Y(_243_) );
NAND2X1 NAND2X1_91 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_244_) );
NAND3X1 NAND3X1_49 ( .A(_237_), .B(_244_), .C(_243_), .Y(_245_) );
AND2X2 AND2X2_48 ( .A(_245_), .B(_239_), .Y(w_C_40_) );
INVX1 INVX1_50 ( .A(i_add2[40]), .Y(_246_) );
INVX1 INVX1_51 ( .A(i_add1[40]), .Y(_247_) );
NAND2X1 NAND2X1_92 ( .A(_246_), .B(_247_), .Y(_248_) );
NAND3X1 NAND3X1_50 ( .A(_239_), .B(_248_), .C(_245_), .Y(_249_) );
OAI21X1 OAI21X1_48 ( .A(_246_), .B(_247_), .C(_249_), .Y(w_C_41_) );
INVX1 INVX1_52 ( .A(i_add2[41]), .Y(_250_) );
INVX1 INVX1_53 ( .A(i_add1[41]), .Y(_251_) );
OAI21X1 OAI21X1_49 ( .A(i_add2[41]), .B(i_add1[41]), .C(w_C_41_), .Y(_252_) );
OAI21X1 OAI21X1_50 ( .A(_250_), .B(_251_), .C(_252_), .Y(w_C_42_) );
INVX1 INVX1_54 ( .A(i_add2[42]), .Y(_253_) );
INVX1 INVX1_55 ( .A(i_add1[42]), .Y(_254_) );
NOR2X1 NOR2X1_48 ( .A(_253_), .B(_254_), .Y(_255_) );
OR2X2 OR2X2_46 ( .A(w_C_42_), .B(_255_), .Y(_256_) );
OAI21X1 OAI21X1_51 ( .A(i_add2[42]), .B(i_add1[42]), .C(_256_), .Y(_257_) );
INVX1 INVX1_56 ( .A(_257_), .Y(w_C_43_) );
NAND2X1 NAND2X1_93 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_258_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_259_) );
OAI21X1 OAI21X1_52 ( .A(_259_), .B(_257_), .C(_258_), .Y(w_C_44_) );
NAND2X1 NAND2X1_94 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_260_) );
INVX1 INVX1_57 ( .A(_259_), .Y(_261_) );
INVX1 INVX1_58 ( .A(_255_), .Y(_262_) );
NAND2X1 NAND2X1_95 ( .A(_250_), .B(_251_), .Y(_263_) );
NAND2X1 NAND2X1_96 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_264_) );
NAND2X1 NAND2X1_97 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_265_) );
NAND3X1 NAND3X1_51 ( .A(_264_), .B(_265_), .C(_249_), .Y(_266_) );
NAND2X1 NAND2X1_98 ( .A(_253_), .B(_254_), .Y(_267_) );
NAND3X1 NAND3X1_52 ( .A(_263_), .B(_267_), .C(_266_), .Y(_268_) );
NAND3X1 NAND3X1_53 ( .A(_262_), .B(_258_), .C(_268_), .Y(_269_) );
OR2X2 OR2X2_47 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_270_) );
NAND3X1 NAND3X1_54 ( .A(_261_), .B(_270_), .C(_269_), .Y(_271_) );
NAND2X1 NAND2X1_99 ( .A(_260_), .B(_271_), .Y(w_C_45_) );
OR2X2 OR2X2_48 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_272_) );
NAND2X1 NAND2X1_100 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_273_) );
NAND3X1 NAND3X1_55 ( .A(_260_), .B(_273_), .C(_271_), .Y(_274_) );
AND2X2 AND2X2_49 ( .A(_274_), .B(_272_), .Y(w_C_46_) );
NAND2X1 NAND2X1_101 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_275_) );
OR2X2 OR2X2_49 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_276_) );
NAND3X1 NAND3X1_56 ( .A(_272_), .B(_276_), .C(_274_), .Y(_277_) );
NAND2X1 NAND2X1_102 ( .A(_275_), .B(_277_), .Y(w_C_47_) );
NAND2X1 NAND2X1_103 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_59 ( .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_104 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_105 ( .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_53 ( .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_60 ( .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_106 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_50 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_51 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_57 ( .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_107 ( .A(_4_), .B(_7_), .Y(w_C_3_) );
INVX1 INVX1_61 ( .A(i_add2[3]), .Y(_8_) );
INVX1 INVX1_62 ( .A(i_add1[3]), .Y(_9_) );
NAND2X1 NAND2X1_108 ( .A(_8_), .B(_9_), .Y(_10_) );
NAND2X1 NAND2X1_109 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_11_) );
NAND3X1 NAND3X1_58 ( .A(_4_), .B(_11_), .C(_7_), .Y(_12_) );
AND2X2 AND2X2_50 ( .A(_12_), .B(_10_), .Y(w_C_4_) );
NAND2X1 NAND2X1_110 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
OR2X2 OR2X2_52 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_14_) );
NAND3X1 NAND3X1_59 ( .A(_10_), .B(_14_), .C(_12_), .Y(_15_) );
NAND2X1 NAND2X1_111 ( .A(_13_), .B(_15_), .Y(w_C_5_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_16_) );
INVX1 INVX1_63 ( .A(_16_), .Y(_17_) );
NAND2X1 NAND2X1_112 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_18_) );
NAND3X1 NAND3X1_60 ( .A(_13_), .B(_18_), .C(_15_), .Y(_19_) );
AND2X2 AND2X2_51 ( .A(_19_), .B(_17_), .Y(w_C_6_) );
INVX1 INVX1_64 ( .A(i_add2[6]), .Y(_20_) );
INVX1 INVX1_65 ( .A(i_add1[6]), .Y(_21_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_66 ( .A(_22_), .Y(_23_) );
NAND3X1 NAND3X1_61 ( .A(_17_), .B(_23_), .C(_19_), .Y(_24_) );
OAI21X1 OAI21X1_54 ( .A(_20_), .B(_21_), .C(_24_), .Y(w_C_7_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_25_) );
INVX1 INVX1_67 ( .A(_25_), .Y(_26_) );
NOR2X1 NOR2X1_53 ( .A(_20_), .B(_21_), .Y(_27_) );
INVX1 INVX1_68 ( .A(_27_), .Y(_28_) );
INVX1 INVX1_69 ( .A(i_add2[7]), .Y(_29_) );
INVX1 INVX1_70 ( .A(i_add1[7]), .Y(_30_) );
NOR2X1 NOR2X1_54 ( .A(_29_), .B(_30_), .Y(_31_) );
INVX1 INVX1_71 ( .A(_31_), .Y(_32_) );
NAND3X1 NAND3X1_62 ( .A(_28_), .B(_32_), .C(_24_), .Y(_33_) );
AND2X2 AND2X2_52 ( .A(_33_), .B(_26_), .Y(w_C_8_) );
INVX1 INVX1_72 ( .A(i_add2[8]), .Y(_34_) );
INVX1 INVX1_73 ( .A(i_add1[8]), .Y(_35_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_36_) );
INVX1 INVX1_74 ( .A(_36_), .Y(_37_) );
NAND3X1 NAND3X1_63 ( .A(_26_), .B(_37_), .C(_33_), .Y(_38_) );
OAI21X1 OAI21X1_55 ( .A(_34_), .B(_35_), .C(_38_), .Y(w_C_9_) );
NOR2X1 NOR2X1_56 ( .A(_34_), .B(_35_), .Y(_39_) );
INVX1 INVX1_75 ( .A(_39_), .Y(_40_) );
AND2X2 AND2X2_53 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_41_) );
INVX1 INVX1_76 ( .A(_41_), .Y(_42_) );
NAND3X1 NAND3X1_64 ( .A(_40_), .B(_42_), .C(_38_), .Y(_43_) );
OAI21X1 OAI21X1_56 ( .A(i_add2[9]), .B(i_add1[9]), .C(_43_), .Y(_44_) );
INVX1 INVX1_77 ( .A(_44_), .Y(w_C_10_) );
INVX1 INVX1_78 ( .A(i_add2[10]), .Y(_45_) );
INVX1 INVX1_79 ( .A(i_add1[10]), .Y(_46_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_47_) );
INVX1 INVX1_80 ( .A(_47_), .Y(_48_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_49_) );
INVX1 INVX1_81 ( .A(_49_), .Y(_50_) );
NAND3X1 NAND3X1_65 ( .A(_48_), .B(_50_), .C(_43_), .Y(_51_) );
OAI21X1 OAI21X1_57 ( .A(_45_), .B(_46_), .C(_51_), .Y(w_C_11_) );
NOR2X1 NOR2X1_59 ( .A(_45_), .B(_46_), .Y(_52_) );
INVX1 INVX1_82 ( .A(_52_), .Y(_53_) );
AND2X2 AND2X2_54 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_54_) );
INVX1 INVX1_83 ( .A(_54_), .Y(_55_) );
NAND3X1 NAND3X1_66 ( .A(_53_), .B(_55_), .C(_51_), .Y(_56_) );
OAI21X1 OAI21X1_58 ( .A(i_add2[11]), .B(i_add1[11]), .C(_56_), .Y(_57_) );
INVX1 INVX1_84 ( .A(_57_), .Y(w_C_12_) );
INVX1 INVX1_85 ( .A(i_add2[12]), .Y(_58_) );
INVX1 INVX1_86 ( .A(i_add1[12]), .Y(_59_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_60_) );
INVX1 INVX1_87 ( .A(_60_), .Y(_61_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_62_) );
INVX1 INVX1_88 ( .A(_62_), .Y(_63_) );
NAND3X1 NAND3X1_67 ( .A(_61_), .B(_63_), .C(_56_), .Y(_64_) );
OAI21X1 OAI21X1_59 ( .A(_58_), .B(_59_), .C(_64_), .Y(w_C_13_) );
NOR2X1 NOR2X1_62 ( .A(_58_), .B(_59_), .Y(_65_) );
INVX1 INVX1_89 ( .A(_65_), .Y(_66_) );
AND2X2 AND2X2_55 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_67_) );
INVX1 INVX1_90 ( .A(_67_), .Y(_68_) );
NAND3X1 NAND3X1_68 ( .A(_66_), .B(_68_), .C(_64_), .Y(_69_) );
OAI21X1 OAI21X1_60 ( .A(i_add2[13]), .B(i_add1[13]), .C(_69_), .Y(_70_) );
INVX1 INVX1_91 ( .A(_70_), .Y(w_C_14_) );
INVX1 INVX1_92 ( .A(i_add2[14]), .Y(_71_) );
INVX1 INVX1_93 ( .A(i_add1[14]), .Y(_72_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_73_) );
INVX1 INVX1_94 ( .A(_73_), .Y(_74_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_75_) );
INVX1 INVX1_95 ( .A(_75_), .Y(_76_) );
NAND3X1 NAND3X1_69 ( .A(_74_), .B(_76_), .C(_69_), .Y(_77_) );
OAI21X1 OAI21X1_61 ( .A(_71_), .B(_72_), .C(_77_), .Y(w_C_15_) );
NOR2X1 NOR2X1_65 ( .A(_71_), .B(_72_), .Y(_78_) );
INVX1 INVX1_96 ( .A(_78_), .Y(_79_) );
AND2X2 AND2X2_56 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_80_) );
INVX1 INVX1_97 ( .A(_80_), .Y(_81_) );
NAND3X1 NAND3X1_70 ( .A(_79_), .B(_81_), .C(_77_), .Y(_82_) );
OAI21X1 OAI21X1_62 ( .A(i_add2[15]), .B(i_add1[15]), .C(_82_), .Y(_83_) );
INVX1 INVX1_98 ( .A(_83_), .Y(w_C_16_) );
INVX1 INVX1_99 ( .A(i_add2[16]), .Y(_84_) );
INVX1 INVX1_100 ( .A(i_add1[16]), .Y(_85_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_86_) );
INVX1 INVX1_101 ( .A(_86_), .Y(_87_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_88_) );
INVX1 INVX1_102 ( .A(_88_), .Y(_89_) );
NAND3X1 NAND3X1_71 ( .A(_87_), .B(_89_), .C(_82_), .Y(_90_) );
OAI21X1 OAI21X1_63 ( .A(_84_), .B(_85_), .C(_90_), .Y(w_C_17_) );
NOR2X1 NOR2X1_68 ( .A(_84_), .B(_85_), .Y(_91_) );
INVX1 INVX1_103 ( .A(_91_), .Y(_92_) );
AND2X2 AND2X2_57 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_93_) );
INVX1 INVX1_104 ( .A(_93_), .Y(_94_) );
NAND3X1 NAND3X1_72 ( .A(_92_), .B(_94_), .C(_90_), .Y(_95_) );
OAI21X1 OAI21X1_64 ( .A(i_add2[17]), .B(i_add1[17]), .C(_95_), .Y(_96_) );
INVX1 INVX1_105 ( .A(_96_), .Y(w_C_18_) );
INVX1 INVX1_106 ( .A(i_add2[18]), .Y(_97_) );
INVX1 INVX1_107 ( .A(i_add1[18]), .Y(_98_) );
NOR2X1 NOR2X1_69 ( .A(_97_), .B(_98_), .Y(_99_) );
INVX1 INVX1_108 ( .A(_99_), .Y(_100_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_101_) );
INVX1 INVX1_109 ( .A(_101_), .Y(_102_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_103_) );
INVX1 INVX1_110 ( .A(_103_), .Y(_104_) );
NAND3X1 NAND3X1_73 ( .A(_102_), .B(_104_), .C(_95_), .Y(_105_) );
AND2X2 AND2X2_58 ( .A(_105_), .B(_100_), .Y(_106_) );
INVX1 INVX1_111 ( .A(_106_), .Y(w_C_19_) );
AND2X2 AND2X2_59 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_107_) );
INVX1 INVX1_112 ( .A(_107_), .Y(_108_) );
NAND3X1 NAND3X1_74 ( .A(_100_), .B(_108_), .C(_105_), .Y(_109_) );
OAI21X1 OAI21X1_65 ( .A(i_add2[19]), .B(i_add1[19]), .C(_109_), .Y(_110_) );
INVX1 INVX1_113 ( .A(_110_), .Y(w_C_20_) );
INVX1 INVX1_114 ( .A(i_add2[20]), .Y(_111_) );
INVX1 INVX1_115 ( .A(i_add1[20]), .Y(_112_) );
NOR2X1 NOR2X1_72 ( .A(_111_), .B(_112_), .Y(_113_) );
INVX1 INVX1_116 ( .A(_113_), .Y(_114_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_115_) );
INVX1 INVX1_117 ( .A(_115_), .Y(_116_) );
NOR2X1 NOR2X1_74 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_117_) );
INVX1 INVX1_118 ( .A(_117_), .Y(_118_) );
NAND3X1 NAND3X1_75 ( .A(_116_), .B(_118_), .C(_109_), .Y(_119_) );
AND2X2 AND2X2_60 ( .A(_119_), .B(_114_), .Y(_120_) );
INVX1 INVX1_119 ( .A(_120_), .Y(w_C_21_) );
AND2X2 AND2X2_61 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_121_) );
INVX1 INVX1_120 ( .A(_121_), .Y(_122_) );
NAND3X1 NAND3X1_76 ( .A(_114_), .B(_122_), .C(_119_), .Y(_123_) );
OAI21X1 OAI21X1_66 ( .A(i_add2[21]), .B(i_add1[21]), .C(_123_), .Y(_124_) );
INVX1 INVX1_121 ( .A(_124_), .Y(w_C_22_) );
INVX1 INVX1_122 ( .A(i_add2[22]), .Y(_125_) );
INVX1 INVX1_123 ( .A(i_add1[22]), .Y(_126_) );
NOR2X1 NOR2X1_75 ( .A(_125_), .B(_126_), .Y(_127_) );
INVX1 INVX1_124 ( .A(_127_), .Y(_128_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_129_) );
INVX1 INVX1_125 ( .A(_129_), .Y(_130_) );
NOR2X1 NOR2X1_77 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_131_) );
INVX1 INVX1_126 ( .A(_131_), .Y(_132_) );
NAND3X1 NAND3X1_77 ( .A(_130_), .B(_132_), .C(_123_), .Y(_133_) );
AND2X2 AND2X2_62 ( .A(_133_), .B(_128_), .Y(_134_) );
INVX1 INVX1_127 ( .A(_134_), .Y(w_C_23_) );
AND2X2 AND2X2_63 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_135_) );
INVX1 INVX1_128 ( .A(_135_), .Y(_136_) );
NAND3X1 NAND3X1_78 ( .A(_128_), .B(_136_), .C(_133_), .Y(_137_) );
OAI21X1 OAI21X1_67 ( .A(i_add2[23]), .B(i_add1[23]), .C(_137_), .Y(_138_) );
INVX1 INVX1_129 ( .A(_138_), .Y(w_C_24_) );
INVX1 INVX1_130 ( .A(i_add2[24]), .Y(_139_) );
INVX1 INVX1_131 ( .A(i_add1[24]), .Y(_140_) );
NOR2X1 NOR2X1_78 ( .A(_139_), .B(_140_), .Y(_141_) );
INVX1 INVX1_132 ( .A(_141_), .Y(_142_) );
NOR2X1 NOR2X1_79 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_143_) );
INVX1 INVX1_133 ( .A(_143_), .Y(_144_) );
NOR2X1 NOR2X1_80 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_145_) );
INVX1 INVX1_134 ( .A(_145_), .Y(_146_) );
NAND3X1 NAND3X1_79 ( .A(_144_), .B(_146_), .C(_137_), .Y(_147_) );
AND2X2 AND2X2_64 ( .A(_147_), .B(_142_), .Y(_148_) );
INVX1 INVX1_135 ( .A(_148_), .Y(w_C_25_) );
AND2X2 AND2X2_65 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_149_) );
INVX1 INVX1_136 ( .A(_149_), .Y(_150_) );
NAND3X1 NAND3X1_80 ( .A(_142_), .B(_150_), .C(_147_), .Y(_151_) );
OAI21X1 OAI21X1_68 ( .A(i_add2[25]), .B(i_add1[25]), .C(_151_), .Y(_152_) );
INVX1 INVX1_137 ( .A(_152_), .Y(w_C_26_) );
INVX1 INVX1_138 ( .A(i_add2[26]), .Y(_153_) );
INVX1 INVX1_139 ( .A(i_add1[26]), .Y(_154_) );
NOR2X1 NOR2X1_81 ( .A(_153_), .B(_154_), .Y(_155_) );
INVX1 INVX1_140 ( .A(_155_), .Y(_156_) );
NOR2X1 NOR2X1_82 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_157_) );
INVX1 INVX1_141 ( .A(_157_), .Y(_158_) );
NOR2X1 NOR2X1_83 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_159_) );
INVX1 INVX1_142 ( .A(_159_), .Y(_160_) );
NAND3X1 NAND3X1_81 ( .A(_158_), .B(_160_), .C(_151_), .Y(_161_) );
AND2X2 AND2X2_66 ( .A(_161_), .B(_156_), .Y(_162_) );
INVX1 INVX1_143 ( .A(_162_), .Y(w_C_27_) );
AND2X2 AND2X2_67 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_163_) );
INVX1 INVX1_144 ( .A(_163_), .Y(_164_) );
NAND3X1 NAND3X1_82 ( .A(_156_), .B(_164_), .C(_161_), .Y(_165_) );
OAI21X1 OAI21X1_69 ( .A(i_add2[27]), .B(i_add1[27]), .C(_165_), .Y(_166_) );
INVX1 INVX1_145 ( .A(_166_), .Y(w_C_28_) );
INVX1 INVX1_146 ( .A(i_add2[28]), .Y(_167_) );
INVX1 INVX1_147 ( .A(i_add1[28]), .Y(_168_) );
NOR2X1 NOR2X1_84 ( .A(_167_), .B(_168_), .Y(_169_) );
INVX1 INVX1_148 ( .A(_169_), .Y(_170_) );
NOR2X1 NOR2X1_85 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_171_) );
INVX1 INVX1_149 ( .A(_171_), .Y(_172_) );
NOR2X1 NOR2X1_86 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_173_) );
INVX1 INVX1_150 ( .A(_173_), .Y(_174_) );
NAND3X1 NAND3X1_83 ( .A(_172_), .B(_174_), .C(_165_), .Y(_175_) );
AND2X2 AND2X2_68 ( .A(_175_), .B(_170_), .Y(_176_) );
INVX1 INVX1_151 ( .A(_176_), .Y(w_C_29_) );
AND2X2 AND2X2_69 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_177_) );
INVX1 INVX1_152 ( .A(_177_), .Y(_178_) );
NAND3X1 NAND3X1_84 ( .A(_170_), .B(_178_), .C(_175_), .Y(_179_) );
OAI21X1 OAI21X1_70 ( .A(i_add2[29]), .B(i_add1[29]), .C(_179_), .Y(_180_) );
INVX1 INVX1_153 ( .A(_180_), .Y(w_C_30_) );
INVX1 INVX1_154 ( .A(i_add2[30]), .Y(_181_) );
INVX1 INVX1_155 ( .A(i_add1[30]), .Y(_182_) );
NOR2X1 NOR2X1_87 ( .A(_181_), .B(_182_), .Y(_183_) );
INVX1 INVX1_156 ( .A(_183_), .Y(_184_) );
NOR2X1 NOR2X1_88 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_185_) );
INVX1 INVX1_157 ( .A(_185_), .Y(_186_) );
NOR2X1 NOR2X1_89 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_187_) );
INVX1 INVX1_158 ( .A(_187_), .Y(_188_) );
NAND3X1 NAND3X1_85 ( .A(_186_), .B(_188_), .C(_179_), .Y(_189_) );
AND2X2 AND2X2_70 ( .A(_189_), .B(_184_), .Y(_190_) );
INVX1 INVX1_159 ( .A(_190_), .Y(w_C_31_) );
AND2X2 AND2X2_71 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_191_) );
INVX1 INVX1_160 ( .A(_191_), .Y(_192_) );
NAND3X1 NAND3X1_86 ( .A(_184_), .B(_192_), .C(_189_), .Y(_193_) );
OAI21X1 OAI21X1_71 ( .A(i_add2[31]), .B(i_add1[31]), .C(_193_), .Y(_194_) );
INVX1 INVX1_161 ( .A(_194_), .Y(w_C_32_) );
INVX1 INVX1_162 ( .A(i_add2[32]), .Y(_195_) );
INVX1 INVX1_163 ( .A(i_add1[32]), .Y(_196_) );
NOR2X1 NOR2X1_90 ( .A(_195_), .B(_196_), .Y(_197_) );
INVX1 INVX1_164 ( .A(_197_), .Y(_198_) );
NOR2X1 NOR2X1_91 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_199_) );
INVX1 INVX1_165 ( .A(_199_), .Y(_200_) );
NOR2X1 NOR2X1_92 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_201_) );
INVX1 INVX1_166 ( .A(_201_), .Y(_202_) );
NAND3X1 NAND3X1_87 ( .A(_200_), .B(_202_), .C(_193_), .Y(_203_) );
AND2X2 AND2X2_72 ( .A(_203_), .B(_198_), .Y(_204_) );
INVX1 INVX1_167 ( .A(_204_), .Y(w_C_33_) );
AND2X2 AND2X2_73 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_205_) );
INVX1 INVX1_168 ( .A(_205_), .Y(_206_) );
NAND3X1 NAND3X1_88 ( .A(_198_), .B(_206_), .C(_203_), .Y(_207_) );
OAI21X1 OAI21X1_72 ( .A(i_add2[33]), .B(i_add1[33]), .C(_207_), .Y(_208_) );
INVX1 INVX1_169 ( .A(_208_), .Y(w_C_34_) );
INVX1 INVX1_170 ( .A(i_add2[34]), .Y(_209_) );
INVX1 INVX1_171 ( .A(i_add1[34]), .Y(_210_) );
NOR2X1 NOR2X1_93 ( .A(_209_), .B(_210_), .Y(_211_) );
INVX1 INVX1_172 ( .A(_211_), .Y(_212_) );
NOR2X1 NOR2X1_94 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_213_) );
INVX1 INVX1_173 ( .A(_213_), .Y(_214_) );
NOR2X1 NOR2X1_95 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_215_) );
INVX1 INVX1_174 ( .A(_215_), .Y(_216_) );
NAND3X1 NAND3X1_89 ( .A(_214_), .B(_216_), .C(_207_), .Y(_217_) );
AND2X2 AND2X2_74 ( .A(_217_), .B(_212_), .Y(_218_) );
INVX1 INVX1_175 ( .A(_218_), .Y(w_C_35_) );
AND2X2 AND2X2_75 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_219_) );
INVX1 INVX1_176 ( .A(_219_), .Y(_220_) );
NAND3X1 NAND3X1_90 ( .A(_212_), .B(_220_), .C(_217_), .Y(_221_) );
OAI21X1 OAI21X1_73 ( .A(i_add2[35]), .B(i_add1[35]), .C(_221_), .Y(_222_) );
INVX1 INVX1_177 ( .A(_222_), .Y(w_C_36_) );
INVX1 INVX1_178 ( .A(i_add2[36]), .Y(_223_) );
INVX1 INVX1_179 ( .A(i_add1[36]), .Y(_224_) );
NOR2X1 NOR2X1_96 ( .A(_223_), .B(_224_), .Y(_225_) );
INVX1 INVX1_180 ( .A(_225_), .Y(_226_) );
NOR2X1 NOR2X1_97 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_227_) );
INVX1 INVX1_181 ( .A(_227_), .Y(_228_) );
NOR2X1 NOR2X1_98 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_229_) );
INVX1 INVX1_182 ( .A(_229_), .Y(_230_) );
BUFX2 BUFX2_1 ( .A(_278__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_278__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_278__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_278__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_278__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_278__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_278__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_278__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_278__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_278__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_278__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_278__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_278__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_278__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_278__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_278__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_278__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_278__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_278__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_278__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_278__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_278__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_278__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_278__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_278__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_278__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_278__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_278__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_278__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_278__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_278__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_278__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_278__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_278__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_278__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_278__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_278__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(_278__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .A(_278__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .A(_278__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .A(_278__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .A(_278__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .A(_278__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .A(_278__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .A(_278__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .A(_278__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .A(_278__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .A(w_C_47_), .Y(o_result[47]) );
INVX1 INVX1_183 ( .A(w_C_4_), .Y(_282_) );
OR2X2 OR2X2_53 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_283_) );
NAND2X1 NAND2X1_113 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_284_) );
NAND3X1 NAND3X1_91 ( .A(_282_), .B(_284_), .C(_283_), .Y(_285_) );
NOR2X1 NOR2X1_99 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_279_) );
AND2X2 AND2X2_76 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_280_) );
OAI21X1 OAI21X1_74 ( .A(_279_), .B(_280_), .C(w_C_4_), .Y(_281_) );
NAND2X1 NAND2X1_114 ( .A(_281_), .B(_285_), .Y(_278__4_) );
INVX1 INVX1_184 ( .A(w_C_5_), .Y(_289_) );
OR2X2 OR2X2_54 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_290_) );
NAND2X1 NAND2X1_115 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_291_) );
NAND3X1 NAND3X1_92 ( .A(_289_), .B(_291_), .C(_290_), .Y(_292_) );
NOR2X1 NOR2X1_100 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_286_) );
AND2X2 AND2X2_77 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_287_) );
OAI21X1 OAI21X1_75 ( .A(_286_), .B(_287_), .C(w_C_5_), .Y(_288_) );
NAND2X1 NAND2X1_116 ( .A(_288_), .B(_292_), .Y(_278__5_) );
INVX1 INVX1_185 ( .A(w_C_6_), .Y(_296_) );
OR2X2 OR2X2_55 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_297_) );
NAND2X1 NAND2X1_117 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_298_) );
BUFX2 BUFX2_49 ( .A(w_C_47_), .Y(_278__47_) );
BUFX2 BUFX2_50 ( .A(1'b0), .Y(w_C_0_) );
endmodule
