module cla_57bit (i_add1, i_add2, o_result);

input [56:0] i_add1;
input [56:0] i_add2;
output [57:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

NAND2X1 NAND2X1_1 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_324_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_325_) );
OAI21X1 OAI21X1_1 ( .A(_325_), .B(_323_), .C(_324_), .Y(w_C_54_) );
NAND2X1 NAND2X1_2 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_326_) );
INVX1 INVX1_1 ( .A(_325_), .Y(_327_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_328_) );
INVX1 INVX1_2 ( .A(_328_), .Y(_329_) );
NOR2X1 NOR2X1_3 ( .A(_311_), .B(_312_), .Y(_330_) );
INVX1 INVX1_3 ( .A(_330_), .Y(_331_) );
NAND3X1 NAND3X1_1 ( .A(_331_), .B(_319_), .C(_314_), .Y(_332_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_333_) );
INVX1 INVX1_4 ( .A(_333_), .Y(_334_) );
NAND3X1 NAND3X1_2 ( .A(_329_), .B(_334_), .C(_332_), .Y(_335_) );
NAND3X1 NAND3X1_3 ( .A(_321_), .B(_324_), .C(_335_), .Y(_336_) );
OR2X2 OR2X2_1 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_337_) );
NAND3X1 NAND3X1_4 ( .A(_327_), .B(_337_), .C(_336_), .Y(_338_) );
NAND2X1 NAND2X1_3 ( .A(_326_), .B(_338_), .Y(w_C_55_) );
OR2X2 OR2X2_2 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_339_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_340_) );
NAND3X1 NAND3X1_5 ( .A(_326_), .B(_340_), .C(_338_), .Y(_341_) );
AND2X2 AND2X2_1 ( .A(_341_), .B(_339_), .Y(w_C_56_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_342_) );
OR2X2 OR2X2_3 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_343_) );
NAND3X1 NAND3X1_6 ( .A(_339_), .B(_343_), .C(_341_), .Y(_344_) );
NAND2X1 NAND2X1_6 ( .A(_342_), .B(_344_), .Y(w_C_57_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_5 ( .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_8 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_9 ( .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_2 ( .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_6 ( .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_4 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_5 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_7 ( .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_11 ( .A(_4_), .B(_7_), .Y(w_C_3_) );
INVX1 INVX1_7 ( .A(i_add2[3]), .Y(_8_) );
INVX1 INVX1_8 ( .A(i_add1[3]), .Y(_9_) );
NAND2X1 NAND2X1_12 ( .A(_8_), .B(_9_), .Y(_10_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_11_) );
NAND3X1 NAND3X1_8 ( .A(_4_), .B(_11_), .C(_7_), .Y(_12_) );
AND2X2 AND2X2_2 ( .A(_12_), .B(_10_), .Y(w_C_4_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
OR2X2 OR2X2_6 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_14_) );
NAND3X1 NAND3X1_9 ( .A(_10_), .B(_14_), .C(_12_), .Y(_15_) );
NAND2X1 NAND2X1_15 ( .A(_13_), .B(_15_), .Y(w_C_5_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_16_) );
INVX1 INVX1_9 ( .A(_16_), .Y(_17_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_18_) );
NAND3X1 NAND3X1_10 ( .A(_13_), .B(_18_), .C(_15_), .Y(_19_) );
AND2X2 AND2X2_3 ( .A(_19_), .B(_17_), .Y(w_C_6_) );
INVX1 INVX1_10 ( .A(i_add2[6]), .Y(_20_) );
INVX1 INVX1_11 ( .A(i_add1[6]), .Y(_21_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_12 ( .A(_22_), .Y(_23_) );
NAND3X1 NAND3X1_11 ( .A(_17_), .B(_23_), .C(_19_), .Y(_24_) );
OAI21X1 OAI21X1_3 ( .A(_20_), .B(_21_), .C(_24_), .Y(w_C_7_) );
NOR2X1 NOR2X1_7 ( .A(_20_), .B(_21_), .Y(_25_) );
INVX1 INVX1_13 ( .A(_25_), .Y(_26_) );
AND2X2 AND2X2_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_27_) );
INVX1 INVX1_14 ( .A(_27_), .Y(_28_) );
NAND3X1 NAND3X1_12 ( .A(_26_), .B(_28_), .C(_24_), .Y(_29_) );
OAI21X1 OAI21X1_4 ( .A(i_add2[7]), .B(i_add1[7]), .C(_29_), .Y(_30_) );
INVX1 INVX1_15 ( .A(_30_), .Y(w_C_8_) );
INVX1 INVX1_16 ( .A(i_add2[8]), .Y(_31_) );
INVX1 INVX1_17 ( .A(i_add1[8]), .Y(_32_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_33_) );
INVX1 INVX1_18 ( .A(_33_), .Y(_34_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_35_) );
INVX1 INVX1_19 ( .A(_35_), .Y(_36_) );
NAND3X1 NAND3X1_13 ( .A(_34_), .B(_36_), .C(_29_), .Y(_37_) );
OAI21X1 OAI21X1_5 ( .A(_31_), .B(_32_), .C(_37_), .Y(w_C_9_) );
NOR2X1 NOR2X1_10 ( .A(_31_), .B(_32_), .Y(_38_) );
INVX1 INVX1_20 ( .A(_38_), .Y(_39_) );
AND2X2 AND2X2_5 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_40_) );
INVX1 INVX1_21 ( .A(_40_), .Y(_41_) );
NAND3X1 NAND3X1_14 ( .A(_39_), .B(_41_), .C(_37_), .Y(_42_) );
OAI21X1 OAI21X1_6 ( .A(i_add2[9]), .B(i_add1[9]), .C(_42_), .Y(_43_) );
INVX1 INVX1_22 ( .A(_43_), .Y(w_C_10_) );
INVX1 INVX1_23 ( .A(i_add2[10]), .Y(_44_) );
INVX1 INVX1_24 ( .A(i_add1[10]), .Y(_45_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_46_) );
INVX1 INVX1_25 ( .A(_46_), .Y(_47_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_48_) );
INVX1 INVX1_26 ( .A(_48_), .Y(_49_) );
NAND3X1 NAND3X1_15 ( .A(_47_), .B(_49_), .C(_42_), .Y(_50_) );
OAI21X1 OAI21X1_7 ( .A(_44_), .B(_45_), .C(_50_), .Y(w_C_11_) );
NOR2X1 NOR2X1_13 ( .A(_44_), .B(_45_), .Y(_51_) );
INVX1 INVX1_27 ( .A(_51_), .Y(_52_) );
AND2X2 AND2X2_6 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_53_) );
INVX1 INVX1_28 ( .A(_53_), .Y(_54_) );
NAND3X1 NAND3X1_16 ( .A(_52_), .B(_54_), .C(_50_), .Y(_55_) );
OAI21X1 OAI21X1_8 ( .A(i_add2[11]), .B(i_add1[11]), .C(_55_), .Y(_56_) );
INVX1 INVX1_29 ( .A(_56_), .Y(w_C_12_) );
INVX1 INVX1_30 ( .A(i_add2[12]), .Y(_57_) );
INVX1 INVX1_31 ( .A(i_add1[12]), .Y(_58_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_59_) );
INVX1 INVX1_32 ( .A(_59_), .Y(_60_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_61_) );
INVX1 INVX1_33 ( .A(_61_), .Y(_62_) );
NAND3X1 NAND3X1_17 ( .A(_60_), .B(_62_), .C(_55_), .Y(_63_) );
OAI21X1 OAI21X1_9 ( .A(_57_), .B(_58_), .C(_63_), .Y(w_C_13_) );
NOR2X1 NOR2X1_16 ( .A(_57_), .B(_58_), .Y(_64_) );
INVX1 INVX1_34 ( .A(_64_), .Y(_65_) );
AND2X2 AND2X2_7 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_66_) );
INVX1 INVX1_35 ( .A(_66_), .Y(_67_) );
NAND3X1 NAND3X1_18 ( .A(_65_), .B(_67_), .C(_63_), .Y(_68_) );
OAI21X1 OAI21X1_10 ( .A(i_add2[13]), .B(i_add1[13]), .C(_68_), .Y(_69_) );
INVX1 INVX1_36 ( .A(_69_), .Y(w_C_14_) );
INVX1 INVX1_37 ( .A(i_add2[14]), .Y(_70_) );
INVX1 INVX1_38 ( .A(i_add1[14]), .Y(_71_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_72_) );
INVX1 INVX1_39 ( .A(_72_), .Y(_73_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_74_) );
INVX1 INVX1_40 ( .A(_74_), .Y(_75_) );
NAND3X1 NAND3X1_19 ( .A(_73_), .B(_75_), .C(_68_), .Y(_76_) );
OAI21X1 OAI21X1_11 ( .A(_70_), .B(_71_), .C(_76_), .Y(w_C_15_) );
NOR2X1 NOR2X1_19 ( .A(_70_), .B(_71_), .Y(_77_) );
INVX1 INVX1_41 ( .A(_77_), .Y(_78_) );
AND2X2 AND2X2_8 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_79_) );
INVX1 INVX1_42 ( .A(_79_), .Y(_80_) );
NAND3X1 NAND3X1_20 ( .A(_78_), .B(_80_), .C(_76_), .Y(_81_) );
OAI21X1 OAI21X1_12 ( .A(i_add2[15]), .B(i_add1[15]), .C(_81_), .Y(_82_) );
INVX1 INVX1_43 ( .A(_82_), .Y(w_C_16_) );
INVX1 INVX1_44 ( .A(i_add2[16]), .Y(_83_) );
INVX1 INVX1_45 ( .A(i_add1[16]), .Y(_84_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_85_) );
INVX1 INVX1_46 ( .A(_85_), .Y(_86_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_87_) );
INVX1 INVX1_47 ( .A(_87_), .Y(_88_) );
NAND3X1 NAND3X1_21 ( .A(_86_), .B(_88_), .C(_81_), .Y(_89_) );
OAI21X1 OAI21X1_13 ( .A(_83_), .B(_84_), .C(_89_), .Y(w_C_17_) );
NOR2X1 NOR2X1_22 ( .A(_83_), .B(_84_), .Y(_90_) );
INVX1 INVX1_48 ( .A(_90_), .Y(_91_) );
AND2X2 AND2X2_9 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_92_) );
INVX1 INVX1_49 ( .A(_92_), .Y(_93_) );
NAND3X1 NAND3X1_22 ( .A(_91_), .B(_93_), .C(_89_), .Y(_94_) );
OAI21X1 OAI21X1_14 ( .A(i_add2[17]), .B(i_add1[17]), .C(_94_), .Y(_95_) );
INVX1 INVX1_50 ( .A(_95_), .Y(w_C_18_) );
INVX1 INVX1_51 ( .A(i_add2[18]), .Y(_96_) );
INVX1 INVX1_52 ( .A(i_add1[18]), .Y(_97_) );
NOR2X1 NOR2X1_23 ( .A(_96_), .B(_97_), .Y(_98_) );
INVX1 INVX1_53 ( .A(_98_), .Y(_99_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_100_) );
INVX1 INVX1_54 ( .A(_100_), .Y(_101_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_102_) );
INVX1 INVX1_55 ( .A(_102_), .Y(_103_) );
BUFX2 BUFX2_1 ( .A(_345__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_345__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_345__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_345__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_345__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_345__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_345__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_345__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_345__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_345__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_345__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_345__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_345__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_345__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_345__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_345__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_345__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_345__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_345__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_345__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_345__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_345__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_345__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_345__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_345__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_345__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_345__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_345__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_345__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_345__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_345__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_345__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_345__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_345__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_345__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_345__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_345__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(_345__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .A(_345__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .A(_345__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .A(_345__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .A(_345__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .A(_345__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .A(_345__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .A(_345__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .A(_345__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .A(_345__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .A(_345__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .A(_345__48_), .Y(o_result[48]) );
BUFX2 BUFX2_50 ( .A(_345__49_), .Y(o_result[49]) );
BUFX2 BUFX2_51 ( .A(_345__50_), .Y(o_result[50]) );
BUFX2 BUFX2_52 ( .A(_345__51_), .Y(o_result[51]) );
BUFX2 BUFX2_53 ( .A(_345__52_), .Y(o_result[52]) );
BUFX2 BUFX2_54 ( .A(_345__53_), .Y(o_result[53]) );
BUFX2 BUFX2_55 ( .A(_345__54_), .Y(o_result[54]) );
BUFX2 BUFX2_56 ( .A(_345__55_), .Y(o_result[55]) );
BUFX2 BUFX2_57 ( .A(_345__56_), .Y(o_result[56]) );
BUFX2 BUFX2_58 ( .A(w_C_57_), .Y(o_result[57]) );
INVX1 INVX1_56 ( .A(w_C_4_), .Y(_349_) );
OR2X2 OR2X2_7 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_350_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_351_) );
NAND3X1 NAND3X1_23 ( .A(_349_), .B(_351_), .C(_350_), .Y(_352_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_346_) );
AND2X2 AND2X2_10 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_347_) );
OAI21X1 OAI21X1_15 ( .A(_346_), .B(_347_), .C(w_C_4_), .Y(_348_) );
NAND2X1 NAND2X1_18 ( .A(_348_), .B(_352_), .Y(_345__4_) );
INVX1 INVX1_57 ( .A(w_C_5_), .Y(_356_) );
OR2X2 OR2X2_8 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_357_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_358_) );
NAND3X1 NAND3X1_24 ( .A(_356_), .B(_358_), .C(_357_), .Y(_359_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_353_) );
AND2X2 AND2X2_11 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_354_) );
OAI21X1 OAI21X1_16 ( .A(_353_), .B(_354_), .C(w_C_5_), .Y(_355_) );
NAND2X1 NAND2X1_20 ( .A(_355_), .B(_359_), .Y(_345__5_) );
INVX1 INVX1_58 ( .A(w_C_6_), .Y(_363_) );
OR2X2 OR2X2_9 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_364_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_365_) );
NAND3X1 NAND3X1_25 ( .A(_363_), .B(_365_), .C(_364_), .Y(_366_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_360_) );
AND2X2 AND2X2_12 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_361_) );
OAI21X1 OAI21X1_17 ( .A(_360_), .B(_361_), .C(w_C_6_), .Y(_362_) );
NAND2X1 NAND2X1_22 ( .A(_362_), .B(_366_), .Y(_345__6_) );
INVX1 INVX1_59 ( .A(w_C_7_), .Y(_370_) );
OR2X2 OR2X2_10 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_371_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_372_) );
NAND3X1 NAND3X1_26 ( .A(_370_), .B(_372_), .C(_371_), .Y(_373_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_367_) );
AND2X2 AND2X2_13 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_368_) );
OAI21X1 OAI21X1_18 ( .A(_367_), .B(_368_), .C(w_C_7_), .Y(_369_) );
NAND2X1 NAND2X1_24 ( .A(_369_), .B(_373_), .Y(_345__7_) );
INVX1 INVX1_60 ( .A(w_C_8_), .Y(_377_) );
OR2X2 OR2X2_11 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_378_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_379_) );
NAND3X1 NAND3X1_27 ( .A(_377_), .B(_379_), .C(_378_), .Y(_380_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_374_) );
AND2X2 AND2X2_14 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_375_) );
OAI21X1 OAI21X1_19 ( .A(_374_), .B(_375_), .C(w_C_8_), .Y(_376_) );
NAND2X1 NAND2X1_26 ( .A(_376_), .B(_380_), .Y(_345__8_) );
INVX1 INVX1_61 ( .A(w_C_9_), .Y(_384_) );
OR2X2 OR2X2_12 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_385_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_386_) );
NAND3X1 NAND3X1_28 ( .A(_384_), .B(_386_), .C(_385_), .Y(_387_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_381_) );
AND2X2 AND2X2_15 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_382_) );
OAI21X1 OAI21X1_20 ( .A(_381_), .B(_382_), .C(w_C_9_), .Y(_383_) );
NAND2X1 NAND2X1_28 ( .A(_383_), .B(_387_), .Y(_345__9_) );
INVX1 INVX1_62 ( .A(w_C_10_), .Y(_391_) );
OR2X2 OR2X2_13 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_392_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_393_) );
NAND3X1 NAND3X1_29 ( .A(_391_), .B(_393_), .C(_392_), .Y(_394_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_388_) );
AND2X2 AND2X2_16 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_389_) );
OAI21X1 OAI21X1_21 ( .A(_388_), .B(_389_), .C(w_C_10_), .Y(_390_) );
NAND2X1 NAND2X1_30 ( .A(_390_), .B(_394_), .Y(_345__10_) );
INVX1 INVX1_63 ( .A(w_C_11_), .Y(_398_) );
OR2X2 OR2X2_14 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_399_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_400_) );
NAND3X1 NAND3X1_30 ( .A(_398_), .B(_400_), .C(_399_), .Y(_401_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_395_) );
AND2X2 AND2X2_17 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_396_) );
OAI21X1 OAI21X1_22 ( .A(_395_), .B(_396_), .C(w_C_11_), .Y(_397_) );
NAND2X1 NAND2X1_32 ( .A(_397_), .B(_401_), .Y(_345__11_) );
INVX1 INVX1_64 ( .A(w_C_12_), .Y(_405_) );
OR2X2 OR2X2_15 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_406_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_407_) );
NAND3X1 NAND3X1_31 ( .A(_405_), .B(_407_), .C(_406_), .Y(_408_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_402_) );
AND2X2 AND2X2_18 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_403_) );
OAI21X1 OAI21X1_23 ( .A(_402_), .B(_403_), .C(w_C_12_), .Y(_404_) );
NAND2X1 NAND2X1_34 ( .A(_404_), .B(_408_), .Y(_345__12_) );
INVX1 INVX1_65 ( .A(w_C_13_), .Y(_412_) );
OR2X2 OR2X2_16 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_413_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_414_) );
NAND3X1 NAND3X1_32 ( .A(_412_), .B(_414_), .C(_413_), .Y(_415_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_409_) );
AND2X2 AND2X2_19 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_410_) );
OAI21X1 OAI21X1_24 ( .A(_409_), .B(_410_), .C(w_C_13_), .Y(_411_) );
NAND2X1 NAND2X1_36 ( .A(_411_), .B(_415_), .Y(_345__13_) );
INVX1 INVX1_66 ( .A(w_C_14_), .Y(_419_) );
OR2X2 OR2X2_17 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_420_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_421_) );
NAND3X1 NAND3X1_33 ( .A(_419_), .B(_421_), .C(_420_), .Y(_422_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_416_) );
AND2X2 AND2X2_20 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_417_) );
OAI21X1 OAI21X1_25 ( .A(_416_), .B(_417_), .C(w_C_14_), .Y(_418_) );
NAND2X1 NAND2X1_38 ( .A(_418_), .B(_422_), .Y(_345__14_) );
INVX1 INVX1_67 ( .A(w_C_15_), .Y(_426_) );
OR2X2 OR2X2_18 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_427_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_428_) );
NAND3X1 NAND3X1_34 ( .A(_426_), .B(_428_), .C(_427_), .Y(_429_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_423_) );
AND2X2 AND2X2_21 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_424_) );
OAI21X1 OAI21X1_26 ( .A(_423_), .B(_424_), .C(w_C_15_), .Y(_425_) );
NAND2X1 NAND2X1_40 ( .A(_425_), .B(_429_), .Y(_345__15_) );
INVX1 INVX1_68 ( .A(w_C_16_), .Y(_433_) );
OR2X2 OR2X2_19 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_434_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_435_) );
NAND3X1 NAND3X1_35 ( .A(_433_), .B(_435_), .C(_434_), .Y(_436_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_430_) );
AND2X2 AND2X2_22 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_431_) );
OAI21X1 OAI21X1_27 ( .A(_430_), .B(_431_), .C(w_C_16_), .Y(_432_) );
NAND2X1 NAND2X1_42 ( .A(_432_), .B(_436_), .Y(_345__16_) );
INVX1 INVX1_69 ( .A(w_C_17_), .Y(_440_) );
OR2X2 OR2X2_20 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_441_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_442_) );
NAND3X1 NAND3X1_36 ( .A(_440_), .B(_442_), .C(_441_), .Y(_443_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_437_) );
AND2X2 AND2X2_23 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_438_) );
OAI21X1 OAI21X1_28 ( .A(_437_), .B(_438_), .C(w_C_17_), .Y(_439_) );
NAND2X1 NAND2X1_44 ( .A(_439_), .B(_443_), .Y(_345__17_) );
INVX1 INVX1_70 ( .A(w_C_18_), .Y(_447_) );
OR2X2 OR2X2_21 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_448_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_449_) );
NAND3X1 NAND3X1_37 ( .A(_447_), .B(_449_), .C(_448_), .Y(_450_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_444_) );
AND2X2 AND2X2_24 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_445_) );
OAI21X1 OAI21X1_29 ( .A(_444_), .B(_445_), .C(w_C_18_), .Y(_446_) );
NAND2X1 NAND2X1_46 ( .A(_446_), .B(_450_), .Y(_345__18_) );
INVX1 INVX1_71 ( .A(w_C_19_), .Y(_454_) );
OR2X2 OR2X2_22 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_455_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_456_) );
NAND3X1 NAND3X1_38 ( .A(_454_), .B(_456_), .C(_455_), .Y(_457_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_451_) );
AND2X2 AND2X2_25 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_452_) );
OAI21X1 OAI21X1_30 ( .A(_451_), .B(_452_), .C(w_C_19_), .Y(_453_) );
NAND2X1 NAND2X1_48 ( .A(_453_), .B(_457_), .Y(_345__19_) );
INVX1 INVX1_72 ( .A(w_C_20_), .Y(_461_) );
OR2X2 OR2X2_23 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_462_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_463_) );
NAND3X1 NAND3X1_39 ( .A(_461_), .B(_463_), .C(_462_), .Y(_464_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_458_) );
AND2X2 AND2X2_26 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_459_) );
OAI21X1 OAI21X1_31 ( .A(_458_), .B(_459_), .C(w_C_20_), .Y(_460_) );
NAND2X1 NAND2X1_50 ( .A(_460_), .B(_464_), .Y(_345__20_) );
INVX1 INVX1_73 ( .A(w_C_21_), .Y(_468_) );
OR2X2 OR2X2_24 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_469_) );
NAND2X1 NAND2X1_51 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_470_) );
NAND3X1 NAND3X1_40 ( .A(_468_), .B(_470_), .C(_469_), .Y(_471_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_465_) );
AND2X2 AND2X2_27 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_466_) );
OAI21X1 OAI21X1_32 ( .A(_465_), .B(_466_), .C(w_C_21_), .Y(_467_) );
NAND2X1 NAND2X1_52 ( .A(_467_), .B(_471_), .Y(_345__21_) );
INVX1 INVX1_74 ( .A(w_C_22_), .Y(_475_) );
OR2X2 OR2X2_25 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_476_) );
NAND2X1 NAND2X1_53 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_477_) );
NAND3X1 NAND3X1_41 ( .A(_475_), .B(_477_), .C(_476_), .Y(_478_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_472_) );
AND2X2 AND2X2_28 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_473_) );
OAI21X1 OAI21X1_33 ( .A(_472_), .B(_473_), .C(w_C_22_), .Y(_474_) );
NAND2X1 NAND2X1_54 ( .A(_474_), .B(_478_), .Y(_345__22_) );
INVX1 INVX1_75 ( .A(w_C_23_), .Y(_482_) );
OR2X2 OR2X2_26 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_483_) );
NAND2X1 NAND2X1_55 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_484_) );
NAND3X1 NAND3X1_42 ( .A(_482_), .B(_484_), .C(_483_), .Y(_485_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_479_) );
AND2X2 AND2X2_29 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_480_) );
OAI21X1 OAI21X1_34 ( .A(_479_), .B(_480_), .C(w_C_23_), .Y(_481_) );
NAND2X1 NAND2X1_56 ( .A(_481_), .B(_485_), .Y(_345__23_) );
INVX1 INVX1_76 ( .A(w_C_24_), .Y(_489_) );
OR2X2 OR2X2_27 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_490_) );
NAND2X1 NAND2X1_57 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_491_) );
NAND3X1 NAND3X1_43 ( .A(_489_), .B(_491_), .C(_490_), .Y(_492_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_486_) );
AND2X2 AND2X2_30 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_487_) );
OAI21X1 OAI21X1_35 ( .A(_486_), .B(_487_), .C(w_C_24_), .Y(_488_) );
NAND2X1 NAND2X1_58 ( .A(_488_), .B(_492_), .Y(_345__24_) );
INVX1 INVX1_77 ( .A(w_C_25_), .Y(_496_) );
OR2X2 OR2X2_28 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_497_) );
NAND2X1 NAND2X1_59 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_498_) );
NAND3X1 NAND3X1_44 ( .A(_496_), .B(_498_), .C(_497_), .Y(_499_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_493_) );
AND2X2 AND2X2_31 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_494_) );
OAI21X1 OAI21X1_36 ( .A(_493_), .B(_494_), .C(w_C_25_), .Y(_495_) );
NAND2X1 NAND2X1_60 ( .A(_495_), .B(_499_), .Y(_345__25_) );
INVX1 INVX1_78 ( .A(w_C_26_), .Y(_503_) );
OR2X2 OR2X2_29 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_504_) );
NAND2X1 NAND2X1_61 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_505_) );
NAND3X1 NAND3X1_45 ( .A(_503_), .B(_505_), .C(_504_), .Y(_506_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_500_) );
AND2X2 AND2X2_32 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_501_) );
OAI21X1 OAI21X1_37 ( .A(_500_), .B(_501_), .C(w_C_26_), .Y(_502_) );
NAND2X1 NAND2X1_62 ( .A(_502_), .B(_506_), .Y(_345__26_) );
INVX1 INVX1_79 ( .A(w_C_27_), .Y(_510_) );
OR2X2 OR2X2_30 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_511_) );
NAND2X1 NAND2X1_63 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_512_) );
NAND3X1 NAND3X1_46 ( .A(_510_), .B(_512_), .C(_511_), .Y(_513_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_507_) );
AND2X2 AND2X2_33 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_508_) );
OAI21X1 OAI21X1_38 ( .A(_507_), .B(_508_), .C(w_C_27_), .Y(_509_) );
NAND2X1 NAND2X1_64 ( .A(_509_), .B(_513_), .Y(_345__27_) );
INVX1 INVX1_80 ( .A(w_C_28_), .Y(_517_) );
OR2X2 OR2X2_31 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_518_) );
NAND2X1 NAND2X1_65 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_519_) );
NAND3X1 NAND3X1_47 ( .A(_517_), .B(_519_), .C(_518_), .Y(_520_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_514_) );
AND2X2 AND2X2_34 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_515_) );
OAI21X1 OAI21X1_39 ( .A(_514_), .B(_515_), .C(w_C_28_), .Y(_516_) );
NAND2X1 NAND2X1_66 ( .A(_516_), .B(_520_), .Y(_345__28_) );
INVX1 INVX1_81 ( .A(w_C_29_), .Y(_524_) );
OR2X2 OR2X2_32 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_525_) );
NAND2X1 NAND2X1_67 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_526_) );
NAND3X1 NAND3X1_48 ( .A(_524_), .B(_526_), .C(_525_), .Y(_527_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_521_) );
AND2X2 AND2X2_35 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_522_) );
OAI21X1 OAI21X1_40 ( .A(_521_), .B(_522_), .C(w_C_29_), .Y(_523_) );
NAND2X1 NAND2X1_68 ( .A(_523_), .B(_527_), .Y(_345__29_) );
INVX1 INVX1_82 ( .A(w_C_30_), .Y(_531_) );
OR2X2 OR2X2_33 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_532_) );
NAND2X1 NAND2X1_69 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_533_) );
NAND3X1 NAND3X1_49 ( .A(_531_), .B(_533_), .C(_532_), .Y(_534_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_528_) );
AND2X2 AND2X2_36 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_529_) );
OAI21X1 OAI21X1_41 ( .A(_528_), .B(_529_), .C(w_C_30_), .Y(_530_) );
NAND2X1 NAND2X1_70 ( .A(_530_), .B(_534_), .Y(_345__30_) );
INVX1 INVX1_83 ( .A(w_C_31_), .Y(_538_) );
OR2X2 OR2X2_34 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_539_) );
NAND2X1 NAND2X1_71 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_540_) );
NAND3X1 NAND3X1_50 ( .A(_538_), .B(_540_), .C(_539_), .Y(_541_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_535_) );
AND2X2 AND2X2_37 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_536_) );
OAI21X1 OAI21X1_42 ( .A(_535_), .B(_536_), .C(w_C_31_), .Y(_537_) );
NAND2X1 NAND2X1_72 ( .A(_537_), .B(_541_), .Y(_345__31_) );
INVX1 INVX1_84 ( .A(w_C_32_), .Y(_545_) );
OR2X2 OR2X2_35 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_546_) );
NAND2X1 NAND2X1_73 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_547_) );
NAND3X1 NAND3X1_51 ( .A(_545_), .B(_547_), .C(_546_), .Y(_548_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_542_) );
AND2X2 AND2X2_38 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_543_) );
OAI21X1 OAI21X1_43 ( .A(_542_), .B(_543_), .C(w_C_32_), .Y(_544_) );
NAND2X1 NAND2X1_74 ( .A(_544_), .B(_548_), .Y(_345__32_) );
INVX1 INVX1_85 ( .A(w_C_33_), .Y(_552_) );
OR2X2 OR2X2_36 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_553_) );
NAND2X1 NAND2X1_75 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_554_) );
NAND3X1 NAND3X1_52 ( .A(_552_), .B(_554_), .C(_553_), .Y(_555_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_549_) );
AND2X2 AND2X2_39 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_550_) );
OAI21X1 OAI21X1_44 ( .A(_549_), .B(_550_), .C(w_C_33_), .Y(_551_) );
NAND2X1 NAND2X1_76 ( .A(_551_), .B(_555_), .Y(_345__33_) );
INVX1 INVX1_86 ( .A(w_C_34_), .Y(_559_) );
OR2X2 OR2X2_37 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_560_) );
NAND2X1 NAND2X1_77 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_561_) );
NAND3X1 NAND3X1_53 ( .A(_559_), .B(_561_), .C(_560_), .Y(_562_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_556_) );
AND2X2 AND2X2_40 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_557_) );
OAI21X1 OAI21X1_45 ( .A(_556_), .B(_557_), .C(w_C_34_), .Y(_558_) );
NAND2X1 NAND2X1_78 ( .A(_558_), .B(_562_), .Y(_345__34_) );
INVX1 INVX1_87 ( .A(w_C_35_), .Y(_566_) );
OR2X2 OR2X2_38 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_567_) );
NAND2X1 NAND2X1_79 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_568_) );
NAND3X1 NAND3X1_54 ( .A(_566_), .B(_568_), .C(_567_), .Y(_569_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_563_) );
AND2X2 AND2X2_41 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_564_) );
OAI21X1 OAI21X1_46 ( .A(_563_), .B(_564_), .C(w_C_35_), .Y(_565_) );
NAND2X1 NAND2X1_80 ( .A(_565_), .B(_569_), .Y(_345__35_) );
INVX1 INVX1_88 ( .A(w_C_36_), .Y(_573_) );
OR2X2 OR2X2_39 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_574_) );
NAND2X1 NAND2X1_81 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_575_) );
NAND3X1 NAND3X1_55 ( .A(_573_), .B(_575_), .C(_574_), .Y(_576_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_570_) );
AND2X2 AND2X2_42 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_571_) );
OAI21X1 OAI21X1_47 ( .A(_570_), .B(_571_), .C(w_C_36_), .Y(_572_) );
NAND2X1 NAND2X1_82 ( .A(_572_), .B(_576_), .Y(_345__36_) );
INVX1 INVX1_89 ( .A(w_C_37_), .Y(_580_) );
OR2X2 OR2X2_40 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_581_) );
NAND2X1 NAND2X1_83 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_582_) );
NAND3X1 NAND3X1_56 ( .A(_580_), .B(_582_), .C(_581_), .Y(_583_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_577_) );
AND2X2 AND2X2_43 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_578_) );
OAI21X1 OAI21X1_48 ( .A(_577_), .B(_578_), .C(w_C_37_), .Y(_579_) );
NAND2X1 NAND2X1_84 ( .A(_579_), .B(_583_), .Y(_345__37_) );
INVX1 INVX1_90 ( .A(w_C_38_), .Y(_587_) );
OR2X2 OR2X2_41 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_588_) );
NAND2X1 NAND2X1_85 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_589_) );
NAND3X1 NAND3X1_57 ( .A(_587_), .B(_589_), .C(_588_), .Y(_590_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_584_) );
AND2X2 AND2X2_44 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_585_) );
OAI21X1 OAI21X1_49 ( .A(_584_), .B(_585_), .C(w_C_38_), .Y(_586_) );
NAND2X1 NAND2X1_86 ( .A(_586_), .B(_590_), .Y(_345__38_) );
INVX1 INVX1_91 ( .A(w_C_39_), .Y(_594_) );
OR2X2 OR2X2_42 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_595_) );
NAND2X1 NAND2X1_87 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_596_) );
NAND3X1 NAND3X1_58 ( .A(_594_), .B(_596_), .C(_595_), .Y(_597_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_591_) );
AND2X2 AND2X2_45 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_592_) );
OAI21X1 OAI21X1_50 ( .A(_591_), .B(_592_), .C(w_C_39_), .Y(_593_) );
NAND2X1 NAND2X1_88 ( .A(_593_), .B(_597_), .Y(_345__39_) );
INVX1 INVX1_92 ( .A(w_C_40_), .Y(_601_) );
OR2X2 OR2X2_43 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_602_) );
NAND2X1 NAND2X1_89 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_603_) );
NAND3X1 NAND3X1_59 ( .A(_601_), .B(_603_), .C(_602_), .Y(_604_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_598_) );
AND2X2 AND2X2_46 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_599_) );
OAI21X1 OAI21X1_51 ( .A(_598_), .B(_599_), .C(w_C_40_), .Y(_600_) );
NAND2X1 NAND2X1_90 ( .A(_600_), .B(_604_), .Y(_345__40_) );
INVX1 INVX1_93 ( .A(w_C_41_), .Y(_608_) );
OR2X2 OR2X2_44 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_609_) );
NAND2X1 NAND2X1_91 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_610_) );
NAND3X1 NAND3X1_60 ( .A(_608_), .B(_610_), .C(_609_), .Y(_611_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_605_) );
AND2X2 AND2X2_47 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_606_) );
OAI21X1 OAI21X1_52 ( .A(_605_), .B(_606_), .C(w_C_41_), .Y(_607_) );
NAND2X1 NAND2X1_92 ( .A(_607_), .B(_611_), .Y(_345__41_) );
INVX1 INVX1_94 ( .A(w_C_42_), .Y(_615_) );
OR2X2 OR2X2_45 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_616_) );
NAND2X1 NAND2X1_93 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_617_) );
NAND3X1 NAND3X1_61 ( .A(_615_), .B(_617_), .C(_616_), .Y(_618_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_612_) );
AND2X2 AND2X2_48 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_613_) );
OAI21X1 OAI21X1_53 ( .A(_612_), .B(_613_), .C(w_C_42_), .Y(_614_) );
NAND2X1 NAND2X1_94 ( .A(_614_), .B(_618_), .Y(_345__42_) );
INVX1 INVX1_95 ( .A(w_C_43_), .Y(_622_) );
OR2X2 OR2X2_46 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_623_) );
NAND2X1 NAND2X1_95 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_624_) );
NAND3X1 NAND3X1_62 ( .A(_622_), .B(_624_), .C(_623_), .Y(_625_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_619_) );
AND2X2 AND2X2_49 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_620_) );
OAI21X1 OAI21X1_54 ( .A(_619_), .B(_620_), .C(w_C_43_), .Y(_621_) );
NAND2X1 NAND2X1_96 ( .A(_621_), .B(_625_), .Y(_345__43_) );
INVX1 INVX1_96 ( .A(w_C_44_), .Y(_629_) );
OR2X2 OR2X2_47 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_630_) );
NAND2X1 NAND2X1_97 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_631_) );
NAND3X1 NAND3X1_63 ( .A(_629_), .B(_631_), .C(_630_), .Y(_632_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_626_) );
AND2X2 AND2X2_50 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_627_) );
OAI21X1 OAI21X1_55 ( .A(_626_), .B(_627_), .C(w_C_44_), .Y(_628_) );
NAND2X1 NAND2X1_98 ( .A(_628_), .B(_632_), .Y(_345__44_) );
INVX1 INVX1_97 ( .A(w_C_45_), .Y(_636_) );
OR2X2 OR2X2_48 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_637_) );
NAND2X1 NAND2X1_99 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_638_) );
NAND3X1 NAND3X1_64 ( .A(_636_), .B(_638_), .C(_637_), .Y(_639_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_633_) );
AND2X2 AND2X2_51 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_634_) );
OAI21X1 OAI21X1_56 ( .A(_633_), .B(_634_), .C(w_C_45_), .Y(_635_) );
NAND2X1 NAND2X1_100 ( .A(_635_), .B(_639_), .Y(_345__45_) );
INVX1 INVX1_98 ( .A(w_C_46_), .Y(_643_) );
OR2X2 OR2X2_49 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_644_) );
NAND2X1 NAND2X1_101 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_645_) );
NAND3X1 NAND3X1_65 ( .A(_643_), .B(_645_), .C(_644_), .Y(_646_) );
NOR2X1 NOR2X1_68 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_640_) );
AND2X2 AND2X2_52 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_641_) );
OAI21X1 OAI21X1_57 ( .A(_640_), .B(_641_), .C(w_C_46_), .Y(_642_) );
NAND2X1 NAND2X1_102 ( .A(_642_), .B(_646_), .Y(_345__46_) );
INVX1 INVX1_99 ( .A(w_C_47_), .Y(_650_) );
OR2X2 OR2X2_50 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_651_) );
NAND2X1 NAND2X1_103 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_652_) );
NAND3X1 NAND3X1_66 ( .A(_650_), .B(_652_), .C(_651_), .Y(_653_) );
NOR2X1 NOR2X1_69 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_647_) );
AND2X2 AND2X2_53 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_648_) );
OAI21X1 OAI21X1_58 ( .A(_647_), .B(_648_), .C(w_C_47_), .Y(_649_) );
NAND2X1 NAND2X1_104 ( .A(_649_), .B(_653_), .Y(_345__47_) );
INVX1 INVX1_100 ( .A(w_C_48_), .Y(_657_) );
OR2X2 OR2X2_51 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_658_) );
NAND2X1 NAND2X1_105 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_659_) );
NAND3X1 NAND3X1_67 ( .A(_657_), .B(_659_), .C(_658_), .Y(_660_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_654_) );
AND2X2 AND2X2_54 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_655_) );
OAI21X1 OAI21X1_59 ( .A(_654_), .B(_655_), .C(w_C_48_), .Y(_656_) );
NAND2X1 NAND2X1_106 ( .A(_656_), .B(_660_), .Y(_345__48_) );
INVX1 INVX1_101 ( .A(w_C_49_), .Y(_664_) );
OR2X2 OR2X2_52 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_665_) );
NAND2X1 NAND2X1_107 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_666_) );
NAND3X1 NAND3X1_68 ( .A(_664_), .B(_666_), .C(_665_), .Y(_667_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_661_) );
AND2X2 AND2X2_55 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_662_) );
OAI21X1 OAI21X1_60 ( .A(_661_), .B(_662_), .C(w_C_49_), .Y(_663_) );
NAND2X1 NAND2X1_108 ( .A(_663_), .B(_667_), .Y(_345__49_) );
INVX1 INVX1_102 ( .A(w_C_50_), .Y(_671_) );
OR2X2 OR2X2_53 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_672_) );
NAND2X1 NAND2X1_109 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_673_) );
NAND3X1 NAND3X1_69 ( .A(_671_), .B(_673_), .C(_672_), .Y(_674_) );
NOR2X1 NOR2X1_72 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_668_) );
AND2X2 AND2X2_56 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_669_) );
OAI21X1 OAI21X1_61 ( .A(_668_), .B(_669_), .C(w_C_50_), .Y(_670_) );
NAND2X1 NAND2X1_110 ( .A(_670_), .B(_674_), .Y(_345__50_) );
INVX1 INVX1_103 ( .A(w_C_51_), .Y(_678_) );
OR2X2 OR2X2_54 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_679_) );
NAND2X1 NAND2X1_111 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_680_) );
NAND3X1 NAND3X1_70 ( .A(_678_), .B(_680_), .C(_679_), .Y(_681_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_675_) );
AND2X2 AND2X2_57 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_676_) );
OAI21X1 OAI21X1_62 ( .A(_675_), .B(_676_), .C(w_C_51_), .Y(_677_) );
NAND2X1 NAND2X1_112 ( .A(_677_), .B(_681_), .Y(_345__51_) );
INVX1 INVX1_104 ( .A(w_C_52_), .Y(_685_) );
OR2X2 OR2X2_55 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_686_) );
NAND2X1 NAND2X1_113 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_687_) );
NAND3X1 NAND3X1_71 ( .A(_685_), .B(_687_), .C(_686_), .Y(_688_) );
NOR2X1 NOR2X1_74 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_682_) );
AND2X2 AND2X2_58 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_683_) );
OAI21X1 OAI21X1_63 ( .A(_682_), .B(_683_), .C(w_C_52_), .Y(_684_) );
NAND2X1 NAND2X1_114 ( .A(_684_), .B(_688_), .Y(_345__52_) );
INVX1 INVX1_105 ( .A(w_C_53_), .Y(_692_) );
OR2X2 OR2X2_56 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_693_) );
NAND2X1 NAND2X1_115 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_694_) );
NAND3X1 NAND3X1_72 ( .A(_692_), .B(_694_), .C(_693_), .Y(_695_) );
NOR2X1 NOR2X1_75 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_689_) );
AND2X2 AND2X2_59 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_690_) );
OAI21X1 OAI21X1_64 ( .A(_689_), .B(_690_), .C(w_C_53_), .Y(_691_) );
NAND2X1 NAND2X1_116 ( .A(_691_), .B(_695_), .Y(_345__53_) );
INVX1 INVX1_106 ( .A(w_C_54_), .Y(_699_) );
OR2X2 OR2X2_57 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_700_) );
NAND2X1 NAND2X1_117 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_701_) );
NAND3X1 NAND3X1_73 ( .A(_699_), .B(_701_), .C(_700_), .Y(_702_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_696_) );
AND2X2 AND2X2_60 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_697_) );
OAI21X1 OAI21X1_65 ( .A(_696_), .B(_697_), .C(w_C_54_), .Y(_698_) );
NAND2X1 NAND2X1_118 ( .A(_698_), .B(_702_), .Y(_345__54_) );
INVX1 INVX1_107 ( .A(w_C_55_), .Y(_706_) );
OR2X2 OR2X2_58 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_707_) );
NAND2X1 NAND2X1_119 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_708_) );
NAND3X1 NAND3X1_74 ( .A(_706_), .B(_708_), .C(_707_), .Y(_709_) );
NOR2X1 NOR2X1_77 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_703_) );
AND2X2 AND2X2_61 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_704_) );
OAI21X1 OAI21X1_66 ( .A(_703_), .B(_704_), .C(w_C_55_), .Y(_705_) );
NAND2X1 NAND2X1_120 ( .A(_705_), .B(_709_), .Y(_345__55_) );
INVX1 INVX1_108 ( .A(w_C_56_), .Y(_713_) );
OR2X2 OR2X2_59 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_714_) );
NAND2X1 NAND2X1_121 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_715_) );
NAND3X1 NAND3X1_75 ( .A(_713_), .B(_715_), .C(_714_), .Y(_716_) );
NOR2X1 NOR2X1_78 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_710_) );
AND2X2 AND2X2_62 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_711_) );
OAI21X1 OAI21X1_67 ( .A(_710_), .B(_711_), .C(w_C_56_), .Y(_712_) );
NAND2X1 NAND2X1_122 ( .A(_712_), .B(_716_), .Y(_345__56_) );
INVX1 INVX1_109 ( .A(gnd), .Y(_720_) );
OR2X2 OR2X2_60 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_721_) );
NAND2X1 NAND2X1_123 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_722_) );
NAND3X1 NAND3X1_76 ( .A(_720_), .B(_722_), .C(_721_), .Y(_723_) );
NOR2X1 NOR2X1_79 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_717_) );
AND2X2 AND2X2_63 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_718_) );
OAI21X1 OAI21X1_68 ( .A(_717_), .B(_718_), .C(gnd), .Y(_719_) );
NAND2X1 NAND2X1_124 ( .A(_719_), .B(_723_), .Y(_345__0_) );
INVX1 INVX1_110 ( .A(w_C_1_), .Y(_727_) );
OR2X2 OR2X2_61 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_728_) );
NAND2X1 NAND2X1_125 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_729_) );
NAND3X1 NAND3X1_77 ( .A(_727_), .B(_729_), .C(_728_), .Y(_730_) );
NOR2X1 NOR2X1_80 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_724_) );
AND2X2 AND2X2_64 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_725_) );
OAI21X1 OAI21X1_69 ( .A(_724_), .B(_725_), .C(w_C_1_), .Y(_726_) );
NAND2X1 NAND2X1_126 ( .A(_726_), .B(_730_), .Y(_345__1_) );
INVX1 INVX1_111 ( .A(w_C_2_), .Y(_734_) );
OR2X2 OR2X2_62 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_735_) );
NAND2X1 NAND2X1_127 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_736_) );
NAND3X1 NAND3X1_78 ( .A(_734_), .B(_736_), .C(_735_), .Y(_737_) );
NOR2X1 NOR2X1_81 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_731_) );
AND2X2 AND2X2_65 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_732_) );
OAI21X1 OAI21X1_70 ( .A(_731_), .B(_732_), .C(w_C_2_), .Y(_733_) );
NAND2X1 NAND2X1_128 ( .A(_733_), .B(_737_), .Y(_345__2_) );
INVX1 INVX1_112 ( .A(w_C_3_), .Y(_741_) );
OR2X2 OR2X2_63 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_742_) );
NAND2X1 NAND2X1_129 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_743_) );
NAND3X1 NAND3X1_79 ( .A(_741_), .B(_743_), .C(_742_), .Y(_744_) );
NOR2X1 NOR2X1_82 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_738_) );
AND2X2 AND2X2_66 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_739_) );
OAI21X1 OAI21X1_71 ( .A(_738_), .B(_739_), .C(w_C_3_), .Y(_740_) );
NAND2X1 NAND2X1_130 ( .A(_740_), .B(_744_), .Y(_345__3_) );
NAND3X1 NAND3X1_80 ( .A(_101_), .B(_103_), .C(_94_), .Y(_104_) );
AND2X2 AND2X2_67 ( .A(_104_), .B(_99_), .Y(_105_) );
INVX1 INVX1_113 ( .A(_105_), .Y(w_C_19_) );
AND2X2 AND2X2_68 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_106_) );
INVX1 INVX1_114 ( .A(_106_), .Y(_107_) );
NAND3X1 NAND3X1_81 ( .A(_99_), .B(_107_), .C(_104_), .Y(_108_) );
OAI21X1 OAI21X1_72 ( .A(i_add2[19]), .B(i_add1[19]), .C(_108_), .Y(_109_) );
INVX1 INVX1_115 ( .A(_109_), .Y(w_C_20_) );
INVX1 INVX1_116 ( .A(i_add2[20]), .Y(_110_) );
INVX1 INVX1_117 ( .A(i_add1[20]), .Y(_111_) );
NOR2X1 NOR2X1_83 ( .A(_110_), .B(_111_), .Y(_112_) );
INVX1 INVX1_118 ( .A(_112_), .Y(_113_) );
NOR2X1 NOR2X1_84 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_114_) );
INVX1 INVX1_119 ( .A(_114_), .Y(_115_) );
NOR2X1 NOR2X1_85 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_116_) );
INVX1 INVX1_120 ( .A(_116_), .Y(_117_) );
NAND3X1 NAND3X1_82 ( .A(_115_), .B(_117_), .C(_108_), .Y(_118_) );
AND2X2 AND2X2_69 ( .A(_118_), .B(_113_), .Y(_119_) );
INVX1 INVX1_121 ( .A(_119_), .Y(w_C_21_) );
AND2X2 AND2X2_70 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_120_) );
INVX1 INVX1_122 ( .A(_120_), .Y(_121_) );
NAND3X1 NAND3X1_83 ( .A(_113_), .B(_121_), .C(_118_), .Y(_122_) );
OAI21X1 OAI21X1_73 ( .A(i_add2[21]), .B(i_add1[21]), .C(_122_), .Y(_123_) );
INVX1 INVX1_123 ( .A(_123_), .Y(w_C_22_) );
INVX1 INVX1_124 ( .A(i_add2[22]), .Y(_124_) );
INVX1 INVX1_125 ( .A(i_add1[22]), .Y(_125_) );
NOR2X1 NOR2X1_86 ( .A(_124_), .B(_125_), .Y(_126_) );
INVX1 INVX1_126 ( .A(_126_), .Y(_127_) );
NOR2X1 NOR2X1_87 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_128_) );
INVX1 INVX1_127 ( .A(_128_), .Y(_129_) );
NOR2X1 NOR2X1_88 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_130_) );
INVX1 INVX1_128 ( .A(_130_), .Y(_131_) );
NAND3X1 NAND3X1_84 ( .A(_129_), .B(_131_), .C(_122_), .Y(_132_) );
AND2X2 AND2X2_71 ( .A(_132_), .B(_127_), .Y(_133_) );
INVX1 INVX1_129 ( .A(_133_), .Y(w_C_23_) );
AND2X2 AND2X2_72 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_134_) );
INVX1 INVX1_130 ( .A(_134_), .Y(_135_) );
NAND3X1 NAND3X1_85 ( .A(_127_), .B(_135_), .C(_132_), .Y(_136_) );
OAI21X1 OAI21X1_74 ( .A(i_add2[23]), .B(i_add1[23]), .C(_136_), .Y(_137_) );
INVX1 INVX1_131 ( .A(_137_), .Y(w_C_24_) );
INVX1 INVX1_132 ( .A(i_add2[24]), .Y(_138_) );
INVX1 INVX1_133 ( .A(i_add1[24]), .Y(_139_) );
NOR2X1 NOR2X1_89 ( .A(_138_), .B(_139_), .Y(_140_) );
INVX1 INVX1_134 ( .A(_140_), .Y(_141_) );
NOR2X1 NOR2X1_90 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_142_) );
INVX1 INVX1_135 ( .A(_142_), .Y(_143_) );
NOR2X1 NOR2X1_91 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_144_) );
INVX1 INVX1_136 ( .A(_144_), .Y(_145_) );
NAND3X1 NAND3X1_86 ( .A(_143_), .B(_145_), .C(_136_), .Y(_146_) );
AND2X2 AND2X2_73 ( .A(_146_), .B(_141_), .Y(_147_) );
INVX1 INVX1_137 ( .A(_147_), .Y(w_C_25_) );
AND2X2 AND2X2_74 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_148_) );
INVX1 INVX1_138 ( .A(_148_), .Y(_149_) );
NAND3X1 NAND3X1_87 ( .A(_141_), .B(_149_), .C(_146_), .Y(_150_) );
OAI21X1 OAI21X1_75 ( .A(i_add2[25]), .B(i_add1[25]), .C(_150_), .Y(_151_) );
INVX1 INVX1_139 ( .A(_151_), .Y(w_C_26_) );
INVX1 INVX1_140 ( .A(i_add2[26]), .Y(_152_) );
INVX1 INVX1_141 ( .A(i_add1[26]), .Y(_153_) );
NOR2X1 NOR2X1_92 ( .A(_152_), .B(_153_), .Y(_154_) );
INVX1 INVX1_142 ( .A(_154_), .Y(_155_) );
NOR2X1 NOR2X1_93 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_156_) );
INVX1 INVX1_143 ( .A(_156_), .Y(_157_) );
NOR2X1 NOR2X1_94 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_158_) );
INVX1 INVX1_144 ( .A(_158_), .Y(_159_) );
NAND3X1 NAND3X1_88 ( .A(_157_), .B(_159_), .C(_150_), .Y(_160_) );
AND2X2 AND2X2_75 ( .A(_160_), .B(_155_), .Y(_161_) );
INVX1 INVX1_145 ( .A(_161_), .Y(w_C_27_) );
AND2X2 AND2X2_76 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_162_) );
INVX1 INVX1_146 ( .A(_162_), .Y(_163_) );
NAND3X1 NAND3X1_89 ( .A(_155_), .B(_163_), .C(_160_), .Y(_164_) );
OAI21X1 OAI21X1_76 ( .A(i_add2[27]), .B(i_add1[27]), .C(_164_), .Y(_165_) );
INVX1 INVX1_147 ( .A(_165_), .Y(w_C_28_) );
INVX1 INVX1_148 ( .A(i_add2[28]), .Y(_166_) );
INVX1 INVX1_149 ( .A(i_add1[28]), .Y(_167_) );
NOR2X1 NOR2X1_95 ( .A(_166_), .B(_167_), .Y(_168_) );
INVX1 INVX1_150 ( .A(_168_), .Y(_169_) );
NOR2X1 NOR2X1_96 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_170_) );
INVX1 INVX1_151 ( .A(_170_), .Y(_171_) );
NOR2X1 NOR2X1_97 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_172_) );
INVX1 INVX1_152 ( .A(_172_), .Y(_173_) );
NAND3X1 NAND3X1_90 ( .A(_171_), .B(_173_), .C(_164_), .Y(_174_) );
AND2X2 AND2X2_77 ( .A(_174_), .B(_169_), .Y(_175_) );
INVX1 INVX1_153 ( .A(_175_), .Y(w_C_29_) );
AND2X2 AND2X2_78 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_176_) );
INVX1 INVX1_154 ( .A(_176_), .Y(_177_) );
NAND3X1 NAND3X1_91 ( .A(_169_), .B(_177_), .C(_174_), .Y(_178_) );
OAI21X1 OAI21X1_77 ( .A(i_add2[29]), .B(i_add1[29]), .C(_178_), .Y(_179_) );
INVX1 INVX1_155 ( .A(_179_), .Y(w_C_30_) );
INVX1 INVX1_156 ( .A(i_add2[30]), .Y(_180_) );
INVX1 INVX1_157 ( .A(i_add1[30]), .Y(_181_) );
NOR2X1 NOR2X1_98 ( .A(_180_), .B(_181_), .Y(_182_) );
INVX1 INVX1_158 ( .A(_182_), .Y(_183_) );
NOR2X1 NOR2X1_99 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_184_) );
INVX1 INVX1_159 ( .A(_184_), .Y(_185_) );
NOR2X1 NOR2X1_100 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_186_) );
INVX1 INVX1_160 ( .A(_186_), .Y(_187_) );
NAND3X1 NAND3X1_92 ( .A(_185_), .B(_187_), .C(_178_), .Y(_188_) );
AND2X2 AND2X2_79 ( .A(_188_), .B(_183_), .Y(_189_) );
INVX1 INVX1_161 ( .A(_189_), .Y(w_C_31_) );
AND2X2 AND2X2_80 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_190_) );
INVX1 INVX1_162 ( .A(_190_), .Y(_191_) );
NAND3X1 NAND3X1_93 ( .A(_183_), .B(_191_), .C(_188_), .Y(_192_) );
OAI21X1 OAI21X1_78 ( .A(i_add2[31]), .B(i_add1[31]), .C(_192_), .Y(_193_) );
INVX1 INVX1_163 ( .A(_193_), .Y(w_C_32_) );
INVX1 INVX1_164 ( .A(i_add2[32]), .Y(_194_) );
INVX1 INVX1_165 ( .A(i_add1[32]), .Y(_195_) );
NOR2X1 NOR2X1_101 ( .A(_194_), .B(_195_), .Y(_196_) );
INVX1 INVX1_166 ( .A(_196_), .Y(_197_) );
NOR2X1 NOR2X1_102 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_198_) );
INVX1 INVX1_167 ( .A(_198_), .Y(_199_) );
NOR2X1 NOR2X1_103 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_200_) );
INVX1 INVX1_168 ( .A(_200_), .Y(_201_) );
NAND3X1 NAND3X1_94 ( .A(_199_), .B(_201_), .C(_192_), .Y(_202_) );
AND2X2 AND2X2_81 ( .A(_202_), .B(_197_), .Y(_203_) );
INVX1 INVX1_169 ( .A(_203_), .Y(w_C_33_) );
AND2X2 AND2X2_82 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_204_) );
INVX1 INVX1_170 ( .A(_204_), .Y(_205_) );
NAND3X1 NAND3X1_95 ( .A(_197_), .B(_205_), .C(_202_), .Y(_206_) );
OAI21X1 OAI21X1_79 ( .A(i_add2[33]), .B(i_add1[33]), .C(_206_), .Y(_207_) );
INVX1 INVX1_171 ( .A(_207_), .Y(w_C_34_) );
INVX1 INVX1_172 ( .A(i_add2[34]), .Y(_208_) );
INVX1 INVX1_173 ( .A(i_add1[34]), .Y(_209_) );
NOR2X1 NOR2X1_104 ( .A(_208_), .B(_209_), .Y(_210_) );
INVX1 INVX1_174 ( .A(_210_), .Y(_211_) );
NOR2X1 NOR2X1_105 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_212_) );
INVX1 INVX1_175 ( .A(_212_), .Y(_213_) );
NOR2X1 NOR2X1_106 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_214_) );
INVX1 INVX1_176 ( .A(_214_), .Y(_215_) );
NAND3X1 NAND3X1_96 ( .A(_213_), .B(_215_), .C(_206_), .Y(_216_) );
AND2X2 AND2X2_83 ( .A(_216_), .B(_211_), .Y(_217_) );
INVX1 INVX1_177 ( .A(_217_), .Y(w_C_35_) );
AND2X2 AND2X2_84 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_218_) );
INVX1 INVX1_178 ( .A(_218_), .Y(_219_) );
NAND3X1 NAND3X1_97 ( .A(_211_), .B(_219_), .C(_216_), .Y(_220_) );
OAI21X1 OAI21X1_80 ( .A(i_add2[35]), .B(i_add1[35]), .C(_220_), .Y(_221_) );
INVX1 INVX1_179 ( .A(_221_), .Y(w_C_36_) );
INVX1 INVX1_180 ( .A(i_add2[36]), .Y(_222_) );
INVX1 INVX1_181 ( .A(i_add1[36]), .Y(_223_) );
NOR2X1 NOR2X1_107 ( .A(_222_), .B(_223_), .Y(_224_) );
INVX1 INVX1_182 ( .A(_224_), .Y(_225_) );
NOR2X1 NOR2X1_108 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_226_) );
INVX1 INVX1_183 ( .A(_226_), .Y(_227_) );
NOR2X1 NOR2X1_109 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_228_) );
INVX1 INVX1_184 ( .A(_228_), .Y(_229_) );
NAND3X1 NAND3X1_98 ( .A(_227_), .B(_229_), .C(_220_), .Y(_230_) );
AND2X2 AND2X2_85 ( .A(_230_), .B(_225_), .Y(_231_) );
INVX1 INVX1_185 ( .A(_231_), .Y(w_C_37_) );
AND2X2 AND2X2_86 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_232_) );
INVX1 INVX1_186 ( .A(_232_), .Y(_233_) );
NAND3X1 NAND3X1_99 ( .A(_225_), .B(_233_), .C(_230_), .Y(_234_) );
OAI21X1 OAI21X1_81 ( .A(i_add2[37]), .B(i_add1[37]), .C(_234_), .Y(_235_) );
INVX1 INVX1_187 ( .A(_235_), .Y(w_C_38_) );
INVX1 INVX1_188 ( .A(i_add2[38]), .Y(_236_) );
INVX1 INVX1_189 ( .A(i_add1[38]), .Y(_237_) );
NOR2X1 NOR2X1_110 ( .A(_236_), .B(_237_), .Y(_238_) );
INVX1 INVX1_190 ( .A(_238_), .Y(_239_) );
NOR2X1 NOR2X1_111 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_240_) );
INVX1 INVX1_191 ( .A(_240_), .Y(_241_) );
NOR2X1 NOR2X1_112 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_242_) );
INVX1 INVX1_192 ( .A(_242_), .Y(_243_) );
NAND3X1 NAND3X1_100 ( .A(_241_), .B(_243_), .C(_234_), .Y(_244_) );
AND2X2 AND2X2_87 ( .A(_244_), .B(_239_), .Y(_245_) );
INVX1 INVX1_193 ( .A(_245_), .Y(w_C_39_) );
AND2X2 AND2X2_88 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_246_) );
INVX1 INVX1_194 ( .A(_246_), .Y(_247_) );
NAND3X1 NAND3X1_101 ( .A(_239_), .B(_247_), .C(_244_), .Y(_248_) );
OAI21X1 OAI21X1_82 ( .A(i_add2[39]), .B(i_add1[39]), .C(_248_), .Y(_249_) );
INVX1 INVX1_195 ( .A(_249_), .Y(w_C_40_) );
INVX1 INVX1_196 ( .A(i_add2[40]), .Y(_250_) );
INVX1 INVX1_197 ( .A(i_add1[40]), .Y(_251_) );
NOR2X1 NOR2X1_113 ( .A(_250_), .B(_251_), .Y(_252_) );
INVX1 INVX1_198 ( .A(_252_), .Y(_253_) );
NOR2X1 NOR2X1_114 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_254_) );
INVX1 INVX1_199 ( .A(_254_), .Y(_255_) );
NOR2X1 NOR2X1_115 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_256_) );
INVX1 INVX1_200 ( .A(_256_), .Y(_257_) );
NAND3X1 NAND3X1_102 ( .A(_255_), .B(_257_), .C(_248_), .Y(_258_) );
AND2X2 AND2X2_89 ( .A(_258_), .B(_253_), .Y(_259_) );
INVX1 INVX1_201 ( .A(_259_), .Y(w_C_41_) );
AND2X2 AND2X2_90 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_260_) );
INVX1 INVX1_202 ( .A(_260_), .Y(_261_) );
NAND3X1 NAND3X1_103 ( .A(_253_), .B(_261_), .C(_258_), .Y(_262_) );
OAI21X1 OAI21X1_83 ( .A(i_add2[41]), .B(i_add1[41]), .C(_262_), .Y(_263_) );
INVX1 INVX1_203 ( .A(_263_), .Y(w_C_42_) );
INVX1 INVX1_204 ( .A(i_add2[42]), .Y(_264_) );
INVX1 INVX1_205 ( .A(i_add1[42]), .Y(_265_) );
NOR2X1 NOR2X1_116 ( .A(_264_), .B(_265_), .Y(_266_) );
INVX1 INVX1_206 ( .A(_266_), .Y(_267_) );
NOR2X1 NOR2X1_117 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_268_) );
INVX1 INVX1_207 ( .A(_268_), .Y(_269_) );
NOR2X1 NOR2X1_118 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_270_) );
INVX1 INVX1_208 ( .A(_270_), .Y(_271_) );
NAND3X1 NAND3X1_104 ( .A(_269_), .B(_271_), .C(_262_), .Y(_272_) );
AND2X2 AND2X2_91 ( .A(_272_), .B(_267_), .Y(_273_) );
INVX1 INVX1_209 ( .A(_273_), .Y(w_C_43_) );
AND2X2 AND2X2_92 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_274_) );
INVX1 INVX1_210 ( .A(_274_), .Y(_275_) );
NAND3X1 NAND3X1_105 ( .A(_267_), .B(_275_), .C(_272_), .Y(_276_) );
OAI21X1 OAI21X1_84 ( .A(i_add2[43]), .B(i_add1[43]), .C(_276_), .Y(_277_) );
INVX1 INVX1_211 ( .A(_277_), .Y(w_C_44_) );
INVX1 INVX1_212 ( .A(i_add2[44]), .Y(_278_) );
INVX1 INVX1_213 ( .A(i_add1[44]), .Y(_279_) );
NOR2X1 NOR2X1_119 ( .A(_278_), .B(_279_), .Y(_280_) );
INVX1 INVX1_214 ( .A(_280_), .Y(_281_) );
NOR2X1 NOR2X1_120 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_282_) );
INVX1 INVX1_215 ( .A(_282_), .Y(_283_) );
NOR2X1 NOR2X1_121 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_284_) );
INVX1 INVX1_216 ( .A(_284_), .Y(_285_) );
NAND3X1 NAND3X1_106 ( .A(_283_), .B(_285_), .C(_276_), .Y(_286_) );
AND2X2 AND2X2_93 ( .A(_286_), .B(_281_), .Y(_287_) );
INVX1 INVX1_217 ( .A(_287_), .Y(w_C_45_) );
AND2X2 AND2X2_94 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_288_) );
INVX1 INVX1_218 ( .A(_288_), .Y(_289_) );
NAND3X1 NAND3X1_107 ( .A(_281_), .B(_289_), .C(_286_), .Y(_290_) );
OAI21X1 OAI21X1_85 ( .A(i_add2[45]), .B(i_add1[45]), .C(_290_), .Y(_291_) );
INVX1 INVX1_219 ( .A(_291_), .Y(w_C_46_) );
NAND2X1 NAND2X1_131 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_292_) );
NOR2X1 NOR2X1_122 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_293_) );
OAI21X1 OAI21X1_86 ( .A(_293_), .B(_291_), .C(_292_), .Y(w_C_47_) );
OR2X2 OR2X2_64 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_294_) );
NOR2X1 NOR2X1_123 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_295_) );
INVX1 INVX1_220 ( .A(_295_), .Y(_296_) );
INVX1 INVX1_221 ( .A(_293_), .Y(_297_) );
NAND3X1 NAND3X1_108 ( .A(_296_), .B(_297_), .C(_290_), .Y(_298_) );
NAND2X1 NAND2X1_132 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_299_) );
NAND3X1 NAND3X1_109 ( .A(_292_), .B(_299_), .C(_298_), .Y(_300_) );
AND2X2 AND2X2_95 ( .A(_300_), .B(_294_), .Y(w_C_48_) );
INVX1 INVX1_222 ( .A(i_add2[48]), .Y(_301_) );
INVX1 INVX1_223 ( .A(i_add1[48]), .Y(_302_) );
NAND2X1 NAND2X1_133 ( .A(_301_), .B(_302_), .Y(_303_) );
NAND3X1 NAND3X1_110 ( .A(_294_), .B(_303_), .C(_300_), .Y(_304_) );
OAI21X1 OAI21X1_87 ( .A(_301_), .B(_302_), .C(_304_), .Y(w_C_49_) );
INVX1 INVX1_224 ( .A(i_add2[49]), .Y(_305_) );
INVX1 INVX1_225 ( .A(i_add1[49]), .Y(_306_) );
NAND2X1 NAND2X1_134 ( .A(_305_), .B(_306_), .Y(_307_) );
NAND2X1 NAND2X1_135 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_308_) );
NAND2X1 NAND2X1_136 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_309_) );
NAND3X1 NAND3X1_111 ( .A(_308_), .B(_309_), .C(_304_), .Y(_310_) );
AND2X2 AND2X2_96 ( .A(_310_), .B(_307_), .Y(w_C_50_) );
INVX1 INVX1_226 ( .A(i_add2[50]), .Y(_311_) );
INVX1 INVX1_227 ( .A(i_add1[50]), .Y(_312_) );
NAND2X1 NAND2X1_137 ( .A(_311_), .B(_312_), .Y(_313_) );
NAND3X1 NAND3X1_112 ( .A(_307_), .B(_313_), .C(_310_), .Y(_314_) );
OAI21X1 OAI21X1_88 ( .A(_311_), .B(_312_), .C(_314_), .Y(w_C_51_) );
INVX1 INVX1_228 ( .A(i_add2[51]), .Y(_315_) );
INVX1 INVX1_229 ( .A(i_add1[51]), .Y(_316_) );
OAI21X1 OAI21X1_89 ( .A(i_add2[51]), .B(i_add1[51]), .C(w_C_51_), .Y(_317_) );
OAI21X1 OAI21X1_90 ( .A(_315_), .B(_316_), .C(_317_), .Y(w_C_52_) );
NOR2X1 NOR2X1_124 ( .A(_315_), .B(_316_), .Y(_318_) );
INVX1 INVX1_230 ( .A(_318_), .Y(_319_) );
AND2X2 AND2X2_97 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_320_) );
INVX1 INVX1_231 ( .A(_320_), .Y(_321_) );
NAND3X1 NAND3X1_113 ( .A(_319_), .B(_321_), .C(_317_), .Y(_322_) );
OAI21X1 OAI21X1_91 ( .A(i_add2[52]), .B(i_add1[52]), .C(_322_), .Y(_323_) );
INVX1 INVX1_232 ( .A(_323_), .Y(w_C_53_) );
BUFX2 BUFX2_59 ( .A(w_C_57_), .Y(_345__57_) );
BUFX2 BUFX2_60 ( .A(gnd), .Y(w_C_0_) );
endmodule
