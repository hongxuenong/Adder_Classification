module cla_56bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add1[19], i_add1[20], i_add1[21], i_add1[22], i_add1[23], i_add1[24], i_add1[25], i_add1[26], i_add1[27], i_add1[28], i_add1[29], i_add1[30], i_add1[31], i_add1[32], i_add1[33], i_add1[34], i_add1[35], i_add1[36], i_add1[37], i_add1[38], i_add1[39], i_add1[40], i_add1[41], i_add1[42], i_add1[43], i_add1[44], i_add1[45], i_add1[46], i_add1[47], i_add1[48], i_add1[49], i_add1[50], i_add1[51], i_add1[52], i_add1[53], i_add1[54], i_add1[55], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], i_add2[19], i_add2[20], i_add2[21], i_add2[22], i_add2[23], i_add2[24], i_add2[25], i_add2[26], i_add2[27], i_add2[28], i_add2[29], i_add2[30], i_add2[31], i_add2[32], i_add2[33], i_add2[34], i_add2[35], i_add2[36], i_add2[37], i_add2[38], i_add2[39], i_add2[40], i_add2[41], i_add2[42], i_add2[43], i_add2[44], i_add2[45], i_add2[46], i_add2[47], i_add2[48], i_add2[49], i_add2[50], i_add2[51], i_add2[52], i_add2[53], i_add2[54], i_add2[55], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21], o_result[22], o_result[23], o_result[24], o_result[25], o_result[26], o_result[27], o_result[28], o_result[29], o_result[30], o_result[31], o_result[32], o_result[33], o_result[34], o_result[35], o_result[36], o_result[37], o_result[38], o_result[39], o_result[40], o_result[41], o_result[42], o_result[43], o_result[44], o_result[45], o_result[46], o_result[47], o_result[48], o_result[49], o_result[50], o_result[51], o_result[52], o_result[53], o_result[54], o_result[55], o_result[56]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add1[19];
input i_add1[20];
input i_add1[21];
input i_add1[22];
input i_add1[23];
input i_add1[24];
input i_add1[25];
input i_add1[26];
input i_add1[27];
input i_add1[28];
input i_add1[29];
input i_add1[30];
input i_add1[31];
input i_add1[32];
input i_add1[33];
input i_add1[34];
input i_add1[35];
input i_add1[36];
input i_add1[37];
input i_add1[38];
input i_add1[39];
input i_add1[40];
input i_add1[41];
input i_add1[42];
input i_add1[43];
input i_add1[44];
input i_add1[45];
input i_add1[46];
input i_add1[47];
input i_add1[48];
input i_add1[49];
input i_add1[50];
input i_add1[51];
input i_add1[52];
input i_add1[53];
input i_add1[54];
input i_add1[55];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
input i_add2[19];
input i_add2[20];
input i_add2[21];
input i_add2[22];
input i_add2[23];
input i_add2[24];
input i_add2[25];
input i_add2[26];
input i_add2[27];
input i_add2[28];
input i_add2[29];
input i_add2[30];
input i_add2[31];
input i_add2[32];
input i_add2[33];
input i_add2[34];
input i_add2[35];
input i_add2[36];
input i_add2[37];
input i_add2[38];
input i_add2[39];
input i_add2[40];
input i_add2[41];
input i_add2[42];
input i_add2[43];
input i_add2[44];
input i_add2[45];
input i_add2[46];
input i_add2[47];
input i_add2[48];
input i_add2[49];
input i_add2[50];
input i_add2[51];
input i_add2[52];
input i_add2[53];
input i_add2[54];
input i_add2[55];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];
output o_result[22];
output o_result[23];
output o_result[24];
output o_result[25];
output o_result[26];
output o_result[27];
output o_result[28];
output o_result[29];
output o_result[30];
output o_result[31];
output o_result[32];
output o_result[33];
output o_result[34];
output o_result[35];
output o_result[36];
output o_result[37];
output o_result[38];
output o_result[39];
output o_result[40];
output o_result[41];
output o_result[42];
output o_result[43];
output o_result[44];
output o_result[45];
output o_result[46];
output o_result[47];
output o_result[48];
output o_result[49];
output o_result[50];
output o_result[51];
output o_result[52];
output o_result[53];
output o_result[54];
output o_result[55];
output o_result[56];

INVX1 INVX1_1 ( .A(_21_), .Y(w_C_6_) );
AND2X2 AND2X2_1 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_2 ( .A(_22_), .Y(_23_) );
NAND3X1 NAND3X1_1 ( .A(_15_), .B(_23_), .C(_20_), .Y(_24_) );
OAI21X1 OAI21X1_1 ( .A(i_add2[6]), .B(i_add1[6]), .C(_24_), .Y(_25_) );
INVX1 INVX1_3 ( .A(_25_), .Y(w_C_7_) );
INVX1 INVX1_4 ( .A(i_add2[7]), .Y(_26_) );
INVX1 INVX1_5 ( .A(i_add1[7]), .Y(_27_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_28_) );
INVX1 INVX1_6 ( .A(_28_), .Y(_29_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_30_) );
INVX1 INVX1_7 ( .A(_30_), .Y(_31_) );
NAND3X1 NAND3X1_2 ( .A(_29_), .B(_31_), .C(_24_), .Y(_32_) );
OAI21X1 OAI21X1_2 ( .A(_26_), .B(_27_), .C(_32_), .Y(w_C_8_) );
NOR2X1 NOR2X1_3 ( .A(_26_), .B(_27_), .Y(_33_) );
INVX1 INVX1_8 ( .A(_33_), .Y(_34_) );
AND2X2 AND2X2_2 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_35_) );
INVX1 INVX1_9 ( .A(_35_), .Y(_36_) );
NAND3X1 NAND3X1_3 ( .A(_34_), .B(_36_), .C(_32_), .Y(_37_) );
OAI21X1 OAI21X1_3 ( .A(i_add2[8]), .B(i_add1[8]), .C(_37_), .Y(_38_) );
INVX1 INVX1_10 ( .A(_38_), .Y(w_C_9_) );
INVX1 INVX1_11 ( .A(i_add2[9]), .Y(_39_) );
INVX1 INVX1_12 ( .A(i_add1[9]), .Y(_40_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_41_) );
INVX1 INVX1_13 ( .A(_41_), .Y(_42_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_43_) );
INVX1 INVX1_14 ( .A(_43_), .Y(_44_) );
NAND3X1 NAND3X1_4 ( .A(_42_), .B(_44_), .C(_37_), .Y(_45_) );
OAI21X1 OAI21X1_4 ( .A(_39_), .B(_40_), .C(_45_), .Y(w_C_10_) );
NOR2X1 NOR2X1_6 ( .A(_39_), .B(_40_), .Y(_46_) );
INVX1 INVX1_15 ( .A(_46_), .Y(_47_) );
AND2X2 AND2X2_3 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_48_) );
INVX1 INVX1_16 ( .A(_48_), .Y(_49_) );
NAND3X1 NAND3X1_5 ( .A(_47_), .B(_49_), .C(_45_), .Y(_50_) );
OAI21X1 OAI21X1_5 ( .A(i_add2[10]), .B(i_add1[10]), .C(_50_), .Y(_51_) );
INVX1 INVX1_17 ( .A(_51_), .Y(w_C_11_) );
INVX1 INVX1_18 ( .A(i_add2[11]), .Y(_52_) );
INVX1 INVX1_19 ( .A(i_add1[11]), .Y(_53_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_54_) );
INVX1 INVX1_20 ( .A(_54_), .Y(_55_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_56_) );
INVX1 INVX1_21 ( .A(_56_), .Y(_57_) );
NAND3X1 NAND3X1_6 ( .A(_55_), .B(_57_), .C(_50_), .Y(_58_) );
OAI21X1 OAI21X1_6 ( .A(_52_), .B(_53_), .C(_58_), .Y(w_C_12_) );
NOR2X1 NOR2X1_9 ( .A(_52_), .B(_53_), .Y(_59_) );
INVX1 INVX1_22 ( .A(_59_), .Y(_60_) );
AND2X2 AND2X2_4 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_61_) );
INVX1 INVX1_23 ( .A(_61_), .Y(_62_) );
NAND3X1 NAND3X1_7 ( .A(_60_), .B(_62_), .C(_58_), .Y(_63_) );
OAI21X1 OAI21X1_7 ( .A(i_add2[12]), .B(i_add1[12]), .C(_63_), .Y(_64_) );
INVX1 INVX1_24 ( .A(_64_), .Y(w_C_13_) );
INVX1 INVX1_25 ( .A(i_add2[13]), .Y(_65_) );
INVX1 INVX1_26 ( .A(i_add1[13]), .Y(_66_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_67_) );
INVX1 INVX1_27 ( .A(_67_), .Y(_68_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_69_) );
INVX1 INVX1_28 ( .A(_69_), .Y(_70_) );
NAND3X1 NAND3X1_8 ( .A(_68_), .B(_70_), .C(_63_), .Y(_71_) );
OAI21X1 OAI21X1_8 ( .A(_65_), .B(_66_), .C(_71_), .Y(w_C_14_) );
NOR2X1 NOR2X1_12 ( .A(_65_), .B(_66_), .Y(_72_) );
INVX1 INVX1_29 ( .A(_72_), .Y(_73_) );
AND2X2 AND2X2_5 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_74_) );
INVX1 INVX1_30 ( .A(_74_), .Y(_75_) );
NAND3X1 NAND3X1_9 ( .A(_73_), .B(_75_), .C(_71_), .Y(_76_) );
OAI21X1 OAI21X1_9 ( .A(i_add2[14]), .B(i_add1[14]), .C(_76_), .Y(_77_) );
INVX1 INVX1_31 ( .A(_77_), .Y(w_C_15_) );
INVX1 INVX1_32 ( .A(i_add2[15]), .Y(_78_) );
INVX1 INVX1_33 ( .A(i_add1[15]), .Y(_79_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_80_) );
INVX1 INVX1_34 ( .A(_80_), .Y(_81_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_82_) );
INVX1 INVX1_35 ( .A(_82_), .Y(_83_) );
NAND3X1 NAND3X1_10 ( .A(_81_), .B(_83_), .C(_76_), .Y(_84_) );
OAI21X1 OAI21X1_10 ( .A(_78_), .B(_79_), .C(_84_), .Y(w_C_16_) );
NOR2X1 NOR2X1_15 ( .A(_78_), .B(_79_), .Y(_85_) );
INVX1 INVX1_36 ( .A(_85_), .Y(_86_) );
AND2X2 AND2X2_6 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_87_) );
INVX1 INVX1_37 ( .A(_87_), .Y(_88_) );
NAND3X1 NAND3X1_11 ( .A(_86_), .B(_88_), .C(_84_), .Y(_89_) );
OAI21X1 OAI21X1_11 ( .A(i_add2[16]), .B(i_add1[16]), .C(_89_), .Y(_90_) );
INVX1 INVX1_38 ( .A(_90_), .Y(w_C_17_) );
INVX1 INVX1_39 ( .A(i_add2[17]), .Y(_91_) );
INVX1 INVX1_40 ( .A(i_add1[17]), .Y(_92_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_93_) );
INVX1 INVX1_41 ( .A(_93_), .Y(_94_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_95_) );
INVX1 INVX1_42 ( .A(_95_), .Y(_96_) );
NAND3X1 NAND3X1_12 ( .A(_94_), .B(_96_), .C(_89_), .Y(_97_) );
OAI21X1 OAI21X1_12 ( .A(_91_), .B(_92_), .C(_97_), .Y(w_C_18_) );
NOR2X1 NOR2X1_18 ( .A(_91_), .B(_92_), .Y(_98_) );
INVX1 INVX1_43 ( .A(_98_), .Y(_99_) );
AND2X2 AND2X2_7 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_100_) );
INVX1 INVX1_44 ( .A(_100_), .Y(_101_) );
NAND3X1 NAND3X1_13 ( .A(_99_), .B(_101_), .C(_97_), .Y(_102_) );
OAI21X1 OAI21X1_13 ( .A(i_add2[18]), .B(i_add1[18]), .C(_102_), .Y(_103_) );
INVX1 INVX1_45 ( .A(_103_), .Y(w_C_19_) );
INVX1 INVX1_46 ( .A(i_add2[19]), .Y(_104_) );
INVX1 INVX1_47 ( .A(i_add1[19]), .Y(_105_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_106_) );
INVX1 INVX1_48 ( .A(_106_), .Y(_107_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_108_) );
INVX1 INVX1_49 ( .A(_108_), .Y(_109_) );
NAND3X1 NAND3X1_14 ( .A(_107_), .B(_109_), .C(_102_), .Y(_110_) );
OAI21X1 OAI21X1_14 ( .A(_104_), .B(_105_), .C(_110_), .Y(w_C_20_) );
NOR2X1 NOR2X1_21 ( .A(_104_), .B(_105_), .Y(_111_) );
INVX1 INVX1_50 ( .A(_111_), .Y(_112_) );
AND2X2 AND2X2_8 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_113_) );
INVX1 INVX1_51 ( .A(_113_), .Y(_114_) );
NAND3X1 NAND3X1_15 ( .A(_112_), .B(_114_), .C(_110_), .Y(_115_) );
BUFX2 BUFX2_1 ( .A(_330__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_330__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_330__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_330__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_330__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_330__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_330__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_330__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_330__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_330__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_330__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_330__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_330__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_330__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_330__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_330__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_330__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_330__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_330__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_330__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_330__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_330__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_330__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_330__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_330__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_330__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_330__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_330__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_330__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_330__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_330__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_330__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_330__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_330__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_330__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_330__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_330__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(_330__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .A(_330__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .A(_330__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .A(_330__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .A(_330__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .A(_330__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .A(_330__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .A(_330__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .A(_330__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .A(_330__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .A(_330__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .A(_330__48_), .Y(o_result[48]) );
BUFX2 BUFX2_50 ( .A(_330__49_), .Y(o_result[49]) );
BUFX2 BUFX2_51 ( .A(_330__50_), .Y(o_result[50]) );
BUFX2 BUFX2_52 ( .A(_330__51_), .Y(o_result[51]) );
BUFX2 BUFX2_53 ( .A(_330__52_), .Y(o_result[52]) );
BUFX2 BUFX2_54 ( .A(_330__53_), .Y(o_result[53]) );
BUFX2 BUFX2_55 ( .A(_330__54_), .Y(o_result[54]) );
BUFX2 BUFX2_56 ( .A(_330__55_), .Y(o_result[55]) );
BUFX2 BUFX2_57 ( .A(w_C_56_), .Y(o_result[56]) );
INVX1 INVX1_52 ( .A(w_C_4_), .Y(_334_) );
OR2X2 OR2X2_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_335_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_336_) );
NAND3X1 NAND3X1_16 ( .A(_334_), .B(_336_), .C(_335_), .Y(_337_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_331_) );
AND2X2 AND2X2_9 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_332_) );
OAI21X1 OAI21X1_15 ( .A(_331_), .B(_332_), .C(w_C_4_), .Y(_333_) );
NAND2X1 NAND2X1_2 ( .A(_333_), .B(_337_), .Y(_330__4_) );
INVX1 INVX1_53 ( .A(w_C_5_), .Y(_341_) );
OR2X2 OR2X2_2 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_342_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_343_) );
NAND3X1 NAND3X1_17 ( .A(_341_), .B(_343_), .C(_342_), .Y(_344_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_338_) );
AND2X2 AND2X2_10 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_339_) );
OAI21X1 OAI21X1_16 ( .A(_338_), .B(_339_), .C(w_C_5_), .Y(_340_) );
NAND2X1 NAND2X1_4 ( .A(_340_), .B(_344_), .Y(_330__5_) );
INVX1 INVX1_54 ( .A(w_C_6_), .Y(_348_) );
OR2X2 OR2X2_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_349_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_350_) );
NAND3X1 NAND3X1_18 ( .A(_348_), .B(_350_), .C(_349_), .Y(_351_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_345_) );
AND2X2 AND2X2_11 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_346_) );
OAI21X1 OAI21X1_17 ( .A(_345_), .B(_346_), .C(w_C_6_), .Y(_347_) );
NAND2X1 NAND2X1_6 ( .A(_347_), .B(_351_), .Y(_330__6_) );
INVX1 INVX1_55 ( .A(w_C_7_), .Y(_355_) );
OR2X2 OR2X2_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_356_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_357_) );
NAND3X1 NAND3X1_19 ( .A(_355_), .B(_357_), .C(_356_), .Y(_358_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_352_) );
AND2X2 AND2X2_12 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_353_) );
OAI21X1 OAI21X1_18 ( .A(_352_), .B(_353_), .C(w_C_7_), .Y(_354_) );
NAND2X1 NAND2X1_8 ( .A(_354_), .B(_358_), .Y(_330__7_) );
INVX1 INVX1_56 ( .A(w_C_8_), .Y(_362_) );
OR2X2 OR2X2_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_363_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_364_) );
NAND3X1 NAND3X1_20 ( .A(_362_), .B(_364_), .C(_363_), .Y(_365_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_359_) );
AND2X2 AND2X2_13 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_360_) );
OAI21X1 OAI21X1_19 ( .A(_359_), .B(_360_), .C(w_C_8_), .Y(_361_) );
NAND2X1 NAND2X1_10 ( .A(_361_), .B(_365_), .Y(_330__8_) );
INVX1 INVX1_57 ( .A(w_C_9_), .Y(_369_) );
OR2X2 OR2X2_6 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_370_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_371_) );
NAND3X1 NAND3X1_21 ( .A(_369_), .B(_371_), .C(_370_), .Y(_372_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_366_) );
AND2X2 AND2X2_14 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_367_) );
OAI21X1 OAI21X1_20 ( .A(_366_), .B(_367_), .C(w_C_9_), .Y(_368_) );
NAND2X1 NAND2X1_12 ( .A(_368_), .B(_372_), .Y(_330__9_) );
INVX1 INVX1_58 ( .A(w_C_10_), .Y(_376_) );
OR2X2 OR2X2_7 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_377_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_378_) );
NAND3X1 NAND3X1_22 ( .A(_376_), .B(_378_), .C(_377_), .Y(_379_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_373_) );
AND2X2 AND2X2_15 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_374_) );
OAI21X1 OAI21X1_21 ( .A(_373_), .B(_374_), .C(w_C_10_), .Y(_375_) );
NAND2X1 NAND2X1_14 ( .A(_375_), .B(_379_), .Y(_330__10_) );
INVX1 INVX1_59 ( .A(w_C_11_), .Y(_383_) );
OR2X2 OR2X2_8 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_384_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_385_) );
NAND3X1 NAND3X1_23 ( .A(_383_), .B(_385_), .C(_384_), .Y(_386_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_380_) );
AND2X2 AND2X2_16 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_381_) );
OAI21X1 OAI21X1_22 ( .A(_380_), .B(_381_), .C(w_C_11_), .Y(_382_) );
NAND2X1 NAND2X1_16 ( .A(_382_), .B(_386_), .Y(_330__11_) );
INVX1 INVX1_60 ( .A(w_C_12_), .Y(_390_) );
OR2X2 OR2X2_9 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_391_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_392_) );
NAND3X1 NAND3X1_24 ( .A(_390_), .B(_392_), .C(_391_), .Y(_393_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_387_) );
AND2X2 AND2X2_17 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_388_) );
OAI21X1 OAI21X1_23 ( .A(_387_), .B(_388_), .C(w_C_12_), .Y(_389_) );
NAND2X1 NAND2X1_18 ( .A(_389_), .B(_393_), .Y(_330__12_) );
INVX1 INVX1_61 ( .A(w_C_13_), .Y(_397_) );
OR2X2 OR2X2_10 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_398_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_399_) );
NAND3X1 NAND3X1_25 ( .A(_397_), .B(_399_), .C(_398_), .Y(_400_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_394_) );
AND2X2 AND2X2_18 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_395_) );
OAI21X1 OAI21X1_24 ( .A(_394_), .B(_395_), .C(w_C_13_), .Y(_396_) );
NAND2X1 NAND2X1_20 ( .A(_396_), .B(_400_), .Y(_330__13_) );
INVX1 INVX1_62 ( .A(w_C_14_), .Y(_404_) );
OR2X2 OR2X2_11 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_405_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_406_) );
NAND3X1 NAND3X1_26 ( .A(_404_), .B(_406_), .C(_405_), .Y(_407_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_401_) );
AND2X2 AND2X2_19 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_402_) );
OAI21X1 OAI21X1_25 ( .A(_401_), .B(_402_), .C(w_C_14_), .Y(_403_) );
NAND2X1 NAND2X1_22 ( .A(_403_), .B(_407_), .Y(_330__14_) );
INVX1 INVX1_63 ( .A(w_C_15_), .Y(_411_) );
OR2X2 OR2X2_12 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_412_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_413_) );
NAND3X1 NAND3X1_27 ( .A(_411_), .B(_413_), .C(_412_), .Y(_414_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_408_) );
AND2X2 AND2X2_20 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_409_) );
OAI21X1 OAI21X1_26 ( .A(_408_), .B(_409_), .C(w_C_15_), .Y(_410_) );
NAND2X1 NAND2X1_24 ( .A(_410_), .B(_414_), .Y(_330__15_) );
INVX1 INVX1_64 ( .A(w_C_16_), .Y(_418_) );
OR2X2 OR2X2_13 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_419_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_420_) );
NAND3X1 NAND3X1_28 ( .A(_418_), .B(_420_), .C(_419_), .Y(_421_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_415_) );
AND2X2 AND2X2_21 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_416_) );
OAI21X1 OAI21X1_27 ( .A(_415_), .B(_416_), .C(w_C_16_), .Y(_417_) );
NAND2X1 NAND2X1_26 ( .A(_417_), .B(_421_), .Y(_330__16_) );
INVX1 INVX1_65 ( .A(w_C_17_), .Y(_425_) );
OR2X2 OR2X2_14 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_426_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_427_) );
NAND3X1 NAND3X1_29 ( .A(_425_), .B(_427_), .C(_426_), .Y(_428_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_422_) );
AND2X2 AND2X2_22 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_423_) );
OAI21X1 OAI21X1_28 ( .A(_422_), .B(_423_), .C(w_C_17_), .Y(_424_) );
NAND2X1 NAND2X1_28 ( .A(_424_), .B(_428_), .Y(_330__17_) );
INVX1 INVX1_66 ( .A(w_C_18_), .Y(_432_) );
OR2X2 OR2X2_15 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_433_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_434_) );
NAND3X1 NAND3X1_30 ( .A(_432_), .B(_434_), .C(_433_), .Y(_435_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_429_) );
AND2X2 AND2X2_23 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_430_) );
OAI21X1 OAI21X1_29 ( .A(_429_), .B(_430_), .C(w_C_18_), .Y(_431_) );
NAND2X1 NAND2X1_30 ( .A(_431_), .B(_435_), .Y(_330__18_) );
INVX1 INVX1_67 ( .A(w_C_19_), .Y(_439_) );
OR2X2 OR2X2_16 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_440_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_441_) );
NAND3X1 NAND3X1_31 ( .A(_439_), .B(_441_), .C(_440_), .Y(_442_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_436_) );
AND2X2 AND2X2_24 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_437_) );
OAI21X1 OAI21X1_30 ( .A(_436_), .B(_437_), .C(w_C_19_), .Y(_438_) );
NAND2X1 NAND2X1_32 ( .A(_438_), .B(_442_), .Y(_330__19_) );
INVX1 INVX1_68 ( .A(w_C_20_), .Y(_446_) );
OR2X2 OR2X2_17 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_447_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_448_) );
NAND3X1 NAND3X1_32 ( .A(_446_), .B(_448_), .C(_447_), .Y(_449_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_443_) );
AND2X2 AND2X2_25 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_444_) );
OAI21X1 OAI21X1_31 ( .A(_443_), .B(_444_), .C(w_C_20_), .Y(_445_) );
NAND2X1 NAND2X1_34 ( .A(_445_), .B(_449_), .Y(_330__20_) );
INVX1 INVX1_69 ( .A(w_C_21_), .Y(_453_) );
OR2X2 OR2X2_18 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_454_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_455_) );
NAND3X1 NAND3X1_33 ( .A(_453_), .B(_455_), .C(_454_), .Y(_456_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_450_) );
AND2X2 AND2X2_26 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_451_) );
OAI21X1 OAI21X1_32 ( .A(_450_), .B(_451_), .C(w_C_21_), .Y(_452_) );
NAND2X1 NAND2X1_36 ( .A(_452_), .B(_456_), .Y(_330__21_) );
INVX1 INVX1_70 ( .A(w_C_22_), .Y(_460_) );
OR2X2 OR2X2_19 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_461_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_462_) );
NAND3X1 NAND3X1_34 ( .A(_460_), .B(_462_), .C(_461_), .Y(_463_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_457_) );
AND2X2 AND2X2_27 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_458_) );
OAI21X1 OAI21X1_33 ( .A(_457_), .B(_458_), .C(w_C_22_), .Y(_459_) );
NAND2X1 NAND2X1_38 ( .A(_459_), .B(_463_), .Y(_330__22_) );
INVX1 INVX1_71 ( .A(w_C_23_), .Y(_467_) );
OR2X2 OR2X2_20 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_468_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_469_) );
NAND3X1 NAND3X1_35 ( .A(_467_), .B(_469_), .C(_468_), .Y(_470_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_464_) );
AND2X2 AND2X2_28 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_465_) );
OAI21X1 OAI21X1_34 ( .A(_464_), .B(_465_), .C(w_C_23_), .Y(_466_) );
NAND2X1 NAND2X1_40 ( .A(_466_), .B(_470_), .Y(_330__23_) );
INVX1 INVX1_72 ( .A(w_C_24_), .Y(_474_) );
OR2X2 OR2X2_21 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_475_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_476_) );
NAND3X1 NAND3X1_36 ( .A(_474_), .B(_476_), .C(_475_), .Y(_477_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_471_) );
AND2X2 AND2X2_29 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_472_) );
OAI21X1 OAI21X1_35 ( .A(_471_), .B(_472_), .C(w_C_24_), .Y(_473_) );
NAND2X1 NAND2X1_42 ( .A(_473_), .B(_477_), .Y(_330__24_) );
INVX1 INVX1_73 ( .A(w_C_25_), .Y(_481_) );
OR2X2 OR2X2_22 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_482_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_483_) );
NAND3X1 NAND3X1_37 ( .A(_481_), .B(_483_), .C(_482_), .Y(_484_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_478_) );
AND2X2 AND2X2_30 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_479_) );
OAI21X1 OAI21X1_36 ( .A(_478_), .B(_479_), .C(w_C_25_), .Y(_480_) );
NAND2X1 NAND2X1_44 ( .A(_480_), .B(_484_), .Y(_330__25_) );
INVX1 INVX1_74 ( .A(w_C_26_), .Y(_488_) );
OR2X2 OR2X2_23 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_489_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_490_) );
NAND3X1 NAND3X1_38 ( .A(_488_), .B(_490_), .C(_489_), .Y(_491_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_485_) );
AND2X2 AND2X2_31 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_486_) );
OAI21X1 OAI21X1_37 ( .A(_485_), .B(_486_), .C(w_C_26_), .Y(_487_) );
NAND2X1 NAND2X1_46 ( .A(_487_), .B(_491_), .Y(_330__26_) );
INVX1 INVX1_75 ( .A(w_C_27_), .Y(_495_) );
OR2X2 OR2X2_24 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_496_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_497_) );
NAND3X1 NAND3X1_39 ( .A(_495_), .B(_497_), .C(_496_), .Y(_498_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_492_) );
AND2X2 AND2X2_32 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_493_) );
OAI21X1 OAI21X1_38 ( .A(_492_), .B(_493_), .C(w_C_27_), .Y(_494_) );
NAND2X1 NAND2X1_48 ( .A(_494_), .B(_498_), .Y(_330__27_) );
INVX1 INVX1_76 ( .A(w_C_28_), .Y(_502_) );
OR2X2 OR2X2_25 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_503_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_504_) );
NAND3X1 NAND3X1_40 ( .A(_502_), .B(_504_), .C(_503_), .Y(_505_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_499_) );
AND2X2 AND2X2_33 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_500_) );
OAI21X1 OAI21X1_39 ( .A(_499_), .B(_500_), .C(w_C_28_), .Y(_501_) );
NAND2X1 NAND2X1_50 ( .A(_501_), .B(_505_), .Y(_330__28_) );
INVX1 INVX1_77 ( .A(w_C_29_), .Y(_509_) );
OR2X2 OR2X2_26 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_510_) );
NAND2X1 NAND2X1_51 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_511_) );
NAND3X1 NAND3X1_41 ( .A(_509_), .B(_511_), .C(_510_), .Y(_512_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_506_) );
AND2X2 AND2X2_34 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_507_) );
OAI21X1 OAI21X1_40 ( .A(_506_), .B(_507_), .C(w_C_29_), .Y(_508_) );
NAND2X1 NAND2X1_52 ( .A(_508_), .B(_512_), .Y(_330__29_) );
INVX1 INVX1_78 ( .A(w_C_30_), .Y(_516_) );
OR2X2 OR2X2_27 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_517_) );
NAND2X1 NAND2X1_53 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_518_) );
NAND3X1 NAND3X1_42 ( .A(_516_), .B(_518_), .C(_517_), .Y(_519_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_513_) );
AND2X2 AND2X2_35 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_514_) );
OAI21X1 OAI21X1_41 ( .A(_513_), .B(_514_), .C(w_C_30_), .Y(_515_) );
NAND2X1 NAND2X1_54 ( .A(_515_), .B(_519_), .Y(_330__30_) );
INVX1 INVX1_79 ( .A(w_C_31_), .Y(_523_) );
OR2X2 OR2X2_28 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_524_) );
NAND2X1 NAND2X1_55 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_525_) );
NAND3X1 NAND3X1_43 ( .A(_523_), .B(_525_), .C(_524_), .Y(_526_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_520_) );
AND2X2 AND2X2_36 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_521_) );
OAI21X1 OAI21X1_42 ( .A(_520_), .B(_521_), .C(w_C_31_), .Y(_522_) );
NAND2X1 NAND2X1_56 ( .A(_522_), .B(_526_), .Y(_330__31_) );
INVX1 INVX1_80 ( .A(w_C_32_), .Y(_530_) );
OR2X2 OR2X2_29 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_531_) );
NAND2X1 NAND2X1_57 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_532_) );
NAND3X1 NAND3X1_44 ( .A(_530_), .B(_532_), .C(_531_), .Y(_533_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_527_) );
AND2X2 AND2X2_37 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_528_) );
OAI21X1 OAI21X1_43 ( .A(_527_), .B(_528_), .C(w_C_32_), .Y(_529_) );
NAND2X1 NAND2X1_58 ( .A(_529_), .B(_533_), .Y(_330__32_) );
INVX1 INVX1_81 ( .A(w_C_33_), .Y(_537_) );
OR2X2 OR2X2_30 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_538_) );
NAND2X1 NAND2X1_59 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_539_) );
NAND3X1 NAND3X1_45 ( .A(_537_), .B(_539_), .C(_538_), .Y(_540_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_534_) );
AND2X2 AND2X2_38 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_535_) );
OAI21X1 OAI21X1_44 ( .A(_534_), .B(_535_), .C(w_C_33_), .Y(_536_) );
NAND2X1 NAND2X1_60 ( .A(_536_), .B(_540_), .Y(_330__33_) );
INVX1 INVX1_82 ( .A(w_C_34_), .Y(_544_) );
OR2X2 OR2X2_31 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_545_) );
NAND2X1 NAND2X1_61 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_546_) );
NAND3X1 NAND3X1_46 ( .A(_544_), .B(_546_), .C(_545_), .Y(_547_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_541_) );
AND2X2 AND2X2_39 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_542_) );
OAI21X1 OAI21X1_45 ( .A(_541_), .B(_542_), .C(w_C_34_), .Y(_543_) );
NAND2X1 NAND2X1_62 ( .A(_543_), .B(_547_), .Y(_330__34_) );
INVX1 INVX1_83 ( .A(w_C_35_), .Y(_551_) );
OR2X2 OR2X2_32 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_552_) );
NAND2X1 NAND2X1_63 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_553_) );
NAND3X1 NAND3X1_47 ( .A(_551_), .B(_553_), .C(_552_), .Y(_554_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_548_) );
AND2X2 AND2X2_40 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_549_) );
OAI21X1 OAI21X1_46 ( .A(_548_), .B(_549_), .C(w_C_35_), .Y(_550_) );
NAND2X1 NAND2X1_64 ( .A(_550_), .B(_554_), .Y(_330__35_) );
INVX1 INVX1_84 ( .A(w_C_36_), .Y(_558_) );
OR2X2 OR2X2_33 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_559_) );
NAND2X1 NAND2X1_65 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_560_) );
NAND3X1 NAND3X1_48 ( .A(_558_), .B(_560_), .C(_559_), .Y(_561_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_555_) );
AND2X2 AND2X2_41 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_556_) );
OAI21X1 OAI21X1_47 ( .A(_555_), .B(_556_), .C(w_C_36_), .Y(_557_) );
NAND2X1 NAND2X1_66 ( .A(_557_), .B(_561_), .Y(_330__36_) );
INVX1 INVX1_85 ( .A(w_C_37_), .Y(_565_) );
OR2X2 OR2X2_34 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_566_) );
NAND2X1 NAND2X1_67 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_567_) );
NAND3X1 NAND3X1_49 ( .A(_565_), .B(_567_), .C(_566_), .Y(_568_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_562_) );
AND2X2 AND2X2_42 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_563_) );
OAI21X1 OAI21X1_48 ( .A(_562_), .B(_563_), .C(w_C_37_), .Y(_564_) );
NAND2X1 NAND2X1_68 ( .A(_564_), .B(_568_), .Y(_330__37_) );
INVX1 INVX1_86 ( .A(w_C_38_), .Y(_572_) );
OR2X2 OR2X2_35 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_573_) );
NAND2X1 NAND2X1_69 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_574_) );
NAND3X1 NAND3X1_50 ( .A(_572_), .B(_574_), .C(_573_), .Y(_575_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_569_) );
AND2X2 AND2X2_43 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_570_) );
OAI21X1 OAI21X1_49 ( .A(_569_), .B(_570_), .C(w_C_38_), .Y(_571_) );
NAND2X1 NAND2X1_70 ( .A(_571_), .B(_575_), .Y(_330__38_) );
INVX1 INVX1_87 ( .A(w_C_39_), .Y(_579_) );
OR2X2 OR2X2_36 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_580_) );
NAND2X1 NAND2X1_71 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_581_) );
NAND3X1 NAND3X1_51 ( .A(_579_), .B(_581_), .C(_580_), .Y(_582_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_576_) );
AND2X2 AND2X2_44 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_577_) );
OAI21X1 OAI21X1_50 ( .A(_576_), .B(_577_), .C(w_C_39_), .Y(_578_) );
NAND2X1 NAND2X1_72 ( .A(_578_), .B(_582_), .Y(_330__39_) );
INVX1 INVX1_88 ( .A(w_C_40_), .Y(_586_) );
OR2X2 OR2X2_37 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_587_) );
NAND2X1 NAND2X1_73 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_588_) );
NAND3X1 NAND3X1_52 ( .A(_586_), .B(_588_), .C(_587_), .Y(_589_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_583_) );
AND2X2 AND2X2_45 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_584_) );
OAI21X1 OAI21X1_51 ( .A(_583_), .B(_584_), .C(w_C_40_), .Y(_585_) );
NAND2X1 NAND2X1_74 ( .A(_585_), .B(_589_), .Y(_330__40_) );
INVX1 INVX1_89 ( .A(w_C_41_), .Y(_593_) );
OR2X2 OR2X2_38 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_594_) );
NAND2X1 NAND2X1_75 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_595_) );
NAND3X1 NAND3X1_53 ( .A(_593_), .B(_595_), .C(_594_), .Y(_596_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_590_) );
AND2X2 AND2X2_46 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_591_) );
OAI21X1 OAI21X1_52 ( .A(_590_), .B(_591_), .C(w_C_41_), .Y(_592_) );
NAND2X1 NAND2X1_76 ( .A(_592_), .B(_596_), .Y(_330__41_) );
INVX1 INVX1_90 ( .A(w_C_42_), .Y(_600_) );
OR2X2 OR2X2_39 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_601_) );
NAND2X1 NAND2X1_77 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_602_) );
NAND3X1 NAND3X1_54 ( .A(_600_), .B(_602_), .C(_601_), .Y(_603_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_597_) );
AND2X2 AND2X2_47 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_598_) );
OAI21X1 OAI21X1_53 ( .A(_597_), .B(_598_), .C(w_C_42_), .Y(_599_) );
NAND2X1 NAND2X1_78 ( .A(_599_), .B(_603_), .Y(_330__42_) );
INVX1 INVX1_91 ( .A(w_C_43_), .Y(_607_) );
OR2X2 OR2X2_40 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_608_) );
NAND2X1 NAND2X1_79 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_609_) );
NAND3X1 NAND3X1_55 ( .A(_607_), .B(_609_), .C(_608_), .Y(_610_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_604_) );
AND2X2 AND2X2_48 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_605_) );
OAI21X1 OAI21X1_54 ( .A(_604_), .B(_605_), .C(w_C_43_), .Y(_606_) );
NAND2X1 NAND2X1_80 ( .A(_606_), .B(_610_), .Y(_330__43_) );
INVX1 INVX1_92 ( .A(w_C_44_), .Y(_614_) );
OR2X2 OR2X2_41 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_615_) );
NAND2X1 NAND2X1_81 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_616_) );
NAND3X1 NAND3X1_56 ( .A(_614_), .B(_616_), .C(_615_), .Y(_617_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_611_) );
AND2X2 AND2X2_49 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_612_) );
OAI21X1 OAI21X1_55 ( .A(_611_), .B(_612_), .C(w_C_44_), .Y(_613_) );
NAND2X1 NAND2X1_82 ( .A(_613_), .B(_617_), .Y(_330__44_) );
INVX1 INVX1_93 ( .A(w_C_45_), .Y(_621_) );
OR2X2 OR2X2_42 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_622_) );
NAND2X1 NAND2X1_83 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_623_) );
NAND3X1 NAND3X1_57 ( .A(_621_), .B(_623_), .C(_622_), .Y(_624_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_618_) );
AND2X2 AND2X2_50 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_619_) );
OAI21X1 OAI21X1_56 ( .A(_618_), .B(_619_), .C(w_C_45_), .Y(_620_) );
NAND2X1 NAND2X1_84 ( .A(_620_), .B(_624_), .Y(_330__45_) );
INVX1 INVX1_94 ( .A(w_C_46_), .Y(_628_) );
OR2X2 OR2X2_43 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_629_) );
NAND2X1 NAND2X1_85 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_630_) );
NAND3X1 NAND3X1_58 ( .A(_628_), .B(_630_), .C(_629_), .Y(_631_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_625_) );
AND2X2 AND2X2_51 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_626_) );
OAI21X1 OAI21X1_57 ( .A(_625_), .B(_626_), .C(w_C_46_), .Y(_627_) );
NAND2X1 NAND2X1_86 ( .A(_627_), .B(_631_), .Y(_330__46_) );
INVX1 INVX1_95 ( .A(w_C_47_), .Y(_635_) );
OR2X2 OR2X2_44 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_636_) );
NAND2X1 NAND2X1_87 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_637_) );
NAND3X1 NAND3X1_59 ( .A(_635_), .B(_637_), .C(_636_), .Y(_638_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_632_) );
AND2X2 AND2X2_52 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_633_) );
OAI21X1 OAI21X1_58 ( .A(_632_), .B(_633_), .C(w_C_47_), .Y(_634_) );
NAND2X1 NAND2X1_88 ( .A(_634_), .B(_638_), .Y(_330__47_) );
INVX1 INVX1_96 ( .A(w_C_48_), .Y(_642_) );
OR2X2 OR2X2_45 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_643_) );
NAND2X1 NAND2X1_89 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_644_) );
NAND3X1 NAND3X1_60 ( .A(_642_), .B(_644_), .C(_643_), .Y(_645_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_639_) );
AND2X2 AND2X2_53 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_640_) );
OAI21X1 OAI21X1_59 ( .A(_639_), .B(_640_), .C(w_C_48_), .Y(_641_) );
NAND2X1 NAND2X1_90 ( .A(_641_), .B(_645_), .Y(_330__48_) );
INVX1 INVX1_97 ( .A(w_C_49_), .Y(_649_) );
OR2X2 OR2X2_46 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_650_) );
NAND2X1 NAND2X1_91 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_651_) );
NAND3X1 NAND3X1_61 ( .A(_649_), .B(_651_), .C(_650_), .Y(_652_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_646_) );
AND2X2 AND2X2_54 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_647_) );
OAI21X1 OAI21X1_60 ( .A(_646_), .B(_647_), .C(w_C_49_), .Y(_648_) );
NAND2X1 NAND2X1_92 ( .A(_648_), .B(_652_), .Y(_330__49_) );
INVX1 INVX1_98 ( .A(w_C_50_), .Y(_656_) );
OR2X2 OR2X2_47 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_657_) );
NAND2X1 NAND2X1_93 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_658_) );
NAND3X1 NAND3X1_62 ( .A(_656_), .B(_658_), .C(_657_), .Y(_659_) );
NOR2X1 NOR2X1_68 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_653_) );
AND2X2 AND2X2_55 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_654_) );
OAI21X1 OAI21X1_61 ( .A(_653_), .B(_654_), .C(w_C_50_), .Y(_655_) );
NAND2X1 NAND2X1_94 ( .A(_655_), .B(_659_), .Y(_330__50_) );
INVX1 INVX1_99 ( .A(w_C_51_), .Y(_663_) );
OR2X2 OR2X2_48 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_664_) );
NAND2X1 NAND2X1_95 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_665_) );
NAND3X1 NAND3X1_63 ( .A(_663_), .B(_665_), .C(_664_), .Y(_666_) );
NOR2X1 NOR2X1_69 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_660_) );
AND2X2 AND2X2_56 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_661_) );
OAI21X1 OAI21X1_62 ( .A(_660_), .B(_661_), .C(w_C_51_), .Y(_662_) );
NAND2X1 NAND2X1_96 ( .A(_662_), .B(_666_), .Y(_330__51_) );
INVX1 INVX1_100 ( .A(w_C_52_), .Y(_670_) );
OR2X2 OR2X2_49 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_671_) );
NAND2X1 NAND2X1_97 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_672_) );
NAND3X1 NAND3X1_64 ( .A(_670_), .B(_672_), .C(_671_), .Y(_673_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_667_) );
AND2X2 AND2X2_57 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_668_) );
OAI21X1 OAI21X1_63 ( .A(_667_), .B(_668_), .C(w_C_52_), .Y(_669_) );
NAND2X1 NAND2X1_98 ( .A(_669_), .B(_673_), .Y(_330__52_) );
INVX1 INVX1_101 ( .A(w_C_53_), .Y(_677_) );
OR2X2 OR2X2_50 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_678_) );
NAND2X1 NAND2X1_99 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_679_) );
NAND3X1 NAND3X1_65 ( .A(_677_), .B(_679_), .C(_678_), .Y(_680_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_674_) );
AND2X2 AND2X2_58 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_675_) );
OAI21X1 OAI21X1_64 ( .A(_674_), .B(_675_), .C(w_C_53_), .Y(_676_) );
NAND2X1 NAND2X1_100 ( .A(_676_), .B(_680_), .Y(_330__53_) );
INVX1 INVX1_102 ( .A(w_C_54_), .Y(_684_) );
OR2X2 OR2X2_51 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_685_) );
NAND2X1 NAND2X1_101 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_686_) );
NAND3X1 NAND3X1_66 ( .A(_684_), .B(_686_), .C(_685_), .Y(_687_) );
NOR2X1 NOR2X1_72 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_681_) );
AND2X2 AND2X2_59 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_682_) );
OAI21X1 OAI21X1_65 ( .A(_681_), .B(_682_), .C(w_C_54_), .Y(_683_) );
NAND2X1 NAND2X1_102 ( .A(_683_), .B(_687_), .Y(_330__54_) );
INVX1 INVX1_103 ( .A(w_C_55_), .Y(_691_) );
OR2X2 OR2X2_52 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_692_) );
NAND2X1 NAND2X1_103 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_693_) );
NAND3X1 NAND3X1_67 ( .A(_691_), .B(_693_), .C(_692_), .Y(_694_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_688_) );
AND2X2 AND2X2_60 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_689_) );
OAI21X1 OAI21X1_66 ( .A(_688_), .B(_689_), .C(w_C_55_), .Y(_690_) );
NAND2X1 NAND2X1_104 ( .A(_690_), .B(_694_), .Y(_330__55_) );
INVX1 INVX1_104 ( .A(1'b0), .Y(_698_) );
OR2X2 OR2X2_53 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_699_) );
NAND2X1 NAND2X1_105 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_700_) );
NAND3X1 NAND3X1_68 ( .A(_698_), .B(_700_), .C(_699_), .Y(_701_) );
NOR2X1 NOR2X1_74 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_695_) );
AND2X2 AND2X2_61 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_696_) );
OAI21X1 OAI21X1_67 ( .A(_695_), .B(_696_), .C(1'b0), .Y(_697_) );
NAND2X1 NAND2X1_106 ( .A(_697_), .B(_701_), .Y(_330__0_) );
INVX1 INVX1_105 ( .A(w_C_1_), .Y(_705_) );
OR2X2 OR2X2_54 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_706_) );
NAND2X1 NAND2X1_107 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_707_) );
NAND3X1 NAND3X1_69 ( .A(_705_), .B(_707_), .C(_706_), .Y(_708_) );
NOR2X1 NOR2X1_75 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_702_) );
AND2X2 AND2X2_62 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_703_) );
OAI21X1 OAI21X1_68 ( .A(_702_), .B(_703_), .C(w_C_1_), .Y(_704_) );
NAND2X1 NAND2X1_108 ( .A(_704_), .B(_708_), .Y(_330__1_) );
INVX1 INVX1_106 ( .A(w_C_2_), .Y(_712_) );
OR2X2 OR2X2_55 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_713_) );
NAND2X1 NAND2X1_109 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_714_) );
NAND3X1 NAND3X1_70 ( .A(_712_), .B(_714_), .C(_713_), .Y(_715_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_709_) );
AND2X2 AND2X2_63 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_710_) );
OAI21X1 OAI21X1_69 ( .A(_709_), .B(_710_), .C(w_C_2_), .Y(_711_) );
NAND2X1 NAND2X1_110 ( .A(_711_), .B(_715_), .Y(_330__2_) );
INVX1 INVX1_107 ( .A(w_C_3_), .Y(_719_) );
OR2X2 OR2X2_56 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_720_) );
NAND2X1 NAND2X1_111 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_721_) );
NAND3X1 NAND3X1_71 ( .A(_719_), .B(_721_), .C(_720_), .Y(_722_) );
NOR2X1 NOR2X1_77 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_716_) );
AND2X2 AND2X2_64 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_717_) );
OAI21X1 OAI21X1_70 ( .A(_716_), .B(_717_), .C(w_C_3_), .Y(_718_) );
NAND2X1 NAND2X1_112 ( .A(_718_), .B(_722_), .Y(_330__3_) );
OAI21X1 OAI21X1_71 ( .A(i_add2[20]), .B(i_add1[20]), .C(_115_), .Y(_116_) );
INVX1 INVX1_108 ( .A(_116_), .Y(w_C_21_) );
INVX1 INVX1_109 ( .A(i_add2[21]), .Y(_117_) );
INVX1 INVX1_110 ( .A(i_add1[21]), .Y(_118_) );
NOR2X1 NOR2X1_78 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_119_) );
INVX1 INVX1_111 ( .A(_119_), .Y(_120_) );
NOR2X1 NOR2X1_79 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_121_) );
INVX1 INVX1_112 ( .A(_121_), .Y(_122_) );
NAND3X1 NAND3X1_72 ( .A(_120_), .B(_122_), .C(_115_), .Y(_123_) );
OAI21X1 OAI21X1_72 ( .A(_117_), .B(_118_), .C(_123_), .Y(w_C_22_) );
NOR2X1 NOR2X1_80 ( .A(_117_), .B(_118_), .Y(_124_) );
INVX1 INVX1_113 ( .A(_124_), .Y(_125_) );
AND2X2 AND2X2_65 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_126_) );
INVX1 INVX1_114 ( .A(_126_), .Y(_127_) );
NAND3X1 NAND3X1_73 ( .A(_125_), .B(_127_), .C(_123_), .Y(_128_) );
OAI21X1 OAI21X1_73 ( .A(i_add2[22]), .B(i_add1[22]), .C(_128_), .Y(_129_) );
INVX1 INVX1_115 ( .A(_129_), .Y(w_C_23_) );
INVX1 INVX1_116 ( .A(i_add2[23]), .Y(_130_) );
INVX1 INVX1_117 ( .A(i_add1[23]), .Y(_131_) );
NOR2X1 NOR2X1_81 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_132_) );
INVX1 INVX1_118 ( .A(_132_), .Y(_133_) );
NOR2X1 NOR2X1_82 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_134_) );
INVX1 INVX1_119 ( .A(_134_), .Y(_135_) );
NAND3X1 NAND3X1_74 ( .A(_133_), .B(_135_), .C(_128_), .Y(_136_) );
OAI21X1 OAI21X1_74 ( .A(_130_), .B(_131_), .C(_136_), .Y(w_C_24_) );
NOR2X1 NOR2X1_83 ( .A(_130_), .B(_131_), .Y(_137_) );
INVX1 INVX1_120 ( .A(_137_), .Y(_138_) );
AND2X2 AND2X2_66 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_139_) );
INVX1 INVX1_121 ( .A(_139_), .Y(_140_) );
NAND3X1 NAND3X1_75 ( .A(_138_), .B(_140_), .C(_136_), .Y(_141_) );
OAI21X1 OAI21X1_75 ( .A(i_add2[24]), .B(i_add1[24]), .C(_141_), .Y(_142_) );
INVX1 INVX1_122 ( .A(_142_), .Y(w_C_25_) );
INVX1 INVX1_123 ( .A(i_add2[25]), .Y(_143_) );
INVX1 INVX1_124 ( .A(i_add1[25]), .Y(_144_) );
NOR2X1 NOR2X1_84 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_145_) );
INVX1 INVX1_125 ( .A(_145_), .Y(_146_) );
NOR2X1 NOR2X1_85 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_147_) );
INVX1 INVX1_126 ( .A(_147_), .Y(_148_) );
NAND3X1 NAND3X1_76 ( .A(_146_), .B(_148_), .C(_141_), .Y(_149_) );
OAI21X1 OAI21X1_76 ( .A(_143_), .B(_144_), .C(_149_), .Y(w_C_26_) );
NOR2X1 NOR2X1_86 ( .A(_143_), .B(_144_), .Y(_150_) );
INVX1 INVX1_127 ( .A(_150_), .Y(_151_) );
AND2X2 AND2X2_67 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_152_) );
INVX1 INVX1_128 ( .A(_152_), .Y(_153_) );
NAND3X1 NAND3X1_77 ( .A(_151_), .B(_153_), .C(_149_), .Y(_154_) );
OAI21X1 OAI21X1_77 ( .A(i_add2[26]), .B(i_add1[26]), .C(_154_), .Y(_155_) );
INVX1 INVX1_129 ( .A(_155_), .Y(w_C_27_) );
INVX1 INVX1_130 ( .A(i_add2[27]), .Y(_156_) );
INVX1 INVX1_131 ( .A(i_add1[27]), .Y(_157_) );
NOR2X1 NOR2X1_87 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_158_) );
INVX1 INVX1_132 ( .A(_158_), .Y(_159_) );
NOR2X1 NOR2X1_88 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_160_) );
INVX1 INVX1_133 ( .A(_160_), .Y(_161_) );
NAND3X1 NAND3X1_78 ( .A(_159_), .B(_161_), .C(_154_), .Y(_162_) );
OAI21X1 OAI21X1_78 ( .A(_156_), .B(_157_), .C(_162_), .Y(w_C_28_) );
NOR2X1 NOR2X1_89 ( .A(_156_), .B(_157_), .Y(_163_) );
INVX1 INVX1_134 ( .A(_163_), .Y(_164_) );
AND2X2 AND2X2_68 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_165_) );
INVX1 INVX1_135 ( .A(_165_), .Y(_166_) );
NAND3X1 NAND3X1_79 ( .A(_164_), .B(_166_), .C(_162_), .Y(_167_) );
OAI21X1 OAI21X1_79 ( .A(i_add2[28]), .B(i_add1[28]), .C(_167_), .Y(_168_) );
INVX1 INVX1_136 ( .A(_168_), .Y(w_C_29_) );
INVX1 INVX1_137 ( .A(i_add2[29]), .Y(_169_) );
INVX1 INVX1_138 ( .A(i_add1[29]), .Y(_170_) );
NOR2X1 NOR2X1_90 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_171_) );
INVX1 INVX1_139 ( .A(_171_), .Y(_172_) );
NOR2X1 NOR2X1_91 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_173_) );
INVX1 INVX1_140 ( .A(_173_), .Y(_174_) );
NAND3X1 NAND3X1_80 ( .A(_172_), .B(_174_), .C(_167_), .Y(_175_) );
OAI21X1 OAI21X1_80 ( .A(_169_), .B(_170_), .C(_175_), .Y(w_C_30_) );
NOR2X1 NOR2X1_92 ( .A(_169_), .B(_170_), .Y(_176_) );
INVX1 INVX1_141 ( .A(_176_), .Y(_177_) );
AND2X2 AND2X2_69 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_178_) );
INVX1 INVX1_142 ( .A(_178_), .Y(_179_) );
NAND3X1 NAND3X1_81 ( .A(_177_), .B(_179_), .C(_175_), .Y(_180_) );
OAI21X1 OAI21X1_81 ( .A(i_add2[30]), .B(i_add1[30]), .C(_180_), .Y(_181_) );
INVX1 INVX1_143 ( .A(_181_), .Y(w_C_31_) );
INVX1 INVX1_144 ( .A(i_add2[31]), .Y(_182_) );
INVX1 INVX1_145 ( .A(i_add1[31]), .Y(_183_) );
NOR2X1 NOR2X1_93 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_184_) );
INVX1 INVX1_146 ( .A(_184_), .Y(_185_) );
NOR2X1 NOR2X1_94 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_186_) );
INVX1 INVX1_147 ( .A(_186_), .Y(_187_) );
NAND3X1 NAND3X1_82 ( .A(_185_), .B(_187_), .C(_180_), .Y(_188_) );
OAI21X1 OAI21X1_82 ( .A(_182_), .B(_183_), .C(_188_), .Y(w_C_32_) );
NOR2X1 NOR2X1_95 ( .A(_182_), .B(_183_), .Y(_189_) );
INVX1 INVX1_148 ( .A(_189_), .Y(_190_) );
AND2X2 AND2X2_70 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_191_) );
INVX1 INVX1_149 ( .A(_191_), .Y(_192_) );
NAND3X1 NAND3X1_83 ( .A(_190_), .B(_192_), .C(_188_), .Y(_193_) );
OAI21X1 OAI21X1_83 ( .A(i_add2[32]), .B(i_add1[32]), .C(_193_), .Y(_194_) );
INVX1 INVX1_150 ( .A(_194_), .Y(w_C_33_) );
INVX1 INVX1_151 ( .A(i_add2[33]), .Y(_195_) );
INVX1 INVX1_152 ( .A(i_add1[33]), .Y(_196_) );
NOR2X1 NOR2X1_96 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_197_) );
INVX1 INVX1_153 ( .A(_197_), .Y(_198_) );
NOR2X1 NOR2X1_97 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_199_) );
INVX1 INVX1_154 ( .A(_199_), .Y(_200_) );
NAND3X1 NAND3X1_84 ( .A(_198_), .B(_200_), .C(_193_), .Y(_201_) );
OAI21X1 OAI21X1_84 ( .A(_195_), .B(_196_), .C(_201_), .Y(w_C_34_) );
NOR2X1 NOR2X1_98 ( .A(_195_), .B(_196_), .Y(_202_) );
INVX1 INVX1_155 ( .A(_202_), .Y(_203_) );
AND2X2 AND2X2_71 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_204_) );
INVX1 INVX1_156 ( .A(_204_), .Y(_205_) );
NAND3X1 NAND3X1_85 ( .A(_203_), .B(_205_), .C(_201_), .Y(_206_) );
OAI21X1 OAI21X1_85 ( .A(i_add2[34]), .B(i_add1[34]), .C(_206_), .Y(_207_) );
INVX1 INVX1_157 ( .A(_207_), .Y(w_C_35_) );
INVX1 INVX1_158 ( .A(i_add2[35]), .Y(_208_) );
INVX1 INVX1_159 ( .A(i_add1[35]), .Y(_209_) );
NOR2X1 NOR2X1_99 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_210_) );
INVX1 INVX1_160 ( .A(_210_), .Y(_211_) );
NOR2X1 NOR2X1_100 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_212_) );
INVX1 INVX1_161 ( .A(_212_), .Y(_213_) );
NAND3X1 NAND3X1_86 ( .A(_211_), .B(_213_), .C(_206_), .Y(_214_) );
OAI21X1 OAI21X1_86 ( .A(_208_), .B(_209_), .C(_214_), .Y(w_C_36_) );
NOR2X1 NOR2X1_101 ( .A(_208_), .B(_209_), .Y(_215_) );
INVX1 INVX1_162 ( .A(_215_), .Y(_216_) );
AND2X2 AND2X2_72 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_217_) );
INVX1 INVX1_163 ( .A(_217_), .Y(_218_) );
NAND3X1 NAND3X1_87 ( .A(_216_), .B(_218_), .C(_214_), .Y(_219_) );
OAI21X1 OAI21X1_87 ( .A(i_add2[36]), .B(i_add1[36]), .C(_219_), .Y(_220_) );
INVX1 INVX1_164 ( .A(_220_), .Y(w_C_37_) );
INVX1 INVX1_165 ( .A(i_add2[37]), .Y(_221_) );
INVX1 INVX1_166 ( .A(i_add1[37]), .Y(_222_) );
NOR2X1 NOR2X1_102 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_223_) );
INVX1 INVX1_167 ( .A(_223_), .Y(_224_) );
NOR2X1 NOR2X1_103 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_225_) );
INVX1 INVX1_168 ( .A(_225_), .Y(_226_) );
NAND3X1 NAND3X1_88 ( .A(_224_), .B(_226_), .C(_219_), .Y(_227_) );
OAI21X1 OAI21X1_88 ( .A(_221_), .B(_222_), .C(_227_), .Y(w_C_38_) );
NOR2X1 NOR2X1_104 ( .A(_221_), .B(_222_), .Y(_228_) );
INVX1 INVX1_169 ( .A(_228_), .Y(_229_) );
AND2X2 AND2X2_73 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_230_) );
INVX1 INVX1_170 ( .A(_230_), .Y(_231_) );
NAND3X1 NAND3X1_89 ( .A(_229_), .B(_231_), .C(_227_), .Y(_232_) );
OAI21X1 OAI21X1_89 ( .A(i_add2[38]), .B(i_add1[38]), .C(_232_), .Y(_233_) );
INVX1 INVX1_171 ( .A(_233_), .Y(w_C_39_) );
INVX1 INVX1_172 ( .A(i_add2[39]), .Y(_234_) );
INVX1 INVX1_173 ( .A(i_add1[39]), .Y(_235_) );
NOR2X1 NOR2X1_105 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_236_) );
INVX1 INVX1_174 ( .A(_236_), .Y(_237_) );
NOR2X1 NOR2X1_106 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_238_) );
INVX1 INVX1_175 ( .A(_238_), .Y(_239_) );
NAND3X1 NAND3X1_90 ( .A(_237_), .B(_239_), .C(_232_), .Y(_240_) );
OAI21X1 OAI21X1_90 ( .A(_234_), .B(_235_), .C(_240_), .Y(w_C_40_) );
NOR2X1 NOR2X1_107 ( .A(_234_), .B(_235_), .Y(_241_) );
INVX1 INVX1_176 ( .A(_241_), .Y(_242_) );
AND2X2 AND2X2_74 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_243_) );
INVX1 INVX1_177 ( .A(_243_), .Y(_244_) );
NAND3X1 NAND3X1_91 ( .A(_242_), .B(_244_), .C(_240_), .Y(_245_) );
OAI21X1 OAI21X1_91 ( .A(i_add2[40]), .B(i_add1[40]), .C(_245_), .Y(_246_) );
INVX1 INVX1_178 ( .A(_246_), .Y(w_C_41_) );
INVX1 INVX1_179 ( .A(i_add2[41]), .Y(_247_) );
INVX1 INVX1_180 ( .A(i_add1[41]), .Y(_248_) );
NOR2X1 NOR2X1_108 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_249_) );
INVX1 INVX1_181 ( .A(_249_), .Y(_250_) );
NOR2X1 NOR2X1_109 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_251_) );
INVX1 INVX1_182 ( .A(_251_), .Y(_252_) );
NAND3X1 NAND3X1_92 ( .A(_250_), .B(_252_), .C(_245_), .Y(_253_) );
OAI21X1 OAI21X1_92 ( .A(_247_), .B(_248_), .C(_253_), .Y(w_C_42_) );
NOR2X1 NOR2X1_110 ( .A(_247_), .B(_248_), .Y(_254_) );
INVX1 INVX1_183 ( .A(_254_), .Y(_255_) );
AND2X2 AND2X2_75 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_256_) );
INVX1 INVX1_184 ( .A(_256_), .Y(_257_) );
NAND3X1 NAND3X1_93 ( .A(_255_), .B(_257_), .C(_253_), .Y(_258_) );
OAI21X1 OAI21X1_93 ( .A(i_add2[42]), .B(i_add1[42]), .C(_258_), .Y(_259_) );
INVX1 INVX1_185 ( .A(_259_), .Y(w_C_43_) );
INVX1 INVX1_186 ( .A(i_add2[43]), .Y(_260_) );
INVX1 INVX1_187 ( .A(i_add1[43]), .Y(_261_) );
NOR2X1 NOR2X1_111 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_262_) );
INVX1 INVX1_188 ( .A(_262_), .Y(_263_) );
NOR2X1 NOR2X1_112 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_264_) );
INVX1 INVX1_189 ( .A(_264_), .Y(_265_) );
NAND3X1 NAND3X1_94 ( .A(_263_), .B(_265_), .C(_258_), .Y(_266_) );
OAI21X1 OAI21X1_94 ( .A(_260_), .B(_261_), .C(_266_), .Y(w_C_44_) );
NOR2X1 NOR2X1_113 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_267_) );
INVX1 INVX1_190 ( .A(_267_), .Y(_268_) );
NOR2X1 NOR2X1_114 ( .A(_260_), .B(_261_), .Y(_269_) );
INVX1 INVX1_191 ( .A(_269_), .Y(_270_) );
NAND2X1 NAND2X1_113 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_271_) );
NAND3X1 NAND3X1_95 ( .A(_270_), .B(_271_), .C(_266_), .Y(_272_) );
AND2X2 AND2X2_76 ( .A(_272_), .B(_268_), .Y(w_C_45_) );
INVX1 INVX1_192 ( .A(i_add2[45]), .Y(_273_) );
INVX1 INVX1_193 ( .A(i_add1[45]), .Y(_274_) );
NAND2X1 NAND2X1_114 ( .A(_273_), .B(_274_), .Y(_275_) );
NAND3X1 NAND3X1_96 ( .A(_268_), .B(_275_), .C(_272_), .Y(_276_) );
OAI21X1 OAI21X1_95 ( .A(_273_), .B(_274_), .C(_276_), .Y(w_C_46_) );
INVX1 INVX1_194 ( .A(i_add2[46]), .Y(_277_) );
INVX1 INVX1_195 ( .A(i_add1[46]), .Y(_278_) );
OAI21X1 OAI21X1_96 ( .A(i_add2[46]), .B(i_add1[46]), .C(w_C_46_), .Y(_279_) );
OAI21X1 OAI21X1_97 ( .A(_277_), .B(_278_), .C(_279_), .Y(w_C_47_) );
INVX1 INVX1_196 ( .A(i_add2[47]), .Y(_280_) );
INVX1 INVX1_197 ( .A(i_add1[47]), .Y(_281_) );
NOR2X1 NOR2X1_115 ( .A(_280_), .B(_281_), .Y(_282_) );
OR2X2 OR2X2_57 ( .A(w_C_47_), .B(_282_), .Y(_283_) );
OAI21X1 OAI21X1_98 ( .A(i_add2[47]), .B(i_add1[47]), .C(_283_), .Y(_284_) );
INVX1 INVX1_198 ( .A(_284_), .Y(w_C_48_) );
NAND2X1 NAND2X1_115 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_285_) );
NOR2X1 NOR2X1_116 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_286_) );
OAI21X1 OAI21X1_99 ( .A(_286_), .B(_284_), .C(_285_), .Y(w_C_49_) );
INVX1 INVX1_199 ( .A(i_add2[49]), .Y(_287_) );
INVX1 INVX1_200 ( .A(i_add1[49]), .Y(_288_) );
INVX1 INVX1_201 ( .A(_286_), .Y(_289_) );
INVX1 INVX1_202 ( .A(_282_), .Y(_290_) );
NAND2X1 NAND2X1_116 ( .A(_277_), .B(_278_), .Y(_291_) );
NAND2X1 NAND2X1_117 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_292_) );
NAND2X1 NAND2X1_118 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_293_) );
NAND3X1 NAND3X1_97 ( .A(_292_), .B(_293_), .C(_276_), .Y(_294_) );
NAND2X1 NAND2X1_119 ( .A(_280_), .B(_281_), .Y(_295_) );
NAND3X1 NAND3X1_98 ( .A(_291_), .B(_295_), .C(_294_), .Y(_296_) );
NAND3X1 NAND3X1_99 ( .A(_290_), .B(_285_), .C(_296_), .Y(_297_) );
NAND2X1 NAND2X1_120 ( .A(_287_), .B(_288_), .Y(_298_) );
NAND3X1 NAND3X1_100 ( .A(_289_), .B(_298_), .C(_297_), .Y(_299_) );
OAI21X1 OAI21X1_100 ( .A(_287_), .B(_288_), .C(_299_), .Y(w_C_50_) );
INVX1 INVX1_203 ( .A(i_add2[50]), .Y(_300_) );
INVX1 INVX1_204 ( .A(i_add1[50]), .Y(_301_) );
OAI21X1 OAI21X1_101 ( .A(i_add2[50]), .B(i_add1[50]), .C(w_C_50_), .Y(_302_) );
OAI21X1 OAI21X1_102 ( .A(_300_), .B(_301_), .C(_302_), .Y(w_C_51_) );
NOR2X1 NOR2X1_117 ( .A(_300_), .B(_301_), .Y(_303_) );
INVX1 INVX1_205 ( .A(_303_), .Y(_304_) );
AND2X2 AND2X2_77 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_305_) );
INVX1 INVX1_206 ( .A(_305_), .Y(_306_) );
NAND3X1 NAND3X1_101 ( .A(_304_), .B(_306_), .C(_302_), .Y(_307_) );
OAI21X1 OAI21X1_103 ( .A(i_add2[51]), .B(i_add1[51]), .C(_307_), .Y(_308_) );
INVX1 INVX1_207 ( .A(_308_), .Y(w_C_52_) );
NAND2X1 NAND2X1_121 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_309_) );
NOR2X1 NOR2X1_118 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_310_) );
OAI21X1 OAI21X1_104 ( .A(_310_), .B(_308_), .C(_309_), .Y(w_C_53_) );
NAND2X1 NAND2X1_122 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_311_) );
INVX1 INVX1_208 ( .A(_310_), .Y(_312_) );
NOR2X1 NOR2X1_119 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_313_) );
INVX1 INVX1_209 ( .A(_313_), .Y(_314_) );
NOR2X1 NOR2X1_120 ( .A(_287_), .B(_288_), .Y(_315_) );
INVX1 INVX1_210 ( .A(_315_), .Y(_316_) );
NAND3X1 NAND3X1_102 ( .A(_316_), .B(_304_), .C(_299_), .Y(_317_) );
NOR2X1 NOR2X1_121 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_318_) );
INVX1 INVX1_211 ( .A(_318_), .Y(_319_) );
NAND3X1 NAND3X1_103 ( .A(_314_), .B(_319_), .C(_317_), .Y(_320_) );
NAND3X1 NAND3X1_104 ( .A(_306_), .B(_309_), .C(_320_), .Y(_321_) );
OR2X2 OR2X2_58 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_322_) );
NAND3X1 NAND3X1_105 ( .A(_312_), .B(_322_), .C(_321_), .Y(_323_) );
NAND2X1 NAND2X1_123 ( .A(_311_), .B(_323_), .Y(w_C_54_) );
OR2X2 OR2X2_59 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_324_) );
NAND2X1 NAND2X1_124 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_325_) );
NAND3X1 NAND3X1_106 ( .A(_311_), .B(_325_), .C(_323_), .Y(_326_) );
AND2X2 AND2X2_78 ( .A(_326_), .B(_324_), .Y(w_C_55_) );
NAND2X1 NAND2X1_125 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_327_) );
OR2X2 OR2X2_60 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_328_) );
NAND3X1 NAND3X1_107 ( .A(_324_), .B(_328_), .C(_326_), .Y(_329_) );
NAND2X1 NAND2X1_126 ( .A(_327_), .B(_329_), .Y(w_C_56_) );
NAND2X1 NAND2X1_127 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_212 ( .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_122 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_123 ( .A(_1_), .B(_2_), .Y(w_C_2_) );
INVX1 INVX1_213 ( .A(i_add2[2]), .Y(_3_) );
INVX1 INVX1_214 ( .A(i_add1[2]), .Y(_4_) );
NAND2X1 NAND2X1_128 ( .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_129 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
OAI21X1 OAI21X1_105 ( .A(_1_), .B(_2_), .C(_6_), .Y(_7_) );
AND2X2 AND2X2_79 ( .A(_7_), .B(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_130 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
OR2X2 OR2X2_61 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_108 ( .A(_5_), .B(_9_), .C(_7_), .Y(_10_) );
AND2X2 AND2X2_80 ( .A(_10_), .B(_8_), .Y(_11_) );
INVX1 INVX1_215 ( .A(_11_), .Y(w_C_4_) );
NAND2X1 NAND2X1_131 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_12_) );
NOR2X1 NOR2X1_124 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
OAI21X1 OAI21X1_106 ( .A(_13_), .B(_11_), .C(_12_), .Y(w_C_5_) );
AND2X2 AND2X2_81 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_14_) );
INVX1 INVX1_216 ( .A(_14_), .Y(_15_) );
INVX1 INVX1_217 ( .A(_13_), .Y(_16_) );
NAND3X1 NAND3X1_109 ( .A(_8_), .B(_12_), .C(_10_), .Y(_17_) );
NOR2X1 NOR2X1_125 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_18_) );
INVX1 INVX1_218 ( .A(_18_), .Y(_19_) );
NAND3X1 NAND3X1_110 ( .A(_16_), .B(_19_), .C(_17_), .Y(_20_) );
AND2X2 AND2X2_82 ( .A(_20_), .B(_15_), .Y(_21_) );
BUFX2 BUFX2_58 ( .A(w_C_56_), .Y(_330__56_) );
BUFX2 BUFX2_59 ( .A(1'b0), .Y(w_C_0_) );
endmodule
