module cla_46bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add1[19], i_add1[20], i_add1[21], i_add1[22], i_add1[23], i_add1[24], i_add1[25], i_add1[26], i_add1[27], i_add1[28], i_add1[29], i_add1[30], i_add1[31], i_add1[32], i_add1[33], i_add1[34], i_add1[35], i_add1[36], i_add1[37], i_add1[38], i_add1[39], i_add1[40], i_add1[41], i_add1[42], i_add1[43], i_add1[44], i_add1[45], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], i_add2[19], i_add2[20], i_add2[21], i_add2[22], i_add2[23], i_add2[24], i_add2[25], i_add2[26], i_add2[27], i_add2[28], i_add2[29], i_add2[30], i_add2[31], i_add2[32], i_add2[33], i_add2[34], i_add2[35], i_add2[36], i_add2[37], i_add2[38], i_add2[39], i_add2[40], i_add2[41], i_add2[42], i_add2[43], i_add2[44], i_add2[45], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21], o_result[22], o_result[23], o_result[24], o_result[25], o_result[26], o_result[27], o_result[28], o_result[29], o_result[30], o_result[31], o_result[32], o_result[33], o_result[34], o_result[35], o_result[36], o_result[37], o_result[38], o_result[39], o_result[40], o_result[41], o_result[42], o_result[43], o_result[44], o_result[45], o_result[46]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add1[19];
input i_add1[20];
input i_add1[21];
input i_add1[22];
input i_add1[23];
input i_add1[24];
input i_add1[25];
input i_add1[26];
input i_add1[27];
input i_add1[28];
input i_add1[29];
input i_add1[30];
input i_add1[31];
input i_add1[32];
input i_add1[33];
input i_add1[34];
input i_add1[35];
input i_add1[36];
input i_add1[37];
input i_add1[38];
input i_add1[39];
input i_add1[40];
input i_add1[41];
input i_add1[42];
input i_add1[43];
input i_add1[44];
input i_add1[45];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
input i_add2[19];
input i_add2[20];
input i_add2[21];
input i_add2[22];
input i_add2[23];
input i_add2[24];
input i_add2[25];
input i_add2[26];
input i_add2[27];
input i_add2[28];
input i_add2[29];
input i_add2[30];
input i_add2[31];
input i_add2[32];
input i_add2[33];
input i_add2[34];
input i_add2[35];
input i_add2[36];
input i_add2[37];
input i_add2[38];
input i_add2[39];
input i_add2[40];
input i_add2[41];
input i_add2[42];
input i_add2[43];
input i_add2[44];
input i_add2[45];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];
output o_result[22];
output o_result[23];
output o_result[24];
output o_result[25];
output o_result[26];
output o_result[27];
output o_result[28];
output o_result[29];
output o_result[30];
output o_result[31];
output o_result[32];
output o_result[33];
output o_result[34];
output o_result[35];
output o_result[36];
output o_result[37];
output o_result[38];
output o_result[39];
output o_result[40];
output o_result[41];
output o_result[42];
output o_result[43];
output o_result[44];
output o_result[45];
output o_result[46];

INVX1 INVX1_1 ( .A(w_C_11_), .Y(_317_) );
OR2X2 OR2X2_1 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_318_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_319_) );
NAND3X1 NAND3X1_1 ( .A(_317_), .B(_319_), .C(_318_), .Y(_320_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_314_) );
AND2X2 AND2X2_1 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_315_) );
OAI21X1 OAI21X1_1 ( .A(_314_), .B(_315_), .C(w_C_11_), .Y(_316_) );
NAND2X1 NAND2X1_2 ( .A(_316_), .B(_320_), .Y(_264__11_) );
INVX1 INVX1_2 ( .A(w_C_12_), .Y(_324_) );
OR2X2 OR2X2_2 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_325_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_326_) );
NAND3X1 NAND3X1_2 ( .A(_324_), .B(_326_), .C(_325_), .Y(_327_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_321_) );
AND2X2 AND2X2_2 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_322_) );
OAI21X1 OAI21X1_2 ( .A(_321_), .B(_322_), .C(w_C_12_), .Y(_323_) );
NAND2X1 NAND2X1_4 ( .A(_323_), .B(_327_), .Y(_264__12_) );
INVX1 INVX1_3 ( .A(w_C_13_), .Y(_331_) );
OR2X2 OR2X2_3 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_332_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_333_) );
NAND3X1 NAND3X1_3 ( .A(_331_), .B(_333_), .C(_332_), .Y(_334_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_328_) );
AND2X2 AND2X2_3 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_329_) );
OAI21X1 OAI21X1_3 ( .A(_328_), .B(_329_), .C(w_C_13_), .Y(_330_) );
NAND2X1 NAND2X1_6 ( .A(_330_), .B(_334_), .Y(_264__13_) );
INVX1 INVX1_4 ( .A(w_C_14_), .Y(_338_) );
OR2X2 OR2X2_4 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_339_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_340_) );
NAND3X1 NAND3X1_4 ( .A(_338_), .B(_340_), .C(_339_), .Y(_341_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_335_) );
AND2X2 AND2X2_4 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_336_) );
OAI21X1 OAI21X1_4 ( .A(_335_), .B(_336_), .C(w_C_14_), .Y(_337_) );
NAND2X1 NAND2X1_8 ( .A(_337_), .B(_341_), .Y(_264__14_) );
INVX1 INVX1_5 ( .A(w_C_15_), .Y(_345_) );
OR2X2 OR2X2_5 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_346_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_347_) );
NAND3X1 NAND3X1_5 ( .A(_345_), .B(_347_), .C(_346_), .Y(_348_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_342_) );
AND2X2 AND2X2_5 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_343_) );
OAI21X1 OAI21X1_5 ( .A(_342_), .B(_343_), .C(w_C_15_), .Y(_344_) );
NAND2X1 NAND2X1_10 ( .A(_344_), .B(_348_), .Y(_264__15_) );
INVX1 INVX1_6 ( .A(w_C_16_), .Y(_352_) );
OR2X2 OR2X2_6 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_353_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_354_) );
NAND3X1 NAND3X1_6 ( .A(_352_), .B(_354_), .C(_353_), .Y(_355_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_349_) );
AND2X2 AND2X2_6 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_350_) );
OAI21X1 OAI21X1_6 ( .A(_349_), .B(_350_), .C(w_C_16_), .Y(_351_) );
NAND2X1 NAND2X1_12 ( .A(_351_), .B(_355_), .Y(_264__16_) );
INVX1 INVX1_7 ( .A(w_C_17_), .Y(_359_) );
OR2X2 OR2X2_7 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_360_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_361_) );
NAND3X1 NAND3X1_7 ( .A(_359_), .B(_361_), .C(_360_), .Y(_362_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_356_) );
AND2X2 AND2X2_7 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_357_) );
OAI21X1 OAI21X1_7 ( .A(_356_), .B(_357_), .C(w_C_17_), .Y(_358_) );
NAND2X1 NAND2X1_14 ( .A(_358_), .B(_362_), .Y(_264__17_) );
INVX1 INVX1_8 ( .A(w_C_18_), .Y(_366_) );
OR2X2 OR2X2_8 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_367_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_368_) );
NAND3X1 NAND3X1_8 ( .A(_366_), .B(_368_), .C(_367_), .Y(_369_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_363_) );
AND2X2 AND2X2_8 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_364_) );
OAI21X1 OAI21X1_8 ( .A(_363_), .B(_364_), .C(w_C_18_), .Y(_365_) );
NAND2X1 NAND2X1_16 ( .A(_365_), .B(_369_), .Y(_264__18_) );
INVX1 INVX1_9 ( .A(w_C_19_), .Y(_373_) );
OR2X2 OR2X2_9 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_374_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_375_) );
NAND3X1 NAND3X1_9 ( .A(_373_), .B(_375_), .C(_374_), .Y(_376_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_370_) );
AND2X2 AND2X2_9 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_371_) );
OAI21X1 OAI21X1_9 ( .A(_370_), .B(_371_), .C(w_C_19_), .Y(_372_) );
NAND2X1 NAND2X1_18 ( .A(_372_), .B(_376_), .Y(_264__19_) );
INVX1 INVX1_10 ( .A(w_C_20_), .Y(_380_) );
OR2X2 OR2X2_10 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_381_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_382_) );
NAND3X1 NAND3X1_10 ( .A(_380_), .B(_382_), .C(_381_), .Y(_383_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_377_) );
AND2X2 AND2X2_10 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_378_) );
OAI21X1 OAI21X1_10 ( .A(_377_), .B(_378_), .C(w_C_20_), .Y(_379_) );
NAND2X1 NAND2X1_20 ( .A(_379_), .B(_383_), .Y(_264__20_) );
INVX1 INVX1_11 ( .A(w_C_21_), .Y(_387_) );
OR2X2 OR2X2_11 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_388_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_389_) );
NAND3X1 NAND3X1_11 ( .A(_387_), .B(_389_), .C(_388_), .Y(_390_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_384_) );
AND2X2 AND2X2_11 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_385_) );
OAI21X1 OAI21X1_11 ( .A(_384_), .B(_385_), .C(w_C_21_), .Y(_386_) );
NAND2X1 NAND2X1_22 ( .A(_386_), .B(_390_), .Y(_264__21_) );
INVX1 INVX1_12 ( .A(w_C_22_), .Y(_394_) );
OR2X2 OR2X2_12 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_395_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_396_) );
NAND3X1 NAND3X1_12 ( .A(_394_), .B(_396_), .C(_395_), .Y(_397_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_391_) );
AND2X2 AND2X2_12 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_392_) );
OAI21X1 OAI21X1_12 ( .A(_391_), .B(_392_), .C(w_C_22_), .Y(_393_) );
NAND2X1 NAND2X1_24 ( .A(_393_), .B(_397_), .Y(_264__22_) );
INVX1 INVX1_13 ( .A(w_C_23_), .Y(_401_) );
OR2X2 OR2X2_13 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_402_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_403_) );
NAND3X1 NAND3X1_13 ( .A(_401_), .B(_403_), .C(_402_), .Y(_404_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_398_) );
AND2X2 AND2X2_13 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_399_) );
OAI21X1 OAI21X1_13 ( .A(_398_), .B(_399_), .C(w_C_23_), .Y(_400_) );
NAND2X1 NAND2X1_26 ( .A(_400_), .B(_404_), .Y(_264__23_) );
INVX1 INVX1_14 ( .A(w_C_24_), .Y(_408_) );
OR2X2 OR2X2_14 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_409_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_410_) );
NAND3X1 NAND3X1_14 ( .A(_408_), .B(_410_), .C(_409_), .Y(_411_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_405_) );
AND2X2 AND2X2_14 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_406_) );
OAI21X1 OAI21X1_14 ( .A(_405_), .B(_406_), .C(w_C_24_), .Y(_407_) );
NAND2X1 NAND2X1_28 ( .A(_407_), .B(_411_), .Y(_264__24_) );
INVX1 INVX1_15 ( .A(w_C_25_), .Y(_415_) );
OR2X2 OR2X2_15 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_416_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_417_) );
NAND3X1 NAND3X1_15 ( .A(_415_), .B(_417_), .C(_416_), .Y(_418_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_412_) );
AND2X2 AND2X2_15 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_413_) );
OAI21X1 OAI21X1_15 ( .A(_412_), .B(_413_), .C(w_C_25_), .Y(_414_) );
NAND2X1 NAND2X1_30 ( .A(_414_), .B(_418_), .Y(_264__25_) );
INVX1 INVX1_16 ( .A(w_C_26_), .Y(_422_) );
OR2X2 OR2X2_16 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_423_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_424_) );
NAND3X1 NAND3X1_16 ( .A(_422_), .B(_424_), .C(_423_), .Y(_425_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_419_) );
AND2X2 AND2X2_16 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_420_) );
OAI21X1 OAI21X1_16 ( .A(_419_), .B(_420_), .C(w_C_26_), .Y(_421_) );
NAND2X1 NAND2X1_32 ( .A(_421_), .B(_425_), .Y(_264__26_) );
INVX1 INVX1_17 ( .A(w_C_27_), .Y(_429_) );
OR2X2 OR2X2_17 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_430_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_431_) );
NAND3X1 NAND3X1_17 ( .A(_429_), .B(_431_), .C(_430_), .Y(_432_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_426_) );
AND2X2 AND2X2_17 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_427_) );
OAI21X1 OAI21X1_17 ( .A(_426_), .B(_427_), .C(w_C_27_), .Y(_428_) );
NAND2X1 NAND2X1_34 ( .A(_428_), .B(_432_), .Y(_264__27_) );
INVX1 INVX1_18 ( .A(w_C_28_), .Y(_436_) );
OR2X2 OR2X2_18 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_437_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_438_) );
NAND3X1 NAND3X1_18 ( .A(_436_), .B(_438_), .C(_437_), .Y(_439_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_433_) );
AND2X2 AND2X2_18 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_434_) );
OAI21X1 OAI21X1_18 ( .A(_433_), .B(_434_), .C(w_C_28_), .Y(_435_) );
NAND2X1 NAND2X1_36 ( .A(_435_), .B(_439_), .Y(_264__28_) );
INVX1 INVX1_19 ( .A(w_C_29_), .Y(_443_) );
OR2X2 OR2X2_19 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_444_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_445_) );
NAND3X1 NAND3X1_19 ( .A(_443_), .B(_445_), .C(_444_), .Y(_446_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_440_) );
AND2X2 AND2X2_19 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_441_) );
OAI21X1 OAI21X1_19 ( .A(_440_), .B(_441_), .C(w_C_29_), .Y(_442_) );
NAND2X1 NAND2X1_38 ( .A(_442_), .B(_446_), .Y(_264__29_) );
INVX1 INVX1_20 ( .A(w_C_30_), .Y(_450_) );
OR2X2 OR2X2_20 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_451_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_452_) );
NAND3X1 NAND3X1_20 ( .A(_450_), .B(_452_), .C(_451_), .Y(_453_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_447_) );
AND2X2 AND2X2_20 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_448_) );
OAI21X1 OAI21X1_20 ( .A(_447_), .B(_448_), .C(w_C_30_), .Y(_449_) );
NAND2X1 NAND2X1_40 ( .A(_449_), .B(_453_), .Y(_264__30_) );
INVX1 INVX1_21 ( .A(w_C_31_), .Y(_457_) );
OR2X2 OR2X2_21 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_458_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_459_) );
NAND3X1 NAND3X1_21 ( .A(_457_), .B(_459_), .C(_458_), .Y(_460_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_454_) );
AND2X2 AND2X2_21 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_455_) );
OAI21X1 OAI21X1_21 ( .A(_454_), .B(_455_), .C(w_C_31_), .Y(_456_) );
NAND2X1 NAND2X1_42 ( .A(_456_), .B(_460_), .Y(_264__31_) );
INVX1 INVX1_22 ( .A(w_C_32_), .Y(_464_) );
OR2X2 OR2X2_22 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_465_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_466_) );
NAND3X1 NAND3X1_22 ( .A(_464_), .B(_466_), .C(_465_), .Y(_467_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_461_) );
AND2X2 AND2X2_22 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_462_) );
OAI21X1 OAI21X1_22 ( .A(_461_), .B(_462_), .C(w_C_32_), .Y(_463_) );
NAND2X1 NAND2X1_44 ( .A(_463_), .B(_467_), .Y(_264__32_) );
INVX1 INVX1_23 ( .A(w_C_33_), .Y(_471_) );
OR2X2 OR2X2_23 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_472_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_473_) );
NAND3X1 NAND3X1_23 ( .A(_471_), .B(_473_), .C(_472_), .Y(_474_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_468_) );
AND2X2 AND2X2_23 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_469_) );
OAI21X1 OAI21X1_23 ( .A(_468_), .B(_469_), .C(w_C_33_), .Y(_470_) );
NAND2X1 NAND2X1_46 ( .A(_470_), .B(_474_), .Y(_264__33_) );
INVX1 INVX1_24 ( .A(w_C_34_), .Y(_478_) );
OR2X2 OR2X2_24 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_479_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_480_) );
NAND3X1 NAND3X1_24 ( .A(_478_), .B(_480_), .C(_479_), .Y(_481_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_475_) );
AND2X2 AND2X2_24 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_476_) );
OAI21X1 OAI21X1_24 ( .A(_475_), .B(_476_), .C(w_C_34_), .Y(_477_) );
NAND2X1 NAND2X1_48 ( .A(_477_), .B(_481_), .Y(_264__34_) );
INVX1 INVX1_25 ( .A(w_C_35_), .Y(_485_) );
OR2X2 OR2X2_25 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_486_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_487_) );
NAND3X1 NAND3X1_25 ( .A(_485_), .B(_487_), .C(_486_), .Y(_488_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_482_) );
AND2X2 AND2X2_25 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_483_) );
OAI21X1 OAI21X1_25 ( .A(_482_), .B(_483_), .C(w_C_35_), .Y(_484_) );
NAND2X1 NAND2X1_50 ( .A(_484_), .B(_488_), .Y(_264__35_) );
INVX1 INVX1_26 ( .A(w_C_36_), .Y(_492_) );
OR2X2 OR2X2_26 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_493_) );
NAND2X1 NAND2X1_51 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_494_) );
NAND3X1 NAND3X1_26 ( .A(_492_), .B(_494_), .C(_493_), .Y(_495_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_489_) );
AND2X2 AND2X2_26 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_490_) );
OAI21X1 OAI21X1_26 ( .A(_489_), .B(_490_), .C(w_C_36_), .Y(_491_) );
NAND2X1 NAND2X1_52 ( .A(_491_), .B(_495_), .Y(_264__36_) );
INVX1 INVX1_27 ( .A(w_C_37_), .Y(_499_) );
OR2X2 OR2X2_27 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_500_) );
NAND2X1 NAND2X1_53 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_501_) );
NAND3X1 NAND3X1_27 ( .A(_499_), .B(_501_), .C(_500_), .Y(_502_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_496_) );
AND2X2 AND2X2_27 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_497_) );
OAI21X1 OAI21X1_27 ( .A(_496_), .B(_497_), .C(w_C_37_), .Y(_498_) );
NAND2X1 NAND2X1_54 ( .A(_498_), .B(_502_), .Y(_264__37_) );
INVX1 INVX1_28 ( .A(w_C_38_), .Y(_506_) );
OR2X2 OR2X2_28 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_507_) );
NAND2X1 NAND2X1_55 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_508_) );
NAND3X1 NAND3X1_28 ( .A(_506_), .B(_508_), .C(_507_), .Y(_509_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_503_) );
AND2X2 AND2X2_28 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_504_) );
OAI21X1 OAI21X1_28 ( .A(_503_), .B(_504_), .C(w_C_38_), .Y(_505_) );
NAND2X1 NAND2X1_56 ( .A(_505_), .B(_509_), .Y(_264__38_) );
INVX1 INVX1_29 ( .A(w_C_39_), .Y(_513_) );
OR2X2 OR2X2_29 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_514_) );
NAND2X1 NAND2X1_57 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_515_) );
NAND3X1 NAND3X1_29 ( .A(_513_), .B(_515_), .C(_514_), .Y(_516_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_510_) );
AND2X2 AND2X2_29 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_511_) );
OAI21X1 OAI21X1_29 ( .A(_510_), .B(_511_), .C(w_C_39_), .Y(_512_) );
NAND2X1 NAND2X1_58 ( .A(_512_), .B(_516_), .Y(_264__39_) );
INVX1 INVX1_30 ( .A(w_C_40_), .Y(_520_) );
OR2X2 OR2X2_30 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_521_) );
NAND2X1 NAND2X1_59 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_522_) );
NAND3X1 NAND3X1_30 ( .A(_520_), .B(_522_), .C(_521_), .Y(_523_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_517_) );
AND2X2 AND2X2_30 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_518_) );
OAI21X1 OAI21X1_30 ( .A(_517_), .B(_518_), .C(w_C_40_), .Y(_519_) );
NAND2X1 NAND2X1_60 ( .A(_519_), .B(_523_), .Y(_264__40_) );
INVX1 INVX1_31 ( .A(w_C_41_), .Y(_527_) );
OR2X2 OR2X2_31 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_528_) );
NAND2X1 NAND2X1_61 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_529_) );
NAND3X1 NAND3X1_31 ( .A(_527_), .B(_529_), .C(_528_), .Y(_530_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_524_) );
AND2X2 AND2X2_31 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_525_) );
OAI21X1 OAI21X1_31 ( .A(_524_), .B(_525_), .C(w_C_41_), .Y(_526_) );
NAND2X1 NAND2X1_62 ( .A(_526_), .B(_530_), .Y(_264__41_) );
INVX1 INVX1_32 ( .A(w_C_42_), .Y(_534_) );
OR2X2 OR2X2_32 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_535_) );
NAND2X1 NAND2X1_63 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_536_) );
NAND3X1 NAND3X1_32 ( .A(_534_), .B(_536_), .C(_535_), .Y(_537_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_531_) );
AND2X2 AND2X2_32 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_532_) );
OAI21X1 OAI21X1_32 ( .A(_531_), .B(_532_), .C(w_C_42_), .Y(_533_) );
NAND2X1 NAND2X1_64 ( .A(_533_), .B(_537_), .Y(_264__42_) );
INVX1 INVX1_33 ( .A(w_C_43_), .Y(_541_) );
OR2X2 OR2X2_33 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_542_) );
NAND2X1 NAND2X1_65 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_543_) );
NAND3X1 NAND3X1_33 ( .A(_541_), .B(_543_), .C(_542_), .Y(_544_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_538_) );
AND2X2 AND2X2_33 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_539_) );
OAI21X1 OAI21X1_33 ( .A(_538_), .B(_539_), .C(w_C_43_), .Y(_540_) );
NAND2X1 NAND2X1_66 ( .A(_540_), .B(_544_), .Y(_264__43_) );
INVX1 INVX1_34 ( .A(w_C_44_), .Y(_548_) );
OR2X2 OR2X2_34 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_549_) );
NAND2X1 NAND2X1_67 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_550_) );
NAND3X1 NAND3X1_34 ( .A(_548_), .B(_550_), .C(_549_), .Y(_551_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_545_) );
AND2X2 AND2X2_34 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_546_) );
OAI21X1 OAI21X1_34 ( .A(_545_), .B(_546_), .C(w_C_44_), .Y(_547_) );
NAND2X1 NAND2X1_68 ( .A(_547_), .B(_551_), .Y(_264__44_) );
INVX1 INVX1_35 ( .A(w_C_45_), .Y(_555_) );
OR2X2 OR2X2_35 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_556_) );
NAND2X1 NAND2X1_69 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_557_) );
NAND3X1 NAND3X1_35 ( .A(_555_), .B(_557_), .C(_556_), .Y(_558_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_552_) );
AND2X2 AND2X2_35 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_553_) );
OAI21X1 OAI21X1_35 ( .A(_552_), .B(_553_), .C(w_C_45_), .Y(_554_) );
NAND2X1 NAND2X1_70 ( .A(_554_), .B(_558_), .Y(_264__45_) );
INVX1 INVX1_36 ( .A(1'b0), .Y(_562_) );
OR2X2 OR2X2_36 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_563_) );
NAND2X1 NAND2X1_71 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_564_) );
NAND3X1 NAND3X1_36 ( .A(_562_), .B(_564_), .C(_563_), .Y(_565_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_559_) );
AND2X2 AND2X2_36 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_560_) );
OAI21X1 OAI21X1_36 ( .A(_559_), .B(_560_), .C(1'b0), .Y(_561_) );
NAND2X1 NAND2X1_72 ( .A(_561_), .B(_565_), .Y(_264__0_) );
INVX1 INVX1_37 ( .A(w_C_1_), .Y(_569_) );
OR2X2 OR2X2_37 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_570_) );
NAND2X1 NAND2X1_73 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_571_) );
NAND3X1 NAND3X1_37 ( .A(_569_), .B(_571_), .C(_570_), .Y(_572_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_566_) );
AND2X2 AND2X2_37 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_567_) );
OAI21X1 OAI21X1_37 ( .A(_566_), .B(_567_), .C(w_C_1_), .Y(_568_) );
NAND2X1 NAND2X1_74 ( .A(_568_), .B(_572_), .Y(_264__1_) );
INVX1 INVX1_38 ( .A(w_C_2_), .Y(_576_) );
OR2X2 OR2X2_38 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_577_) );
NAND2X1 NAND2X1_75 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_578_) );
NAND3X1 NAND3X1_38 ( .A(_576_), .B(_578_), .C(_577_), .Y(_579_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_573_) );
AND2X2 AND2X2_38 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_574_) );
OAI21X1 OAI21X1_38 ( .A(_573_), .B(_574_), .C(w_C_2_), .Y(_575_) );
NAND2X1 NAND2X1_76 ( .A(_575_), .B(_579_), .Y(_264__2_) );
INVX1 INVX1_39 ( .A(w_C_3_), .Y(_583_) );
OR2X2 OR2X2_39 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_584_) );
NAND2X1 NAND2X1_77 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_585_) );
NAND3X1 NAND3X1_39 ( .A(_583_), .B(_585_), .C(_584_), .Y(_586_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_580_) );
AND2X2 AND2X2_39 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_581_) );
OAI21X1 OAI21X1_39 ( .A(_580_), .B(_581_), .C(w_C_3_), .Y(_582_) );
NAND2X1 NAND2X1_78 ( .A(_582_), .B(_586_), .Y(_264__3_) );
INVX1 INVX1_40 ( .A(_240_), .Y(w_C_41_) );
INVX1 INVX1_41 ( .A(i_add2[41]), .Y(_241_) );
INVX1 INVX1_42 ( .A(i_add1[41]), .Y(_242_) );
OAI21X1 OAI21X1_40 ( .A(_241_), .B(_242_), .C(_240_), .Y(_243_) );
OAI21X1 OAI21X1_41 ( .A(i_add2[41]), .B(i_add1[41]), .C(_243_), .Y(_244_) );
INVX1 INVX1_43 ( .A(_244_), .Y(w_C_42_) );
NAND2X1 NAND2X1_79 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_245_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_246_) );
OAI21X1 OAI21X1_42 ( .A(_246_), .B(_244_), .C(_245_), .Y(w_C_43_) );
NAND2X1 NAND2X1_80 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_247_) );
INVX1 INVX1_44 ( .A(_246_), .Y(_248_) );
NOR2X1 NOR2X1_41 ( .A(_241_), .B(_242_), .Y(_249_) );
INVX1 INVX1_45 ( .A(_249_), .Y(_250_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_251_) );
INVX1 INVX1_46 ( .A(_251_), .Y(_252_) );
NAND2X1 NAND2X1_81 ( .A(_241_), .B(_242_), .Y(_253_) );
NAND3X1 NAND3X1_40 ( .A(_252_), .B(_253_), .C(_239_), .Y(_254_) );
NAND3X1 NAND3X1_41 ( .A(_250_), .B(_245_), .C(_254_), .Y(_255_) );
OR2X2 OR2X2_40 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_256_) );
NAND3X1 NAND3X1_42 ( .A(_248_), .B(_256_), .C(_255_), .Y(_257_) );
NAND2X1 NAND2X1_82 ( .A(_247_), .B(_257_), .Y(w_C_44_) );
OR2X2 OR2X2_41 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_258_) );
NAND2X1 NAND2X1_83 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_259_) );
NAND3X1 NAND3X1_43 ( .A(_247_), .B(_259_), .C(_257_), .Y(_260_) );
AND2X2 AND2X2_40 ( .A(_260_), .B(_258_), .Y(w_C_45_) );
NAND2X1 NAND2X1_84 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_261_) );
OR2X2 OR2X2_42 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_262_) );
NAND3X1 NAND3X1_44 ( .A(_258_), .B(_262_), .C(_260_), .Y(_263_) );
NAND2X1 NAND2X1_85 ( .A(_261_), .B(_263_), .Y(w_C_46_) );
NAND2X1 NAND2X1_86 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_47 ( .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_44 ( .A(_1_), .B(_2_), .Y(w_C_2_) );
INVX1 INVX1_48 ( .A(i_add2[2]), .Y(_3_) );
INVX1 INVX1_49 ( .A(i_add1[2]), .Y(_4_) );
NAND2X1 NAND2X1_87 ( .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_88 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
OAI21X1 OAI21X1_43 ( .A(_1_), .B(_2_), .C(_6_), .Y(_7_) );
AND2X2 AND2X2_41 ( .A(_7_), .B(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_89 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
OR2X2 OR2X2_43 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_45 ( .A(_5_), .B(_9_), .C(_7_), .Y(_10_) );
AND2X2 AND2X2_42 ( .A(_10_), .B(_8_), .Y(_11_) );
INVX1 INVX1_50 ( .A(_11_), .Y(w_C_4_) );
NAND2X1 NAND2X1_90 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_12_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
OAI21X1 OAI21X1_44 ( .A(_13_), .B(_11_), .C(_12_), .Y(w_C_5_) );
AND2X2 AND2X2_43 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_14_) );
INVX1 INVX1_51 ( .A(_14_), .Y(_15_) );
INVX1 INVX1_52 ( .A(_13_), .Y(_16_) );
NAND3X1 NAND3X1_46 ( .A(_8_), .B(_12_), .C(_10_), .Y(_17_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_18_) );
INVX1 INVX1_53 ( .A(_18_), .Y(_19_) );
NAND3X1 NAND3X1_47 ( .A(_16_), .B(_19_), .C(_17_), .Y(_20_) );
AND2X2 AND2X2_44 ( .A(_20_), .B(_15_), .Y(_21_) );
INVX1 INVX1_54 ( .A(_21_), .Y(w_C_6_) );
AND2X2 AND2X2_45 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_55 ( .A(_22_), .Y(_23_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_24_) );
OAI21X1 OAI21X1_45 ( .A(_24_), .B(_21_), .C(_23_), .Y(w_C_7_) );
AND2X2 AND2X2_46 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_25_) );
INVX1 INVX1_56 ( .A(_25_), .Y(_26_) );
INVX1 INVX1_57 ( .A(_24_), .Y(_27_) );
NAND3X1 NAND3X1_48 ( .A(_15_), .B(_23_), .C(_20_), .Y(_28_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_29_) );
INVX1 INVX1_58 ( .A(_29_), .Y(_30_) );
NAND3X1 NAND3X1_49 ( .A(_27_), .B(_30_), .C(_28_), .Y(_31_) );
AND2X2 AND2X2_47 ( .A(_31_), .B(_26_), .Y(_32_) );
INVX1 INVX1_59 ( .A(_32_), .Y(w_C_8_) );
AND2X2 AND2X2_48 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_33_) );
INVX1 INVX1_60 ( .A(_33_), .Y(_34_) );
NAND3X1 NAND3X1_50 ( .A(_26_), .B(_34_), .C(_31_), .Y(_35_) );
OAI21X1 OAI21X1_46 ( .A(i_add2[8]), .B(i_add1[8]), .C(_35_), .Y(_36_) );
INVX1 INVX1_61 ( .A(_36_), .Y(w_C_9_) );
INVX1 INVX1_62 ( .A(i_add2[9]), .Y(_37_) );
INVX1 INVX1_63 ( .A(i_add1[9]), .Y(_38_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_39_) );
INVX1 INVX1_64 ( .A(_39_), .Y(_40_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_41_) );
INVX1 INVX1_65 ( .A(_41_), .Y(_42_) );
NAND3X1 NAND3X1_51 ( .A(_40_), .B(_42_), .C(_35_), .Y(_43_) );
OAI21X1 OAI21X1_47 ( .A(_37_), .B(_38_), .C(_43_), .Y(w_C_10_) );
NOR2X1 NOR2X1_51 ( .A(_37_), .B(_38_), .Y(_44_) );
INVX1 INVX1_66 ( .A(_44_), .Y(_45_) );
AND2X2 AND2X2_49 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_46_) );
INVX1 INVX1_67 ( .A(_46_), .Y(_47_) );
NAND3X1 NAND3X1_52 ( .A(_45_), .B(_47_), .C(_43_), .Y(_48_) );
OAI21X1 OAI21X1_48 ( .A(i_add2[10]), .B(i_add1[10]), .C(_48_), .Y(_49_) );
INVX1 INVX1_68 ( .A(_49_), .Y(w_C_11_) );
INVX1 INVX1_69 ( .A(i_add2[11]), .Y(_50_) );
INVX1 INVX1_70 ( .A(i_add1[11]), .Y(_51_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_52_) );
INVX1 INVX1_71 ( .A(_52_), .Y(_53_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_54_) );
INVX1 INVX1_72 ( .A(_54_), .Y(_55_) );
NAND3X1 NAND3X1_53 ( .A(_53_), .B(_55_), .C(_48_), .Y(_56_) );
OAI21X1 OAI21X1_49 ( .A(_50_), .B(_51_), .C(_56_), .Y(w_C_12_) );
NOR2X1 NOR2X1_54 ( .A(_50_), .B(_51_), .Y(_57_) );
INVX1 INVX1_73 ( .A(_57_), .Y(_58_) );
AND2X2 AND2X2_50 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_59_) );
INVX1 INVX1_74 ( .A(_59_), .Y(_60_) );
NAND3X1 NAND3X1_54 ( .A(_58_), .B(_60_), .C(_56_), .Y(_61_) );
OAI21X1 OAI21X1_50 ( .A(i_add2[12]), .B(i_add1[12]), .C(_61_), .Y(_62_) );
INVX1 INVX1_75 ( .A(_62_), .Y(w_C_13_) );
INVX1 INVX1_76 ( .A(i_add2[13]), .Y(_63_) );
INVX1 INVX1_77 ( .A(i_add1[13]), .Y(_64_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_65_) );
INVX1 INVX1_78 ( .A(_65_), .Y(_66_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_67_) );
INVX1 INVX1_79 ( .A(_67_), .Y(_68_) );
NAND3X1 NAND3X1_55 ( .A(_66_), .B(_68_), .C(_61_), .Y(_69_) );
OAI21X1 OAI21X1_51 ( .A(_63_), .B(_64_), .C(_69_), .Y(w_C_14_) );
NOR2X1 NOR2X1_57 ( .A(_63_), .B(_64_), .Y(_70_) );
INVX1 INVX1_80 ( .A(_70_), .Y(_71_) );
AND2X2 AND2X2_51 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_72_) );
INVX1 INVX1_81 ( .A(_72_), .Y(_73_) );
NAND3X1 NAND3X1_56 ( .A(_71_), .B(_73_), .C(_69_), .Y(_74_) );
OAI21X1 OAI21X1_52 ( .A(i_add2[14]), .B(i_add1[14]), .C(_74_), .Y(_75_) );
INVX1 INVX1_82 ( .A(_75_), .Y(w_C_15_) );
INVX1 INVX1_83 ( .A(i_add2[15]), .Y(_76_) );
INVX1 INVX1_84 ( .A(i_add1[15]), .Y(_77_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_78_) );
INVX1 INVX1_85 ( .A(_78_), .Y(_79_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_80_) );
INVX1 INVX1_86 ( .A(_80_), .Y(_81_) );
NAND3X1 NAND3X1_57 ( .A(_79_), .B(_81_), .C(_74_), .Y(_82_) );
OAI21X1 OAI21X1_53 ( .A(_76_), .B(_77_), .C(_82_), .Y(w_C_16_) );
NOR2X1 NOR2X1_60 ( .A(_76_), .B(_77_), .Y(_83_) );
INVX1 INVX1_87 ( .A(_83_), .Y(_84_) );
AND2X2 AND2X2_52 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_85_) );
INVX1 INVX1_88 ( .A(_85_), .Y(_86_) );
NAND3X1 NAND3X1_58 ( .A(_84_), .B(_86_), .C(_82_), .Y(_87_) );
OAI21X1 OAI21X1_54 ( .A(i_add2[16]), .B(i_add1[16]), .C(_87_), .Y(_88_) );
INVX1 INVX1_89 ( .A(_88_), .Y(w_C_17_) );
INVX1 INVX1_90 ( .A(i_add2[17]), .Y(_89_) );
INVX1 INVX1_91 ( .A(i_add1[17]), .Y(_90_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_91_) );
INVX1 INVX1_92 ( .A(_91_), .Y(_92_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_93_) );
INVX1 INVX1_93 ( .A(_93_), .Y(_94_) );
NAND3X1 NAND3X1_59 ( .A(_92_), .B(_94_), .C(_87_), .Y(_95_) );
OAI21X1 OAI21X1_55 ( .A(_89_), .B(_90_), .C(_95_), .Y(w_C_18_) );
NOR2X1 NOR2X1_63 ( .A(_89_), .B(_90_), .Y(_96_) );
INVX1 INVX1_94 ( .A(_96_), .Y(_97_) );
AND2X2 AND2X2_53 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_98_) );
INVX1 INVX1_95 ( .A(_98_), .Y(_99_) );
NAND3X1 NAND3X1_60 ( .A(_97_), .B(_99_), .C(_95_), .Y(_100_) );
OAI21X1 OAI21X1_56 ( .A(i_add2[18]), .B(i_add1[18]), .C(_100_), .Y(_101_) );
INVX1 INVX1_96 ( .A(_101_), .Y(w_C_19_) );
INVX1 INVX1_97 ( .A(i_add2[19]), .Y(_102_) );
INVX1 INVX1_98 ( .A(i_add1[19]), .Y(_103_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_104_) );
INVX1 INVX1_99 ( .A(_104_), .Y(_105_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_106_) );
INVX1 INVX1_100 ( .A(_106_), .Y(_107_) );
NAND3X1 NAND3X1_61 ( .A(_105_), .B(_107_), .C(_100_), .Y(_108_) );
OAI21X1 OAI21X1_57 ( .A(_102_), .B(_103_), .C(_108_), .Y(w_C_20_) );
NOR2X1 NOR2X1_66 ( .A(_102_), .B(_103_), .Y(_109_) );
INVX1 INVX1_101 ( .A(_109_), .Y(_110_) );
AND2X2 AND2X2_54 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_111_) );
INVX1 INVX1_102 ( .A(_111_), .Y(_112_) );
NAND3X1 NAND3X1_62 ( .A(_110_), .B(_112_), .C(_108_), .Y(_113_) );
OAI21X1 OAI21X1_58 ( .A(i_add2[20]), .B(i_add1[20]), .C(_113_), .Y(_114_) );
INVX1 INVX1_103 ( .A(_114_), .Y(w_C_21_) );
INVX1 INVX1_104 ( .A(i_add2[21]), .Y(_115_) );
INVX1 INVX1_105 ( .A(i_add1[21]), .Y(_116_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_117_) );
INVX1 INVX1_106 ( .A(_117_), .Y(_118_) );
NOR2X1 NOR2X1_68 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_119_) );
INVX1 INVX1_107 ( .A(_119_), .Y(_120_) );
NAND3X1 NAND3X1_63 ( .A(_118_), .B(_120_), .C(_113_), .Y(_121_) );
OAI21X1 OAI21X1_59 ( .A(_115_), .B(_116_), .C(_121_), .Y(w_C_22_) );
NOR2X1 NOR2X1_69 ( .A(_115_), .B(_116_), .Y(_122_) );
INVX1 INVX1_108 ( .A(_122_), .Y(_123_) );
AND2X2 AND2X2_55 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_124_) );
INVX1 INVX1_109 ( .A(_124_), .Y(_125_) );
NAND3X1 NAND3X1_64 ( .A(_123_), .B(_125_), .C(_121_), .Y(_126_) );
OAI21X1 OAI21X1_60 ( .A(i_add2[22]), .B(i_add1[22]), .C(_126_), .Y(_127_) );
INVX1 INVX1_110 ( .A(_127_), .Y(w_C_23_) );
INVX1 INVX1_111 ( .A(i_add2[23]), .Y(_128_) );
INVX1 INVX1_112 ( .A(i_add1[23]), .Y(_129_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_130_) );
INVX1 INVX1_113 ( .A(_130_), .Y(_131_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_132_) );
INVX1 INVX1_114 ( .A(_132_), .Y(_133_) );
NAND3X1 NAND3X1_65 ( .A(_131_), .B(_133_), .C(_126_), .Y(_134_) );
OAI21X1 OAI21X1_61 ( .A(_128_), .B(_129_), .C(_134_), .Y(w_C_24_) );
NOR2X1 NOR2X1_72 ( .A(_128_), .B(_129_), .Y(_135_) );
INVX1 INVX1_115 ( .A(_135_), .Y(_136_) );
AND2X2 AND2X2_56 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_137_) );
INVX1 INVX1_116 ( .A(_137_), .Y(_138_) );
NAND3X1 NAND3X1_66 ( .A(_136_), .B(_138_), .C(_134_), .Y(_139_) );
OAI21X1 OAI21X1_62 ( .A(i_add2[24]), .B(i_add1[24]), .C(_139_), .Y(_140_) );
INVX1 INVX1_117 ( .A(_140_), .Y(w_C_25_) );
INVX1 INVX1_118 ( .A(i_add2[25]), .Y(_141_) );
INVX1 INVX1_119 ( .A(i_add1[25]), .Y(_142_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_143_) );
INVX1 INVX1_120 ( .A(_143_), .Y(_144_) );
NOR2X1 NOR2X1_74 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_145_) );
INVX1 INVX1_121 ( .A(_145_), .Y(_146_) );
NAND3X1 NAND3X1_67 ( .A(_144_), .B(_146_), .C(_139_), .Y(_147_) );
OAI21X1 OAI21X1_63 ( .A(_141_), .B(_142_), .C(_147_), .Y(w_C_26_) );
NOR2X1 NOR2X1_75 ( .A(_141_), .B(_142_), .Y(_148_) );
INVX1 INVX1_122 ( .A(_148_), .Y(_149_) );
AND2X2 AND2X2_57 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_150_) );
INVX1 INVX1_123 ( .A(_150_), .Y(_151_) );
NAND3X1 NAND3X1_68 ( .A(_149_), .B(_151_), .C(_147_), .Y(_152_) );
OAI21X1 OAI21X1_64 ( .A(i_add2[26]), .B(i_add1[26]), .C(_152_), .Y(_153_) );
INVX1 INVX1_124 ( .A(_153_), .Y(w_C_27_) );
INVX1 INVX1_125 ( .A(i_add2[27]), .Y(_154_) );
INVX1 INVX1_126 ( .A(i_add1[27]), .Y(_155_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_156_) );
INVX1 INVX1_127 ( .A(_156_), .Y(_157_) );
NOR2X1 NOR2X1_77 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_158_) );
INVX1 INVX1_128 ( .A(_158_), .Y(_159_) );
NAND3X1 NAND3X1_69 ( .A(_157_), .B(_159_), .C(_152_), .Y(_160_) );
OAI21X1 OAI21X1_65 ( .A(_154_), .B(_155_), .C(_160_), .Y(w_C_28_) );
NOR2X1 NOR2X1_78 ( .A(_154_), .B(_155_), .Y(_161_) );
INVX1 INVX1_129 ( .A(_161_), .Y(_162_) );
AND2X2 AND2X2_58 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_163_) );
INVX1 INVX1_130 ( .A(_163_), .Y(_164_) );
NAND3X1 NAND3X1_70 ( .A(_162_), .B(_164_), .C(_160_), .Y(_165_) );
OAI21X1 OAI21X1_66 ( .A(i_add2[28]), .B(i_add1[28]), .C(_165_), .Y(_166_) );
INVX1 INVX1_131 ( .A(_166_), .Y(w_C_29_) );
INVX1 INVX1_132 ( .A(i_add2[29]), .Y(_167_) );
INVX1 INVX1_133 ( .A(i_add1[29]), .Y(_168_) );
NOR2X1 NOR2X1_79 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_169_) );
INVX1 INVX1_134 ( .A(_169_), .Y(_170_) );
NOR2X1 NOR2X1_80 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_171_) );
INVX1 INVX1_135 ( .A(_171_), .Y(_172_) );
NAND3X1 NAND3X1_71 ( .A(_170_), .B(_172_), .C(_165_), .Y(_173_) );
OAI21X1 OAI21X1_67 ( .A(_167_), .B(_168_), .C(_173_), .Y(w_C_30_) );
NOR2X1 NOR2X1_81 ( .A(_167_), .B(_168_), .Y(_174_) );
INVX1 INVX1_136 ( .A(_174_), .Y(_175_) );
AND2X2 AND2X2_59 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_176_) );
INVX1 INVX1_137 ( .A(_176_), .Y(_177_) );
NAND3X1 NAND3X1_72 ( .A(_175_), .B(_177_), .C(_173_), .Y(_178_) );
OAI21X1 OAI21X1_68 ( .A(i_add2[30]), .B(i_add1[30]), .C(_178_), .Y(_179_) );
INVX1 INVX1_138 ( .A(_179_), .Y(w_C_31_) );
INVX1 INVX1_139 ( .A(i_add2[31]), .Y(_180_) );
INVX1 INVX1_140 ( .A(i_add1[31]), .Y(_181_) );
NOR2X1 NOR2X1_82 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_182_) );
INVX1 INVX1_141 ( .A(_182_), .Y(_183_) );
NOR2X1 NOR2X1_83 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_184_) );
INVX1 INVX1_142 ( .A(_184_), .Y(_185_) );
NAND3X1 NAND3X1_73 ( .A(_183_), .B(_185_), .C(_178_), .Y(_186_) );
OAI21X1 OAI21X1_69 ( .A(_180_), .B(_181_), .C(_186_), .Y(w_C_32_) );
NOR2X1 NOR2X1_84 ( .A(_180_), .B(_181_), .Y(_187_) );
INVX1 INVX1_143 ( .A(_187_), .Y(_188_) );
AND2X2 AND2X2_60 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_189_) );
INVX1 INVX1_144 ( .A(_189_), .Y(_190_) );
NAND3X1 NAND3X1_74 ( .A(_188_), .B(_190_), .C(_186_), .Y(_191_) );
OAI21X1 OAI21X1_70 ( .A(i_add2[32]), .B(i_add1[32]), .C(_191_), .Y(_192_) );
INVX1 INVX1_145 ( .A(_192_), .Y(w_C_33_) );
INVX1 INVX1_146 ( .A(i_add2[33]), .Y(_193_) );
INVX1 INVX1_147 ( .A(i_add1[33]), .Y(_194_) );
NOR2X1 NOR2X1_85 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_195_) );
INVX1 INVX1_148 ( .A(_195_), .Y(_196_) );
NOR2X1 NOR2X1_86 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_197_) );
INVX1 INVX1_149 ( .A(_197_), .Y(_198_) );
NAND3X1 NAND3X1_75 ( .A(_196_), .B(_198_), .C(_191_), .Y(_199_) );
OAI21X1 OAI21X1_71 ( .A(_193_), .B(_194_), .C(_199_), .Y(w_C_34_) );
NOR2X1 NOR2X1_87 ( .A(_193_), .B(_194_), .Y(_200_) );
INVX1 INVX1_150 ( .A(_200_), .Y(_201_) );
AND2X2 AND2X2_61 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_202_) );
INVX1 INVX1_151 ( .A(_202_), .Y(_203_) );
NAND3X1 NAND3X1_76 ( .A(_201_), .B(_203_), .C(_199_), .Y(_204_) );
OAI21X1 OAI21X1_72 ( .A(i_add2[34]), .B(i_add1[34]), .C(_204_), .Y(_205_) );
INVX1 INVX1_152 ( .A(_205_), .Y(w_C_35_) );
INVX1 INVX1_153 ( .A(i_add2[35]), .Y(_206_) );
INVX1 INVX1_154 ( .A(i_add1[35]), .Y(_207_) );
NOR2X1 NOR2X1_88 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_208_) );
INVX1 INVX1_155 ( .A(_208_), .Y(_209_) );
NOR2X1 NOR2X1_89 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_210_) );
INVX1 INVX1_156 ( .A(_210_), .Y(_211_) );
NAND3X1 NAND3X1_77 ( .A(_209_), .B(_211_), .C(_204_), .Y(_212_) );
OAI21X1 OAI21X1_73 ( .A(_206_), .B(_207_), .C(_212_), .Y(w_C_36_) );
NOR2X1 NOR2X1_90 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_213_) );
INVX1 INVX1_157 ( .A(_213_), .Y(_214_) );
NOR2X1 NOR2X1_91 ( .A(_206_), .B(_207_), .Y(_215_) );
INVX1 INVX1_158 ( .A(_215_), .Y(_216_) );
NAND2X1 NAND2X1_91 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_217_) );
NAND3X1 NAND3X1_78 ( .A(_216_), .B(_217_), .C(_212_), .Y(_218_) );
AND2X2 AND2X2_62 ( .A(_218_), .B(_214_), .Y(w_C_37_) );
INVX1 INVX1_159 ( .A(i_add2[37]), .Y(_219_) );
INVX1 INVX1_160 ( .A(i_add1[37]), .Y(_220_) );
NAND2X1 NAND2X1_92 ( .A(_219_), .B(_220_), .Y(_221_) );
NAND3X1 NAND3X1_79 ( .A(_214_), .B(_221_), .C(_218_), .Y(_222_) );
OAI21X1 OAI21X1_74 ( .A(_219_), .B(_220_), .C(_222_), .Y(w_C_38_) );
INVX1 INVX1_161 ( .A(i_add2[38]), .Y(_223_) );
INVX1 INVX1_162 ( .A(i_add1[38]), .Y(_224_) );
OAI21X1 OAI21X1_75 ( .A(i_add2[38]), .B(i_add1[38]), .C(w_C_38_), .Y(_225_) );
OAI21X1 OAI21X1_76 ( .A(_223_), .B(_224_), .C(_225_), .Y(w_C_39_) );
INVX1 INVX1_163 ( .A(i_add2[39]), .Y(_226_) );
INVX1 INVX1_164 ( .A(i_add1[39]), .Y(_227_) );
NOR2X1 NOR2X1_92 ( .A(_226_), .B(_227_), .Y(_228_) );
OR2X2 OR2X2_44 ( .A(w_C_39_), .B(_228_), .Y(_229_) );
OAI21X1 OAI21X1_77 ( .A(i_add2[39]), .B(i_add1[39]), .C(_229_), .Y(_230_) );
INVX1 INVX1_165 ( .A(_230_), .Y(w_C_40_) );
INVX1 INVX1_166 ( .A(_228_), .Y(_231_) );
NAND2X1 NAND2X1_93 ( .A(_223_), .B(_224_), .Y(_232_) );
NAND2X1 NAND2X1_94 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_233_) );
NAND2X1 NAND2X1_95 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_234_) );
NAND3X1 NAND3X1_80 ( .A(_233_), .B(_234_), .C(_222_), .Y(_235_) );
NAND2X1 NAND2X1_96 ( .A(_226_), .B(_227_), .Y(_236_) );
NAND3X1 NAND3X1_81 ( .A(_232_), .B(_236_), .C(_235_), .Y(_237_) );
NAND2X1 NAND2X1_97 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_238_) );
NAND3X1 NAND3X1_82 ( .A(_231_), .B(_238_), .C(_237_), .Y(_239_) );
OAI21X1 OAI21X1_78 ( .A(i_add2[40]), .B(i_add1[40]), .C(_239_), .Y(_240_) );
BUFX2 BUFX2_1 ( .A(_264__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_264__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_264__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_264__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_264__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_264__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_264__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_264__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_264__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_264__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_264__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_264__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_264__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_264__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_264__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_264__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_264__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_264__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_264__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_264__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_264__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_264__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_264__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_264__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_264__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_264__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_264__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_264__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_264__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_264__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_264__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_264__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_264__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_264__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_264__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_264__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_264__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(_264__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .A(_264__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .A(_264__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .A(_264__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .A(_264__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .A(_264__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .A(_264__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .A(_264__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .A(_264__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .A(w_C_46_), .Y(o_result[46]) );
INVX1 INVX1_167 ( .A(w_C_4_), .Y(_268_) );
OR2X2 OR2X2_45 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_269_) );
NAND2X1 NAND2X1_98 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_270_) );
NAND3X1 NAND3X1_83 ( .A(_268_), .B(_270_), .C(_269_), .Y(_271_) );
NOR2X1 NOR2X1_93 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_265_) );
AND2X2 AND2X2_63 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_266_) );
OAI21X1 OAI21X1_79 ( .A(_265_), .B(_266_), .C(w_C_4_), .Y(_267_) );
NAND2X1 NAND2X1_99 ( .A(_267_), .B(_271_), .Y(_264__4_) );
INVX1 INVX1_168 ( .A(w_C_5_), .Y(_275_) );
OR2X2 OR2X2_46 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_276_) );
NAND2X1 NAND2X1_100 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_277_) );
NAND3X1 NAND3X1_84 ( .A(_275_), .B(_277_), .C(_276_), .Y(_278_) );
NOR2X1 NOR2X1_94 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_272_) );
AND2X2 AND2X2_64 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_273_) );
OAI21X1 OAI21X1_80 ( .A(_272_), .B(_273_), .C(w_C_5_), .Y(_274_) );
NAND2X1 NAND2X1_101 ( .A(_274_), .B(_278_), .Y(_264__5_) );
INVX1 INVX1_169 ( .A(w_C_6_), .Y(_282_) );
OR2X2 OR2X2_47 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_283_) );
NAND2X1 NAND2X1_102 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_284_) );
NAND3X1 NAND3X1_85 ( .A(_282_), .B(_284_), .C(_283_), .Y(_285_) );
NOR2X1 NOR2X1_95 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_279_) );
AND2X2 AND2X2_65 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_280_) );
OAI21X1 OAI21X1_81 ( .A(_279_), .B(_280_), .C(w_C_6_), .Y(_281_) );
NAND2X1 NAND2X1_103 ( .A(_281_), .B(_285_), .Y(_264__6_) );
INVX1 INVX1_170 ( .A(w_C_7_), .Y(_289_) );
OR2X2 OR2X2_48 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_290_) );
NAND2X1 NAND2X1_104 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_291_) );
NAND3X1 NAND3X1_86 ( .A(_289_), .B(_291_), .C(_290_), .Y(_292_) );
NOR2X1 NOR2X1_96 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_286_) );
AND2X2 AND2X2_66 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_287_) );
OAI21X1 OAI21X1_82 ( .A(_286_), .B(_287_), .C(w_C_7_), .Y(_288_) );
NAND2X1 NAND2X1_105 ( .A(_288_), .B(_292_), .Y(_264__7_) );
INVX1 INVX1_171 ( .A(w_C_8_), .Y(_296_) );
OR2X2 OR2X2_49 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_297_) );
NAND2X1 NAND2X1_106 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_298_) );
NAND3X1 NAND3X1_87 ( .A(_296_), .B(_298_), .C(_297_), .Y(_299_) );
NOR2X1 NOR2X1_97 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_293_) );
AND2X2 AND2X2_67 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_294_) );
OAI21X1 OAI21X1_83 ( .A(_293_), .B(_294_), .C(w_C_8_), .Y(_295_) );
NAND2X1 NAND2X1_107 ( .A(_295_), .B(_299_), .Y(_264__8_) );
INVX1 INVX1_172 ( .A(w_C_9_), .Y(_303_) );
OR2X2 OR2X2_50 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_304_) );
NAND2X1 NAND2X1_108 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_305_) );
NAND3X1 NAND3X1_88 ( .A(_303_), .B(_305_), .C(_304_), .Y(_306_) );
NOR2X1 NOR2X1_98 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_300_) );
AND2X2 AND2X2_68 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_301_) );
OAI21X1 OAI21X1_84 ( .A(_300_), .B(_301_), .C(w_C_9_), .Y(_302_) );
NAND2X1 NAND2X1_109 ( .A(_302_), .B(_306_), .Y(_264__9_) );
INVX1 INVX1_173 ( .A(w_C_10_), .Y(_310_) );
OR2X2 OR2X2_51 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_311_) );
NAND2X1 NAND2X1_110 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_312_) );
NAND3X1 NAND3X1_89 ( .A(_310_), .B(_312_), .C(_311_), .Y(_313_) );
NOR2X1 NOR2X1_99 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_307_) );
AND2X2 AND2X2_69 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_308_) );
OAI21X1 OAI21X1_85 ( .A(_307_), .B(_308_), .C(w_C_10_), .Y(_309_) );
NAND2X1 NAND2X1_111 ( .A(_309_), .B(_313_), .Y(_264__10_) );
BUFX2 BUFX2_48 ( .A(w_C_46_), .Y(_264__46_) );
BUFX2 BUFX2_49 ( .A(1'b0), .Y(w_C_0_) );
endmodule
