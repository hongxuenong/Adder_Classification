module CSkipA_31bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_7_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_15_) );
OAI21X1 OAI21X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .C(1'b0), .Y(_16_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_17_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_18_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_19_) );
NAND3X1 NAND3X1_1 ( .A(_17_), .B(_18_), .C(_19_), .Y(_20_) );
OAI21X1 OAI21X1_2 ( .A(_16_), .B(_20_), .C(_15_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3_), .Y(_21_) );
OAI21X1 OAI21X1_3 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .C(1'b0), .Y(_22_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_23_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_24_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_25_) );
NAND3X1 NAND3X1_2 ( .A(_23_), .B(_24_), .C(_25_), .Y(_26_) );
OAI21X1 OAI21X1_4 ( .A(_22_), .B(_26_), .C(_21_), .Y(w_cout_2_) );
INVX1 INVX1_3 ( .A(_5_), .Y(_27_) );
OAI21X1 OAI21X1_5 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .C(1'b0), .Y(_28_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_29_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_30_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_31_) );
NAND3X1 NAND3X1_3 ( .A(_29_), .B(_30_), .C(_31_), .Y(_32_) );
OAI21X1 OAI21X1_6 ( .A(_28_), .B(_32_), .C(_27_), .Y(w_cout_3_) );
INVX1 INVX1_4 ( .A(_7_), .Y(_33_) );
OAI21X1 OAI21X1_7 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .C(1'b0), .Y(_34_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_35_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_36_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_37_) );
NAND3X1 NAND3X1_4 ( .A(_35_), .B(_36_), .C(_37_), .Y(_38_) );
OAI21X1 OAI21X1_8 ( .A(_34_), .B(_38_), .C(_33_), .Y(w_cout_4_) );
INVX1 INVX1_5 ( .A(_9_), .Y(_39_) );
OAI21X1 OAI21X1_9 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .C(1'b0), .Y(_40_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_41_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_42_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_43_) );
NAND3X1 NAND3X1_5 ( .A(_41_), .B(_42_), .C(_43_), .Y(_44_) );
OAI21X1 OAI21X1_10 ( .A(_40_), .B(_44_), .C(_39_), .Y(w_cout_5_) );
INVX1 INVX1_6 ( .A(_11_), .Y(_45_) );
OAI21X1 OAI21X1_11 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .C(1'b0), .Y(_46_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_47_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_48_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_49_) );
NAND3X1 NAND3X1_6 ( .A(_47_), .B(_48_), .C(_49_), .Y(_50_) );
OAI21X1 OAI21X1_12 ( .A(_46_), .B(_50_), .C(_45_), .Y(w_cout_6_) );
INVX1 INVX1_7 ( .A(_13_), .Y(_51_) );
OAI21X1 OAI21X1_13 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .C(1'b0), .Y(_52_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_53_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_54_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_55_) );
NAND3X1 NAND3X1_7 ( .A(_53_), .B(_54_), .C(_55_), .Y(_56_) );
OAI21X1 OAI21X1_14 ( .A(_52_), .B(_56_), .C(_51_), .Y(w_cout_7_) );
INVX1 INVX1_8 ( .A(skip0_cin_next), .Y(_60_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_61_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_62_) );
NAND3X1 NAND3X1_8 ( .A(_60_), .B(_62_), .C(_61_), .Y(_63_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_57_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_58_) );
OAI21X1 OAI21X1_15 ( .A(_57_), .B(_58_), .C(skip0_cin_next), .Y(_59_) );
NAND2X1 NAND2X1_2 ( .A(_59_), .B(_63_), .Y(_0__4_) );
OAI21X1 OAI21X1_16 ( .A(_60_), .B(_57_), .C(_62_), .Y(_2__1_) );
INVX1 INVX1_9 ( .A(_2__1_), .Y(_67_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_68_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_69_) );
NAND3X1 NAND3X1_9 ( .A(_67_), .B(_69_), .C(_68_), .Y(_70_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_64_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_65_) );
OAI21X1 OAI21X1_17 ( .A(_64_), .B(_65_), .C(_2__1_), .Y(_66_) );
NAND2X1 NAND2X1_4 ( .A(_66_), .B(_70_), .Y(_0__5_) );
OAI21X1 OAI21X1_18 ( .A(_67_), .B(_64_), .C(_69_), .Y(_2__2_) );
INVX1 INVX1_10 ( .A(_2__2_), .Y(_74_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_75_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_76_) );
NAND3X1 NAND3X1_10 ( .A(_74_), .B(_76_), .C(_75_), .Y(_77_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_71_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_72_) );
OAI21X1 OAI21X1_19 ( .A(_71_), .B(_72_), .C(_2__2_), .Y(_73_) );
NAND2X1 NAND2X1_6 ( .A(_73_), .B(_77_), .Y(_0__6_) );
OAI21X1 OAI21X1_20 ( .A(_74_), .B(_71_), .C(_76_), .Y(_2__3_) );
INVX1 INVX1_11 ( .A(_2__3_), .Y(_81_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_82_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_83_) );
NAND3X1 NAND3X1_11 ( .A(_81_), .B(_83_), .C(_82_), .Y(_84_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_78_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_79_) );
OAI21X1 OAI21X1_21 ( .A(_78_), .B(_79_), .C(_2__3_), .Y(_80_) );
NAND2X1 NAND2X1_8 ( .A(_80_), .B(_84_), .Y(_0__7_) );
OAI21X1 OAI21X1_22 ( .A(_81_), .B(_78_), .C(_83_), .Y(_1_) );
INVX1 INVX1_12 ( .A(w_cout_1_), .Y(_88_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_89_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_90_) );
NAND3X1 NAND3X1_12 ( .A(_88_), .B(_90_), .C(_89_), .Y(_91_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_85_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_86_) );
OAI21X1 OAI21X1_23 ( .A(_85_), .B(_86_), .C(w_cout_1_), .Y(_87_) );
NAND2X1 NAND2X1_10 ( .A(_87_), .B(_91_), .Y(_0__8_) );
OAI21X1 OAI21X1_24 ( .A(_88_), .B(_85_), .C(_90_), .Y(_4__1_) );
INVX1 INVX1_13 ( .A(_4__1_), .Y(_95_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_96_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_97_) );
NAND3X1 NAND3X1_13 ( .A(_95_), .B(_97_), .C(_96_), .Y(_98_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_92_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_93_) );
OAI21X1 OAI21X1_25 ( .A(_92_), .B(_93_), .C(_4__1_), .Y(_94_) );
NAND2X1 NAND2X1_12 ( .A(_94_), .B(_98_), .Y(_0__9_) );
OAI21X1 OAI21X1_26 ( .A(_95_), .B(_92_), .C(_97_), .Y(_4__2_) );
INVX1 INVX1_14 ( .A(_4__2_), .Y(_102_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_103_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_104_) );
NAND3X1 NAND3X1_14 ( .A(_102_), .B(_104_), .C(_103_), .Y(_105_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_99_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_100_) );
OAI21X1 OAI21X1_27 ( .A(_99_), .B(_100_), .C(_4__2_), .Y(_101_) );
NAND2X1 NAND2X1_14 ( .A(_101_), .B(_105_), .Y(_0__10_) );
OAI21X1 OAI21X1_28 ( .A(_102_), .B(_99_), .C(_104_), .Y(_4__3_) );
INVX1 INVX1_15 ( .A(_4__3_), .Y(_109_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_110_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_111_) );
NAND3X1 NAND3X1_15 ( .A(_109_), .B(_111_), .C(_110_), .Y(_112_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_106_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_107_) );
OAI21X1 OAI21X1_29 ( .A(_106_), .B(_107_), .C(_4__3_), .Y(_108_) );
NAND2X1 NAND2X1_16 ( .A(_108_), .B(_112_), .Y(_0__11_) );
OAI21X1 OAI21X1_30 ( .A(_109_), .B(_106_), .C(_111_), .Y(_3_) );
INVX1 INVX1_16 ( .A(w_cout_2_), .Y(_116_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_117_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_118_) );
NAND3X1 NAND3X1_16 ( .A(_116_), .B(_118_), .C(_117_), .Y(_119_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_113_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_114_) );
OAI21X1 OAI21X1_31 ( .A(_113_), .B(_114_), .C(w_cout_2_), .Y(_115_) );
NAND2X1 NAND2X1_18 ( .A(_115_), .B(_119_), .Y(_0__12_) );
OAI21X1 OAI21X1_32 ( .A(_116_), .B(_113_), .C(_118_), .Y(_6__1_) );
INVX1 INVX1_17 ( .A(_6__1_), .Y(_123_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_124_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_125_) );
NAND3X1 NAND3X1_17 ( .A(_123_), .B(_125_), .C(_124_), .Y(_126_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_120_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_121_) );
OAI21X1 OAI21X1_33 ( .A(_120_), .B(_121_), .C(_6__1_), .Y(_122_) );
NAND2X1 NAND2X1_20 ( .A(_122_), .B(_126_), .Y(_0__13_) );
OAI21X1 OAI21X1_34 ( .A(_123_), .B(_120_), .C(_125_), .Y(_6__2_) );
INVX1 INVX1_18 ( .A(_6__2_), .Y(_130_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_131_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_132_) );
NAND3X1 NAND3X1_18 ( .A(_130_), .B(_132_), .C(_131_), .Y(_133_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_127_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_128_) );
OAI21X1 OAI21X1_35 ( .A(_127_), .B(_128_), .C(_6__2_), .Y(_129_) );
NAND2X1 NAND2X1_22 ( .A(_129_), .B(_133_), .Y(_0__14_) );
OAI21X1 OAI21X1_36 ( .A(_130_), .B(_127_), .C(_132_), .Y(_6__3_) );
INVX1 INVX1_19 ( .A(_6__3_), .Y(_137_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_138_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_139_) );
NAND3X1 NAND3X1_19 ( .A(_137_), .B(_139_), .C(_138_), .Y(_140_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_134_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_135_) );
OAI21X1 OAI21X1_37 ( .A(_134_), .B(_135_), .C(_6__3_), .Y(_136_) );
NAND2X1 NAND2X1_24 ( .A(_136_), .B(_140_), .Y(_0__15_) );
OAI21X1 OAI21X1_38 ( .A(_137_), .B(_134_), .C(_139_), .Y(_5_) );
INVX1 INVX1_20 ( .A(w_cout_3_), .Y(_144_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_145_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_146_) );
NAND3X1 NAND3X1_20 ( .A(_144_), .B(_146_), .C(_145_), .Y(_147_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_141_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_142_) );
OAI21X1 OAI21X1_39 ( .A(_141_), .B(_142_), .C(w_cout_3_), .Y(_143_) );
NAND2X1 NAND2X1_26 ( .A(_143_), .B(_147_), .Y(_0__16_) );
OAI21X1 OAI21X1_40 ( .A(_144_), .B(_141_), .C(_146_), .Y(_8__1_) );
INVX1 INVX1_21 ( .A(_8__1_), .Y(_151_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_152_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_153_) );
NAND3X1 NAND3X1_21 ( .A(_151_), .B(_153_), .C(_152_), .Y(_154_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_148_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_149_) );
OAI21X1 OAI21X1_41 ( .A(_148_), .B(_149_), .C(_8__1_), .Y(_150_) );
NAND2X1 NAND2X1_28 ( .A(_150_), .B(_154_), .Y(_0__17_) );
OAI21X1 OAI21X1_42 ( .A(_151_), .B(_148_), .C(_153_), .Y(_8__2_) );
INVX1 INVX1_22 ( .A(_8__2_), .Y(_158_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_159_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_160_) );
NAND3X1 NAND3X1_22 ( .A(_158_), .B(_160_), .C(_159_), .Y(_161_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_155_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_156_) );
OAI21X1 OAI21X1_43 ( .A(_155_), .B(_156_), .C(_8__2_), .Y(_157_) );
NAND2X1 NAND2X1_30 ( .A(_157_), .B(_161_), .Y(_0__18_) );
OAI21X1 OAI21X1_44 ( .A(_158_), .B(_155_), .C(_160_), .Y(_8__3_) );
INVX1 INVX1_23 ( .A(_8__3_), .Y(_165_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_166_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_167_) );
NAND3X1 NAND3X1_23 ( .A(_165_), .B(_167_), .C(_166_), .Y(_168_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_162_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_163_) );
OAI21X1 OAI21X1_45 ( .A(_162_), .B(_163_), .C(_8__3_), .Y(_164_) );
NAND2X1 NAND2X1_32 ( .A(_164_), .B(_168_), .Y(_0__19_) );
OAI21X1 OAI21X1_46 ( .A(_165_), .B(_162_), .C(_167_), .Y(_7_) );
INVX1 INVX1_24 ( .A(w_cout_4_), .Y(_172_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_173_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_174_) );
NAND3X1 NAND3X1_24 ( .A(_172_), .B(_174_), .C(_173_), .Y(_175_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_169_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_170_) );
OAI21X1 OAI21X1_47 ( .A(_169_), .B(_170_), .C(w_cout_4_), .Y(_171_) );
NAND2X1 NAND2X1_34 ( .A(_171_), .B(_175_), .Y(_0__20_) );
OAI21X1 OAI21X1_48 ( .A(_172_), .B(_169_), .C(_174_), .Y(_10__1_) );
INVX1 INVX1_25 ( .A(_10__1_), .Y(_179_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_180_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_181_) );
NAND3X1 NAND3X1_25 ( .A(_179_), .B(_181_), .C(_180_), .Y(_182_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_176_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_177_) );
OAI21X1 OAI21X1_49 ( .A(_176_), .B(_177_), .C(_10__1_), .Y(_178_) );
NAND2X1 NAND2X1_36 ( .A(_178_), .B(_182_), .Y(_0__21_) );
OAI21X1 OAI21X1_50 ( .A(_179_), .B(_176_), .C(_181_), .Y(_10__2_) );
INVX1 INVX1_26 ( .A(_10__2_), .Y(_186_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_187_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_188_) );
NAND3X1 NAND3X1_26 ( .A(_186_), .B(_188_), .C(_187_), .Y(_189_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_183_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_184_) );
OAI21X1 OAI21X1_51 ( .A(_183_), .B(_184_), .C(_10__2_), .Y(_185_) );
NAND2X1 NAND2X1_38 ( .A(_185_), .B(_189_), .Y(_0__22_) );
OAI21X1 OAI21X1_52 ( .A(_186_), .B(_183_), .C(_188_), .Y(_10__3_) );
INVX1 INVX1_27 ( .A(_10__3_), .Y(_193_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_194_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_195_) );
NAND3X1 NAND3X1_27 ( .A(_193_), .B(_195_), .C(_194_), .Y(_196_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_190_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_191_) );
OAI21X1 OAI21X1_53 ( .A(_190_), .B(_191_), .C(_10__3_), .Y(_192_) );
NAND2X1 NAND2X1_40 ( .A(_192_), .B(_196_), .Y(_0__23_) );
OAI21X1 OAI21X1_54 ( .A(_193_), .B(_190_), .C(_195_), .Y(_9_) );
INVX1 INVX1_28 ( .A(w_cout_5_), .Y(_200_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_201_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_202_) );
NAND3X1 NAND3X1_28 ( .A(_200_), .B(_202_), .C(_201_), .Y(_203_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_197_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_198_) );
OAI21X1 OAI21X1_55 ( .A(_197_), .B(_198_), .C(w_cout_5_), .Y(_199_) );
NAND2X1 NAND2X1_42 ( .A(_199_), .B(_203_), .Y(_0__24_) );
OAI21X1 OAI21X1_56 ( .A(_200_), .B(_197_), .C(_202_), .Y(_12__1_) );
INVX1 INVX1_29 ( .A(_12__1_), .Y(_207_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_208_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_209_) );
NAND3X1 NAND3X1_29 ( .A(_207_), .B(_209_), .C(_208_), .Y(_210_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_204_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_205_) );
OAI21X1 OAI21X1_57 ( .A(_204_), .B(_205_), .C(_12__1_), .Y(_206_) );
NAND2X1 NAND2X1_44 ( .A(_206_), .B(_210_), .Y(_0__25_) );
OAI21X1 OAI21X1_58 ( .A(_207_), .B(_204_), .C(_209_), .Y(_12__2_) );
INVX1 INVX1_30 ( .A(_12__2_), .Y(_214_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_215_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_216_) );
NAND3X1 NAND3X1_30 ( .A(_214_), .B(_216_), .C(_215_), .Y(_217_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_211_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_212_) );
OAI21X1 OAI21X1_59 ( .A(_211_), .B(_212_), .C(_12__2_), .Y(_213_) );
NAND2X1 NAND2X1_46 ( .A(_213_), .B(_217_), .Y(_0__26_) );
OAI21X1 OAI21X1_60 ( .A(_214_), .B(_211_), .C(_216_), .Y(_12__3_) );
INVX1 INVX1_31 ( .A(_12__3_), .Y(_221_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_222_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_223_) );
NAND3X1 NAND3X1_31 ( .A(_221_), .B(_223_), .C(_222_), .Y(_224_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_218_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_219_) );
OAI21X1 OAI21X1_61 ( .A(_218_), .B(_219_), .C(_12__3_), .Y(_220_) );
NAND2X1 NAND2X1_48 ( .A(_220_), .B(_224_), .Y(_0__27_) );
OAI21X1 OAI21X1_62 ( .A(_221_), .B(_218_), .C(_223_), .Y(_11_) );
INVX1 INVX1_32 ( .A(w_cout_6_), .Y(_228_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_229_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_230_) );
NAND3X1 NAND3X1_32 ( .A(_228_), .B(_230_), .C(_229_), .Y(_231_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_225_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_226_) );
OAI21X1 OAI21X1_63 ( .A(_225_), .B(_226_), .C(w_cout_6_), .Y(_227_) );
NAND2X1 NAND2X1_50 ( .A(_227_), .B(_231_), .Y(_0__28_) );
OAI21X1 OAI21X1_64 ( .A(_228_), .B(_225_), .C(_230_), .Y(_14__1_) );
INVX1 INVX1_33 ( .A(_14__1_), .Y(_235_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_236_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_237_) );
NAND3X1 NAND3X1_33 ( .A(_235_), .B(_237_), .C(_236_), .Y(_238_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_232_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_233_) );
OAI21X1 OAI21X1_65 ( .A(_232_), .B(_233_), .C(_14__1_), .Y(_234_) );
NAND2X1 NAND2X1_52 ( .A(_234_), .B(_238_), .Y(_0__29_) );
OAI21X1 OAI21X1_66 ( .A(_235_), .B(_232_), .C(_237_), .Y(_14__2_) );
INVX1 INVX1_34 ( .A(_14__2_), .Y(_242_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_243_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_244_) );
NAND3X1 NAND3X1_34 ( .A(_242_), .B(_244_), .C(_243_), .Y(_245_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_239_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_240_) );
OAI21X1 OAI21X1_67 ( .A(_239_), .B(_240_), .C(_14__2_), .Y(_241_) );
NAND2X1 NAND2X1_54 ( .A(_241_), .B(_245_), .Y(_0__30_) );
OAI21X1 OAI21X1_68 ( .A(_242_), .B(_239_), .C(_244_), .Y(_14__3_) );
INVX1 INVX1_35 ( .A(_14__3_), .Y(_249_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_250_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_251_) );
NAND3X1 NAND3X1_35 ( .A(_249_), .B(_251_), .C(_250_), .Y(_252_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_246_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_247_) );
OAI21X1 OAI21X1_69 ( .A(_246_), .B(_247_), .C(_14__3_), .Y(_248_) );
NAND2X1 NAND2X1_56 ( .A(_248_), .B(_252_), .Y(_0__31_) );
OAI21X1 OAI21X1_70 ( .A(_249_), .B(_246_), .C(_251_), .Y(_13_) );
INVX1 INVX1_36 ( .A(1'b0), .Y(_256_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_257_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_258_) );
NAND3X1 NAND3X1_36 ( .A(_256_), .B(_258_), .C(_257_), .Y(_259_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_253_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_254_) );
OAI21X1 OAI21X1_71 ( .A(_253_), .B(_254_), .C(1'b0), .Y(_255_) );
NAND2X1 NAND2X1_58 ( .A(_255_), .B(_259_), .Y(_0__0_) );
OAI21X1 OAI21X1_72 ( .A(_256_), .B(_253_), .C(_258_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_37 ( .A(rca_inst_w_CARRY_1_), .Y(_263_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_264_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_265_) );
NAND3X1 NAND3X1_37 ( .A(_263_), .B(_265_), .C(_264_), .Y(_266_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_260_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_261_) );
OAI21X1 OAI21X1_73 ( .A(_260_), .B(_261_), .C(rca_inst_w_CARRY_1_), .Y(_262_) );
NAND2X1 NAND2X1_60 ( .A(_262_), .B(_266_), .Y(_0__1_) );
OAI21X1 OAI21X1_74 ( .A(_263_), .B(_260_), .C(_265_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_38 ( .A(rca_inst_w_CARRY_2_), .Y(_270_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_271_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_272_) );
NAND3X1 NAND3X1_38 ( .A(_270_), .B(_272_), .C(_271_), .Y(_273_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_267_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_268_) );
OAI21X1 OAI21X1_75 ( .A(_267_), .B(_268_), .C(rca_inst_w_CARRY_2_), .Y(_269_) );
NAND2X1 NAND2X1_62 ( .A(_269_), .B(_273_), .Y(_0__2_) );
OAI21X1 OAI21X1_76 ( .A(_270_), .B(_267_), .C(_272_), .Y(rca_inst_w_CARRY_3_) );
INVX1 INVX1_39 ( .A(rca_inst_w_CARRY_3_), .Y(_277_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_278_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_279_) );
NAND3X1 NAND3X1_39 ( .A(_277_), .B(_279_), .C(_278_), .Y(_280_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_274_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_275_) );
OAI21X1 OAI21X1_77 ( .A(_274_), .B(_275_), .C(rca_inst_w_CARRY_3_), .Y(_276_) );
NAND2X1 NAND2X1_64 ( .A(_276_), .B(_280_), .Y(_0__3_) );
OAI21X1 OAI21X1_78 ( .A(_277_), .B(_274_), .C(_279_), .Y(cout0) );
INVX1 INVX1_40 ( .A(cout0), .Y(_281_) );
OAI21X1 OAI21X1_79 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .C(1'b0), .Y(_282_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_283_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_284_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_285_) );
NAND3X1 NAND3X1_40 ( .A(_283_), .B(_284_), .C(_285_), .Y(_286_) );
OAI21X1 OAI21X1_80 ( .A(_282_), .B(_286_), .C(_281_), .Y(skip0_cin_next) );
BUFX2 BUFX2_34 ( .A(skip0_cin_next), .Y(_2__0_) );
BUFX2 BUFX2_35 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_36 ( .A(w_cout_1_), .Y(_4__0_) );
BUFX2 BUFX2_37 ( .A(_3_), .Y(_4__4_) );
BUFX2 BUFX2_38 ( .A(w_cout_2_), .Y(_6__0_) );
BUFX2 BUFX2_39 ( .A(_5_), .Y(_6__4_) );
BUFX2 BUFX2_40 ( .A(w_cout_3_), .Y(_8__0_) );
BUFX2 BUFX2_41 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_42 ( .A(w_cout_4_), .Y(_10__0_) );
BUFX2 BUFX2_43 ( .A(_9_), .Y(_10__4_) );
BUFX2 BUFX2_44 ( .A(w_cout_5_), .Y(_12__0_) );
BUFX2 BUFX2_45 ( .A(_11_), .Y(_12__4_) );
BUFX2 BUFX2_46 ( .A(w_cout_6_), .Y(_14__0_) );
BUFX2 BUFX2_47 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_48 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_49 ( .A(cout0), .Y(rca_inst_w_CARRY_4_) );
BUFX2 BUFX2_50 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
