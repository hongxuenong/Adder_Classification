module CSkipA_64bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term1[45], i_add_term1[46], i_add_term1[47], i_add_term1[48], i_add_term1[49], i_add_term1[50], i_add_term1[51], i_add_term1[52], i_add_term1[53], i_add_term1[54], i_add_term1[55], i_add_term1[56], i_add_term1[57], i_add_term1[58], i_add_term1[59], i_add_term1[60], i_add_term1[61], i_add_term1[62], i_add_term1[63], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], i_add_term2[45], i_add_term2[46], i_add_term2[47], i_add_term2[48], i_add_term2[49], i_add_term2[50], i_add_term2[51], i_add_term2[52], i_add_term2[53], i_add_term2[54], i_add_term2[55], i_add_term2[56], i_add_term2[57], i_add_term2[58], i_add_term2[59], i_add_term2[60], i_add_term2[61], i_add_term2[62], i_add_term2[63], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], sum[45], sum[46], sum[47], sum[48], sum[49], sum[50], sum[51], sum[52], sum[53], sum[54], sum[55], sum[56], sum[57], sum[58], sum[59], sum[60], sum[61], sum[62], sum[63], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term1[45];
input i_add_term1[46];
input i_add_term1[47];
input i_add_term1[48];
input i_add_term1[49];
input i_add_term1[50];
input i_add_term1[51];
input i_add_term1[52];
input i_add_term1[53];
input i_add_term1[54];
input i_add_term1[55];
input i_add_term1[56];
input i_add_term1[57];
input i_add_term1[58];
input i_add_term1[59];
input i_add_term1[60];
input i_add_term1[61];
input i_add_term1[62];
input i_add_term1[63];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
input i_add_term2[45];
input i_add_term2[46];
input i_add_term2[47];
input i_add_term2[48];
input i_add_term2[49];
input i_add_term2[50];
input i_add_term2[51];
input i_add_term2[52];
input i_add_term2[53];
input i_add_term2[54];
input i_add_term2[55];
input i_add_term2[56];
input i_add_term2[57];
input i_add_term2[58];
input i_add_term2[59];
input i_add_term2[60];
input i_add_term2[61];
input i_add_term2[62];
input i_add_term2[63];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output sum[45];
output sum[46];
output sum[47];
output sum[48];
output sum[49];
output sum[50];
output sum[51];
output sum[52];
output sum[53];
output sum[54];
output sum[55];
output sum[56];
output sum[57];
output sum[58];
output sum[59];
output sum[60];
output sum[61];
output sum[62];
output sum[63];
output cout;

NAND3X1 NAND3X1_1 ( .A(_196_), .B(_197_), .C(_192_), .Y(_193_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_194_) );
OAI21X1 OAI21X1_1 ( .A(_198_), .B(_194_), .C(_11__1_), .Y(_195_) );
NAND2X1 NAND2X1_1 ( .A(_195_), .B(_193_), .Y(_0__17_) );
INVX1 INVX1_1 ( .A(_11__2_), .Y(_203_) );
NAND2X1 NAND2X1_2 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_204_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_205_) );
OAI21X1 OAI21X1_2 ( .A(_203_), .B(_205_), .C(_204_), .Y(_11__3_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_199_) );
NAND3X1 NAND3X1_2 ( .A(_203_), .B(_204_), .C(_199_), .Y(_200_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_201_) );
OAI21X1 OAI21X1_3 ( .A(_205_), .B(_201_), .C(_11__2_), .Y(_202_) );
NAND2X1 NAND2X1_3 ( .A(_202_), .B(_200_), .Y(_0__18_) );
INVX1 INVX1_2 ( .A(i_add_term1[16]), .Y(_206_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[16]), .B(_206_), .Y(_207_) );
INVX1 INVX1_3 ( .A(i_add_term2[16]), .Y(_208_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term1[16]), .B(_208_), .Y(_209_) );
INVX1 INVX1_4 ( .A(i_add_term1[17]), .Y(_210_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[17]), .B(_210_), .Y(_211_) );
INVX1 INVX1_5 ( .A(i_add_term2[17]), .Y(_212_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term1[17]), .B(_212_), .Y(_213_) );
OAI22X1 OAI22X1_1 ( .A(_207_), .B(_209_), .C(_211_), .D(_213_), .Y(_214_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_215_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_216_) );
NOR2X1 NOR2X1_7 ( .A(_215_), .B(_216_), .Y(_217_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_218_) );
NAND2X1 NAND2X1_4 ( .A(_217_), .B(_218_), .Y(_219_) );
NOR2X1 NOR2X1_8 ( .A(_214_), .B(_219_), .Y(_12_) );
INVX1 INVX1_6 ( .A(_10_), .Y(_220_) );
NAND2X1 NAND2X1_5 ( .A(1'b0), .B(_12_), .Y(_221_) );
OAI21X1 OAI21X1_4 ( .A(_12_), .B(_220_), .C(_221_), .Y(w_cout_4_) );
INVX1 INVX1_7 ( .A(w_cout_4_), .Y(_226_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_227_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_228_) );
OAI21X1 OAI21X1_5 ( .A(_226_), .B(_228_), .C(_227_), .Y(_14__1_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_222_) );
NAND3X1 NAND3X1_3 ( .A(_226_), .B(_227_), .C(_222_), .Y(_223_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_224_) );
OAI21X1 OAI21X1_6 ( .A(_228_), .B(_224_), .C(w_cout_4_), .Y(_225_) );
NAND2X1 NAND2X1_7 ( .A(_225_), .B(_223_), .Y(_0__20_) );
INVX1 INVX1_8 ( .A(_14__3_), .Y(_233_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_234_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_235_) );
OAI21X1 OAI21X1_7 ( .A(_233_), .B(_235_), .C(_234_), .Y(_13_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_229_) );
NAND3X1 NAND3X1_4 ( .A(_233_), .B(_234_), .C(_229_), .Y(_230_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_231_) );
OAI21X1 OAI21X1_8 ( .A(_235_), .B(_231_), .C(_14__3_), .Y(_232_) );
NAND2X1 NAND2X1_9 ( .A(_232_), .B(_230_), .Y(_0__23_) );
INVX1 INVX1_9 ( .A(_14__1_), .Y(_240_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_241_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_242_) );
OAI21X1 OAI21X1_9 ( .A(_240_), .B(_242_), .C(_241_), .Y(_14__2_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_236_) );
NAND3X1 NAND3X1_5 ( .A(_240_), .B(_241_), .C(_236_), .Y(_237_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_238_) );
OAI21X1 OAI21X1_10 ( .A(_242_), .B(_238_), .C(_14__1_), .Y(_239_) );
NAND2X1 NAND2X1_11 ( .A(_239_), .B(_237_), .Y(_0__21_) );
INVX1 INVX1_10 ( .A(_14__2_), .Y(_247_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_248_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_249_) );
OAI21X1 OAI21X1_11 ( .A(_247_), .B(_249_), .C(_248_), .Y(_14__3_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_243_) );
NAND3X1 NAND3X1_6 ( .A(_247_), .B(_248_), .C(_243_), .Y(_244_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_245_) );
OAI21X1 OAI21X1_12 ( .A(_249_), .B(_245_), .C(_14__2_), .Y(_246_) );
NAND2X1 NAND2X1_13 ( .A(_246_), .B(_244_), .Y(_0__22_) );
INVX1 INVX1_11 ( .A(i_add_term1[20]), .Y(_250_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[20]), .B(_250_), .Y(_251_) );
INVX1 INVX1_12 ( .A(i_add_term2[20]), .Y(_252_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term1[20]), .B(_252_), .Y(_253_) );
INVX1 INVX1_13 ( .A(i_add_term1[21]), .Y(_254_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[21]), .B(_254_), .Y(_255_) );
INVX1 INVX1_14 ( .A(i_add_term2[21]), .Y(_256_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term1[21]), .B(_256_), .Y(_257_) );
OAI22X1 OAI22X1_2 ( .A(_251_), .B(_253_), .C(_255_), .D(_257_), .Y(_258_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_259_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_260_) );
NOR2X1 NOR2X1_18 ( .A(_259_), .B(_260_), .Y(_261_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_262_) );
NAND2X1 NAND2X1_14 ( .A(_261_), .B(_262_), .Y(_263_) );
NOR2X1 NOR2X1_19 ( .A(_258_), .B(_263_), .Y(_15_) );
INVX1 INVX1_15 ( .A(_13_), .Y(_264_) );
NAND2X1 NAND2X1_15 ( .A(1'b0), .B(_15_), .Y(_265_) );
OAI21X1 OAI21X1_13 ( .A(_15_), .B(_264_), .C(_265_), .Y(w_cout_5_) );
INVX1 INVX1_16 ( .A(w_cout_5_), .Y(_270_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_271_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_272_) );
OAI21X1 OAI21X1_14 ( .A(_270_), .B(_272_), .C(_271_), .Y(_17__1_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_266_) );
NAND3X1 NAND3X1_7 ( .A(_270_), .B(_271_), .C(_266_), .Y(_267_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_268_) );
OAI21X1 OAI21X1_15 ( .A(_272_), .B(_268_), .C(w_cout_5_), .Y(_269_) );
NAND2X1 NAND2X1_17 ( .A(_269_), .B(_267_), .Y(_0__24_) );
INVX1 INVX1_17 ( .A(_17__3_), .Y(_277_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_278_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_279_) );
OAI21X1 OAI21X1_16 ( .A(_277_), .B(_279_), .C(_278_), .Y(_16_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_273_) );
NAND3X1 NAND3X1_8 ( .A(_277_), .B(_278_), .C(_273_), .Y(_274_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_275_) );
OAI21X1 OAI21X1_17 ( .A(_279_), .B(_275_), .C(_17__3_), .Y(_276_) );
NAND2X1 NAND2X1_19 ( .A(_276_), .B(_274_), .Y(_0__27_) );
INVX1 INVX1_18 ( .A(_17__1_), .Y(_284_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_285_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_286_) );
OAI21X1 OAI21X1_18 ( .A(_284_), .B(_286_), .C(_285_), .Y(_17__2_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_280_) );
NAND3X1 NAND3X1_9 ( .A(_284_), .B(_285_), .C(_280_), .Y(_281_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_282_) );
OAI21X1 OAI21X1_19 ( .A(_286_), .B(_282_), .C(_17__1_), .Y(_283_) );
NAND2X1 NAND2X1_21 ( .A(_283_), .B(_281_), .Y(_0__25_) );
INVX1 INVX1_19 ( .A(_17__2_), .Y(_291_) );
NAND2X1 NAND2X1_22 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_292_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_293_) );
OAI21X1 OAI21X1_20 ( .A(_291_), .B(_293_), .C(_292_), .Y(_17__3_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_287_) );
NAND3X1 NAND3X1_10 ( .A(_291_), .B(_292_), .C(_287_), .Y(_288_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_289_) );
OAI21X1 OAI21X1_21 ( .A(_293_), .B(_289_), .C(_17__2_), .Y(_290_) );
NAND2X1 NAND2X1_23 ( .A(_290_), .B(_288_), .Y(_0__26_) );
INVX1 INVX1_20 ( .A(i_add_term1[24]), .Y(_294_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[24]), .B(_294_), .Y(_295_) );
INVX1 INVX1_21 ( .A(i_add_term2[24]), .Y(_296_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term1[24]), .B(_296_), .Y(_297_) );
INVX1 INVX1_22 ( .A(i_add_term1[25]), .Y(_298_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[25]), .B(_298_), .Y(_299_) );
INVX1 INVX1_23 ( .A(i_add_term2[25]), .Y(_300_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term1[25]), .B(_300_), .Y(_301_) );
OAI22X1 OAI22X1_3 ( .A(_295_), .B(_297_), .C(_299_), .D(_301_), .Y(_302_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_303_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_304_) );
NOR2X1 NOR2X1_29 ( .A(_303_), .B(_304_), .Y(_305_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_306_) );
NAND2X1 NAND2X1_24 ( .A(_305_), .B(_306_), .Y(_307_) );
NOR2X1 NOR2X1_30 ( .A(_302_), .B(_307_), .Y(_18_) );
INVX1 INVX1_24 ( .A(_16_), .Y(_308_) );
NAND2X1 NAND2X1_25 ( .A(1'b0), .B(_18_), .Y(_309_) );
OAI21X1 OAI21X1_22 ( .A(_18_), .B(_308_), .C(_309_), .Y(w_cout_6_) );
INVX1 INVX1_25 ( .A(w_cout_6_), .Y(_314_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_315_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_316_) );
OAI21X1 OAI21X1_23 ( .A(_314_), .B(_316_), .C(_315_), .Y(_20__1_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_310_) );
NAND3X1 NAND3X1_11 ( .A(_314_), .B(_315_), .C(_310_), .Y(_311_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_312_) );
OAI21X1 OAI21X1_24 ( .A(_316_), .B(_312_), .C(w_cout_6_), .Y(_313_) );
NAND2X1 NAND2X1_27 ( .A(_313_), .B(_311_), .Y(_0__28_) );
INVX1 INVX1_26 ( .A(_20__3_), .Y(_321_) );
NAND2X1 NAND2X1_28 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_322_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_323_) );
OAI21X1 OAI21X1_25 ( .A(_321_), .B(_323_), .C(_322_), .Y(_19_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_317_) );
NAND3X1 NAND3X1_12 ( .A(_321_), .B(_322_), .C(_317_), .Y(_318_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_319_) );
OAI21X1 OAI21X1_26 ( .A(_323_), .B(_319_), .C(_20__3_), .Y(_320_) );
NAND2X1 NAND2X1_29 ( .A(_320_), .B(_318_), .Y(_0__31_) );
INVX1 INVX1_27 ( .A(_20__1_), .Y(_328_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_329_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_330_) );
OAI21X1 OAI21X1_27 ( .A(_328_), .B(_330_), .C(_329_), .Y(_20__2_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_324_) );
NAND3X1 NAND3X1_13 ( .A(_328_), .B(_329_), .C(_324_), .Y(_325_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_326_) );
OAI21X1 OAI21X1_28 ( .A(_330_), .B(_326_), .C(_20__1_), .Y(_327_) );
NAND2X1 NAND2X1_31 ( .A(_327_), .B(_325_), .Y(_0__29_) );
INVX1 INVX1_28 ( .A(_20__2_), .Y(_335_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_336_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_337_) );
OAI21X1 OAI21X1_29 ( .A(_335_), .B(_337_), .C(_336_), .Y(_20__3_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_331_) );
NAND3X1 NAND3X1_14 ( .A(_335_), .B(_336_), .C(_331_), .Y(_332_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_333_) );
OAI21X1 OAI21X1_30 ( .A(_337_), .B(_333_), .C(_20__2_), .Y(_334_) );
NAND2X1 NAND2X1_33 ( .A(_334_), .B(_332_), .Y(_0__30_) );
INVX1 INVX1_29 ( .A(i_add_term1[28]), .Y(_338_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[28]), .B(_338_), .Y(_339_) );
INVX1 INVX1_30 ( .A(i_add_term2[28]), .Y(_340_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term1[28]), .B(_340_), .Y(_341_) );
INVX1 INVX1_31 ( .A(i_add_term1[29]), .Y(_342_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[29]), .B(_342_), .Y(_343_) );
INVX1 INVX1_32 ( .A(i_add_term2[29]), .Y(_344_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term1[29]), .B(_344_), .Y(_345_) );
OAI22X1 OAI22X1_4 ( .A(_339_), .B(_341_), .C(_343_), .D(_345_), .Y(_346_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_347_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_348_) );
NOR2X1 NOR2X1_40 ( .A(_347_), .B(_348_), .Y(_349_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_350_) );
NAND2X1 NAND2X1_34 ( .A(_349_), .B(_350_), .Y(_351_) );
NOR2X1 NOR2X1_41 ( .A(_346_), .B(_351_), .Y(_21_) );
INVX1 INVX1_33 ( .A(_19_), .Y(_352_) );
NAND2X1 NAND2X1_35 ( .A(1'b0), .B(_21_), .Y(_353_) );
OAI21X1 OAI21X1_31 ( .A(_21_), .B(_352_), .C(_353_), .Y(w_cout_7_) );
INVX1 INVX1_34 ( .A(w_cout_7_), .Y(_358_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_359_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_360_) );
OAI21X1 OAI21X1_32 ( .A(_358_), .B(_360_), .C(_359_), .Y(_23__1_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_354_) );
NAND3X1 NAND3X1_15 ( .A(_358_), .B(_359_), .C(_354_), .Y(_355_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_356_) );
OAI21X1 OAI21X1_33 ( .A(_360_), .B(_356_), .C(w_cout_7_), .Y(_357_) );
NAND2X1 NAND2X1_37 ( .A(_357_), .B(_355_), .Y(_0__32_) );
INVX1 INVX1_35 ( .A(_23__3_), .Y(_365_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_366_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_367_) );
OAI21X1 OAI21X1_34 ( .A(_365_), .B(_367_), .C(_366_), .Y(_22_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_361_) );
NAND3X1 NAND3X1_16 ( .A(_365_), .B(_366_), .C(_361_), .Y(_362_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_363_) );
OAI21X1 OAI21X1_35 ( .A(_367_), .B(_363_), .C(_23__3_), .Y(_364_) );
NAND2X1 NAND2X1_39 ( .A(_364_), .B(_362_), .Y(_0__35_) );
INVX1 INVX1_36 ( .A(_23__1_), .Y(_372_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_373_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_374_) );
OAI21X1 OAI21X1_36 ( .A(_372_), .B(_374_), .C(_373_), .Y(_23__2_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_368_) );
NAND3X1 NAND3X1_17 ( .A(_372_), .B(_373_), .C(_368_), .Y(_369_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_370_) );
OAI21X1 OAI21X1_37 ( .A(_374_), .B(_370_), .C(_23__1_), .Y(_371_) );
NAND2X1 NAND2X1_41 ( .A(_371_), .B(_369_), .Y(_0__33_) );
INVX1 INVX1_37 ( .A(_23__2_), .Y(_379_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_380_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_381_) );
OAI21X1 OAI21X1_38 ( .A(_379_), .B(_381_), .C(_380_), .Y(_23__3_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_375_) );
NAND3X1 NAND3X1_18 ( .A(_379_), .B(_380_), .C(_375_), .Y(_376_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_377_) );
OAI21X1 OAI21X1_39 ( .A(_381_), .B(_377_), .C(_23__2_), .Y(_378_) );
NAND2X1 NAND2X1_43 ( .A(_378_), .B(_376_), .Y(_0__34_) );
INVX1 INVX1_38 ( .A(i_add_term1[32]), .Y(_382_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[32]), .B(_382_), .Y(_383_) );
INVX1 INVX1_39 ( .A(i_add_term2[32]), .Y(_384_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term1[32]), .B(_384_), .Y(_385_) );
INVX1 INVX1_40 ( .A(i_add_term1[33]), .Y(_386_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[33]), .B(_386_), .Y(_387_) );
INVX1 INVX1_41 ( .A(i_add_term2[33]), .Y(_388_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term1[33]), .B(_388_), .Y(_389_) );
OAI22X1 OAI22X1_5 ( .A(_383_), .B(_385_), .C(_387_), .D(_389_), .Y(_390_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_391_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_392_) );
NOR2X1 NOR2X1_51 ( .A(_391_), .B(_392_), .Y(_393_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_394_) );
NAND2X1 NAND2X1_44 ( .A(_393_), .B(_394_), .Y(_395_) );
NOR2X1 NOR2X1_52 ( .A(_390_), .B(_395_), .Y(_24_) );
INVX1 INVX1_42 ( .A(_22_), .Y(_396_) );
NAND2X1 NAND2X1_45 ( .A(1'b0), .B(_24_), .Y(_397_) );
OAI21X1 OAI21X1_40 ( .A(_24_), .B(_396_), .C(_397_), .Y(w_cout_8_) );
INVX1 INVX1_43 ( .A(w_cout_8_), .Y(_402_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_403_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_404_) );
OAI21X1 OAI21X1_41 ( .A(_402_), .B(_404_), .C(_403_), .Y(_26__1_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_398_) );
NAND3X1 NAND3X1_19 ( .A(_402_), .B(_403_), .C(_398_), .Y(_399_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_400_) );
OAI21X1 OAI21X1_42 ( .A(_404_), .B(_400_), .C(w_cout_8_), .Y(_401_) );
NAND2X1 NAND2X1_47 ( .A(_401_), .B(_399_), .Y(_0__36_) );
INVX1 INVX1_44 ( .A(_26__3_), .Y(_409_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_410_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_411_) );
OAI21X1 OAI21X1_43 ( .A(_409_), .B(_411_), .C(_410_), .Y(_25_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_405_) );
NAND3X1 NAND3X1_20 ( .A(_409_), .B(_410_), .C(_405_), .Y(_406_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_407_) );
OAI21X1 OAI21X1_44 ( .A(_411_), .B(_407_), .C(_26__3_), .Y(_408_) );
NAND2X1 NAND2X1_49 ( .A(_408_), .B(_406_), .Y(_0__39_) );
INVX1 INVX1_45 ( .A(_26__1_), .Y(_416_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_417_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_418_) );
OAI21X1 OAI21X1_45 ( .A(_416_), .B(_418_), .C(_417_), .Y(_26__2_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_412_) );
NAND3X1 NAND3X1_21 ( .A(_416_), .B(_417_), .C(_412_), .Y(_413_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_414_) );
OAI21X1 OAI21X1_46 ( .A(_418_), .B(_414_), .C(_26__1_), .Y(_415_) );
NAND2X1 NAND2X1_51 ( .A(_415_), .B(_413_), .Y(_0__37_) );
INVX1 INVX1_46 ( .A(_26__2_), .Y(_423_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_424_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_425_) );
OAI21X1 OAI21X1_47 ( .A(_423_), .B(_425_), .C(_424_), .Y(_26__3_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_419_) );
NAND3X1 NAND3X1_22 ( .A(_423_), .B(_424_), .C(_419_), .Y(_420_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_421_) );
OAI21X1 OAI21X1_48 ( .A(_425_), .B(_421_), .C(_26__2_), .Y(_422_) );
NAND2X1 NAND2X1_53 ( .A(_422_), .B(_420_), .Y(_0__38_) );
INVX1 INVX1_47 ( .A(i_add_term1[36]), .Y(_426_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[36]), .B(_426_), .Y(_427_) );
INVX1 INVX1_48 ( .A(i_add_term2[36]), .Y(_428_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term1[36]), .B(_428_), .Y(_429_) );
INVX1 INVX1_49 ( .A(i_add_term1[37]), .Y(_430_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[37]), .B(_430_), .Y(_431_) );
INVX1 INVX1_50 ( .A(i_add_term2[37]), .Y(_432_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term1[37]), .B(_432_), .Y(_433_) );
OAI22X1 OAI22X1_6 ( .A(_427_), .B(_429_), .C(_431_), .D(_433_), .Y(_434_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_435_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_436_) );
NOR2X1 NOR2X1_62 ( .A(_435_), .B(_436_), .Y(_437_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_438_) );
NAND2X1 NAND2X1_54 ( .A(_437_), .B(_438_), .Y(_439_) );
NOR2X1 NOR2X1_63 ( .A(_434_), .B(_439_), .Y(_27_) );
INVX1 INVX1_51 ( .A(_25_), .Y(_440_) );
NAND2X1 NAND2X1_55 ( .A(1'b0), .B(_27_), .Y(_441_) );
OAI21X1 OAI21X1_49 ( .A(_27_), .B(_440_), .C(_441_), .Y(w_cout_9_) );
INVX1 INVX1_52 ( .A(w_cout_9_), .Y(_446_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_447_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_448_) );
OAI21X1 OAI21X1_50 ( .A(_446_), .B(_448_), .C(_447_), .Y(_29__1_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_442_) );
NAND3X1 NAND3X1_23 ( .A(_446_), .B(_447_), .C(_442_), .Y(_443_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_444_) );
OAI21X1 OAI21X1_51 ( .A(_448_), .B(_444_), .C(w_cout_9_), .Y(_445_) );
NAND2X1 NAND2X1_57 ( .A(_445_), .B(_443_), .Y(_0__40_) );
INVX1 INVX1_53 ( .A(_29__3_), .Y(_453_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_454_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_455_) );
OAI21X1 OAI21X1_52 ( .A(_453_), .B(_455_), .C(_454_), .Y(_28_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_449_) );
NAND3X1 NAND3X1_24 ( .A(_453_), .B(_454_), .C(_449_), .Y(_450_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_451_) );
OAI21X1 OAI21X1_53 ( .A(_455_), .B(_451_), .C(_29__3_), .Y(_452_) );
NAND2X1 NAND2X1_59 ( .A(_452_), .B(_450_), .Y(_0__43_) );
INVX1 INVX1_54 ( .A(_29__1_), .Y(_460_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_461_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_462_) );
OAI21X1 OAI21X1_54 ( .A(_460_), .B(_462_), .C(_461_), .Y(_29__2_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_456_) );
NAND3X1 NAND3X1_25 ( .A(_460_), .B(_461_), .C(_456_), .Y(_457_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_458_) );
OAI21X1 OAI21X1_55 ( .A(_462_), .B(_458_), .C(_29__1_), .Y(_459_) );
NAND2X1 NAND2X1_61 ( .A(_459_), .B(_457_), .Y(_0__41_) );
INVX1 INVX1_55 ( .A(_29__2_), .Y(_467_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_468_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_469_) );
OAI21X1 OAI21X1_56 ( .A(_467_), .B(_469_), .C(_468_), .Y(_29__3_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_463_) );
NAND3X1 NAND3X1_26 ( .A(_467_), .B(_468_), .C(_463_), .Y(_464_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_465_) );
OAI21X1 OAI21X1_57 ( .A(_469_), .B(_465_), .C(_29__2_), .Y(_466_) );
NAND2X1 NAND2X1_63 ( .A(_466_), .B(_464_), .Y(_0__42_) );
INVX1 INVX1_56 ( .A(i_add_term1[40]), .Y(_470_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[40]), .B(_470_), .Y(_471_) );
INVX1 INVX1_57 ( .A(i_add_term2[40]), .Y(_472_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term1[40]), .B(_472_), .Y(_473_) );
INVX1 INVX1_58 ( .A(i_add_term1[41]), .Y(_474_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[41]), .B(_474_), .Y(_475_) );
INVX1 INVX1_59 ( .A(i_add_term2[41]), .Y(_476_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term1[41]), .B(_476_), .Y(_477_) );
OAI22X1 OAI22X1_7 ( .A(_471_), .B(_473_), .C(_475_), .D(_477_), .Y(_478_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_479_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_480_) );
NOR2X1 NOR2X1_73 ( .A(_479_), .B(_480_), .Y(_481_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_482_) );
NAND2X1 NAND2X1_64 ( .A(_481_), .B(_482_), .Y(_483_) );
NOR2X1 NOR2X1_74 ( .A(_478_), .B(_483_), .Y(_30_) );
INVX1 INVX1_60 ( .A(_28_), .Y(_484_) );
NAND2X1 NAND2X1_65 ( .A(1'b0), .B(_30_), .Y(_485_) );
OAI21X1 OAI21X1_58 ( .A(_30_), .B(_484_), .C(_485_), .Y(w_cout_10_) );
INVX1 INVX1_61 ( .A(w_cout_10_), .Y(_490_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_491_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_492_) );
OAI21X1 OAI21X1_59 ( .A(_490_), .B(_492_), .C(_491_), .Y(_32__1_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_486_) );
NAND3X1 NAND3X1_27 ( .A(_490_), .B(_491_), .C(_486_), .Y(_487_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_488_) );
OAI21X1 OAI21X1_60 ( .A(_492_), .B(_488_), .C(w_cout_10_), .Y(_489_) );
NAND2X1 NAND2X1_67 ( .A(_489_), .B(_487_), .Y(_0__44_) );
INVX1 INVX1_62 ( .A(_32__3_), .Y(_497_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_498_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_499_) );
OAI21X1 OAI21X1_61 ( .A(_497_), .B(_499_), .C(_498_), .Y(_31_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_493_) );
NAND3X1 NAND3X1_28 ( .A(_497_), .B(_498_), .C(_493_), .Y(_494_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_495_) );
OAI21X1 OAI21X1_62 ( .A(_499_), .B(_495_), .C(_32__3_), .Y(_496_) );
NAND2X1 NAND2X1_69 ( .A(_496_), .B(_494_), .Y(_0__47_) );
INVX1 INVX1_63 ( .A(_32__1_), .Y(_504_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_505_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_506_) );
OAI21X1 OAI21X1_63 ( .A(_504_), .B(_506_), .C(_505_), .Y(_32__2_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_500_) );
NAND3X1 NAND3X1_29 ( .A(_504_), .B(_505_), .C(_500_), .Y(_501_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_502_) );
OAI21X1 OAI21X1_64 ( .A(_506_), .B(_502_), .C(_32__1_), .Y(_503_) );
NAND2X1 NAND2X1_71 ( .A(_503_), .B(_501_), .Y(_0__45_) );
INVX1 INVX1_64 ( .A(_32__2_), .Y(_511_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_512_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_513_) );
OAI21X1 OAI21X1_65 ( .A(_511_), .B(_513_), .C(_512_), .Y(_32__3_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_507_) );
NAND3X1 NAND3X1_30 ( .A(_511_), .B(_512_), .C(_507_), .Y(_508_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_509_) );
OAI21X1 OAI21X1_66 ( .A(_513_), .B(_509_), .C(_32__2_), .Y(_510_) );
NAND2X1 NAND2X1_73 ( .A(_510_), .B(_508_), .Y(_0__46_) );
INVX1 INVX1_65 ( .A(i_add_term1[44]), .Y(_514_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[44]), .B(_514_), .Y(_515_) );
INVX1 INVX1_66 ( .A(i_add_term2[44]), .Y(_516_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term1[44]), .B(_516_), .Y(_517_) );
INVX1 INVX1_67 ( .A(i_add_term1[45]), .Y(_518_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[45]), .B(_518_), .Y(_519_) );
INVX1 INVX1_68 ( .A(i_add_term2[45]), .Y(_520_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term1[45]), .B(_520_), .Y(_521_) );
OAI22X1 OAI22X1_8 ( .A(_515_), .B(_517_), .C(_519_), .D(_521_), .Y(_522_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_523_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_524_) );
NOR2X1 NOR2X1_84 ( .A(_523_), .B(_524_), .Y(_525_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_526_) );
NAND2X1 NAND2X1_74 ( .A(_525_), .B(_526_), .Y(_527_) );
NOR2X1 NOR2X1_85 ( .A(_522_), .B(_527_), .Y(_33_) );
INVX1 INVX1_69 ( .A(_31_), .Y(_528_) );
NAND2X1 NAND2X1_75 ( .A(1'b0), .B(_33_), .Y(_529_) );
OAI21X1 OAI21X1_67 ( .A(_33_), .B(_528_), .C(_529_), .Y(w_cout_11_) );
INVX1 INVX1_70 ( .A(w_cout_11_), .Y(_534_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_535_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_536_) );
OAI21X1 OAI21X1_68 ( .A(_534_), .B(_536_), .C(_535_), .Y(_35__1_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_530_) );
NAND3X1 NAND3X1_31 ( .A(_534_), .B(_535_), .C(_530_), .Y(_531_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_532_) );
OAI21X1 OAI21X1_69 ( .A(_536_), .B(_532_), .C(w_cout_11_), .Y(_533_) );
NAND2X1 NAND2X1_77 ( .A(_533_), .B(_531_), .Y(_0__48_) );
INVX1 INVX1_71 ( .A(_35__3_), .Y(_541_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_542_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_543_) );
OAI21X1 OAI21X1_70 ( .A(_541_), .B(_543_), .C(_542_), .Y(_34_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_537_) );
NAND3X1 NAND3X1_32 ( .A(_541_), .B(_542_), .C(_537_), .Y(_538_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_539_) );
OAI21X1 OAI21X1_71 ( .A(_543_), .B(_539_), .C(_35__3_), .Y(_540_) );
NAND2X1 NAND2X1_79 ( .A(_540_), .B(_538_), .Y(_0__51_) );
INVX1 INVX1_72 ( .A(_35__1_), .Y(_548_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_549_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_550_) );
OAI21X1 OAI21X1_72 ( .A(_548_), .B(_550_), .C(_549_), .Y(_35__2_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_544_) );
NAND3X1 NAND3X1_33 ( .A(_548_), .B(_549_), .C(_544_), .Y(_545_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_546_) );
OAI21X1 OAI21X1_73 ( .A(_550_), .B(_546_), .C(_35__1_), .Y(_547_) );
NAND2X1 NAND2X1_81 ( .A(_547_), .B(_545_), .Y(_0__49_) );
INVX1 INVX1_73 ( .A(_35__2_), .Y(_555_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_556_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_557_) );
OAI21X1 OAI21X1_74 ( .A(_555_), .B(_557_), .C(_556_), .Y(_35__3_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_551_) );
NAND3X1 NAND3X1_34 ( .A(_555_), .B(_556_), .C(_551_), .Y(_552_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_553_) );
OAI21X1 OAI21X1_75 ( .A(_557_), .B(_553_), .C(_35__2_), .Y(_554_) );
NAND2X1 NAND2X1_83 ( .A(_554_), .B(_552_), .Y(_0__50_) );
INVX1 INVX1_74 ( .A(i_add_term1[48]), .Y(_558_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[48]), .B(_558_), .Y(_559_) );
INVX1 INVX1_75 ( .A(i_add_term2[48]), .Y(_560_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term1[48]), .B(_560_), .Y(_561_) );
INVX1 INVX1_76 ( .A(i_add_term1[49]), .Y(_562_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[49]), .B(_562_), .Y(_563_) );
INVX1 INVX1_77 ( .A(i_add_term2[49]), .Y(_564_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term1[49]), .B(_564_), .Y(_565_) );
OAI22X1 OAI22X1_9 ( .A(_559_), .B(_561_), .C(_563_), .D(_565_), .Y(_566_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_567_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_568_) );
NOR2X1 NOR2X1_95 ( .A(_567_), .B(_568_), .Y(_569_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_570_) );
NAND2X1 NAND2X1_84 ( .A(_569_), .B(_570_), .Y(_571_) );
NOR2X1 NOR2X1_96 ( .A(_566_), .B(_571_), .Y(_36_) );
INVX1 INVX1_78 ( .A(_34_), .Y(_572_) );
NAND2X1 NAND2X1_85 ( .A(1'b0), .B(_36_), .Y(_573_) );
OAI21X1 OAI21X1_76 ( .A(_36_), .B(_572_), .C(_573_), .Y(w_cout_12_) );
INVX1 INVX1_79 ( .A(w_cout_12_), .Y(_578_) );
NAND2X1 NAND2X1_86 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_579_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_580_) );
OAI21X1 OAI21X1_77 ( .A(_578_), .B(_580_), .C(_579_), .Y(_38__1_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_574_) );
NAND3X1 NAND3X1_35 ( .A(_578_), .B(_579_), .C(_574_), .Y(_575_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_576_) );
OAI21X1 OAI21X1_78 ( .A(_580_), .B(_576_), .C(w_cout_12_), .Y(_577_) );
NAND2X1 NAND2X1_87 ( .A(_577_), .B(_575_), .Y(_0__52_) );
INVX1 INVX1_80 ( .A(_38__3_), .Y(_585_) );
NAND2X1 NAND2X1_88 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_586_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_587_) );
OAI21X1 OAI21X1_79 ( .A(_585_), .B(_587_), .C(_586_), .Y(_37_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_581_) );
NAND3X1 NAND3X1_36 ( .A(_585_), .B(_586_), .C(_581_), .Y(_582_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_583_) );
OAI21X1 OAI21X1_80 ( .A(_587_), .B(_583_), .C(_38__3_), .Y(_584_) );
NAND2X1 NAND2X1_89 ( .A(_584_), .B(_582_), .Y(_0__55_) );
INVX1 INVX1_81 ( .A(_38__1_), .Y(_592_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_593_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_594_) );
OAI21X1 OAI21X1_81 ( .A(_592_), .B(_594_), .C(_593_), .Y(_38__2_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_588_) );
NAND3X1 NAND3X1_37 ( .A(_592_), .B(_593_), .C(_588_), .Y(_589_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_590_) );
OAI21X1 OAI21X1_82 ( .A(_594_), .B(_590_), .C(_38__1_), .Y(_591_) );
NAND2X1 NAND2X1_91 ( .A(_591_), .B(_589_), .Y(_0__53_) );
INVX1 INVX1_82 ( .A(_38__2_), .Y(_599_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_600_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_601_) );
OAI21X1 OAI21X1_83 ( .A(_599_), .B(_601_), .C(_600_), .Y(_38__3_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_595_) );
NAND3X1 NAND3X1_38 ( .A(_599_), .B(_600_), .C(_595_), .Y(_596_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_597_) );
OAI21X1 OAI21X1_84 ( .A(_601_), .B(_597_), .C(_38__2_), .Y(_598_) );
NAND2X1 NAND2X1_93 ( .A(_598_), .B(_596_), .Y(_0__54_) );
INVX1 INVX1_83 ( .A(i_add_term1[52]), .Y(_602_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[52]), .B(_602_), .Y(_603_) );
INVX1 INVX1_84 ( .A(i_add_term2[52]), .Y(_604_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term1[52]), .B(_604_), .Y(_605_) );
INVX1 INVX1_85 ( .A(i_add_term1[53]), .Y(_606_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[53]), .B(_606_), .Y(_607_) );
INVX1 INVX1_86 ( .A(i_add_term2[53]), .Y(_608_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term1[53]), .B(_608_), .Y(_609_) );
OAI22X1 OAI22X1_10 ( .A(_603_), .B(_605_), .C(_607_), .D(_609_), .Y(_610_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_611_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_612_) );
NOR2X1 NOR2X1_106 ( .A(_611_), .B(_612_), .Y(_613_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_614_) );
NAND2X1 NAND2X1_94 ( .A(_613_), .B(_614_), .Y(_615_) );
NOR2X1 NOR2X1_107 ( .A(_610_), .B(_615_), .Y(_39_) );
INVX1 INVX1_87 ( .A(_37_), .Y(_616_) );
NAND2X1 NAND2X1_95 ( .A(1'b0), .B(_39_), .Y(_617_) );
OAI21X1 OAI21X1_85 ( .A(_39_), .B(_616_), .C(_617_), .Y(w_cout_13_) );
INVX1 INVX1_88 ( .A(w_cout_13_), .Y(_622_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_623_) );
NOR2X1 NOR2X1_108 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_624_) );
OAI21X1 OAI21X1_86 ( .A(_622_), .B(_624_), .C(_623_), .Y(_41__1_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_618_) );
NAND3X1 NAND3X1_39 ( .A(_622_), .B(_623_), .C(_618_), .Y(_619_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_620_) );
OAI21X1 OAI21X1_87 ( .A(_624_), .B(_620_), .C(w_cout_13_), .Y(_621_) );
NAND2X1 NAND2X1_97 ( .A(_621_), .B(_619_), .Y(_0__56_) );
INVX1 INVX1_89 ( .A(_41__3_), .Y(_629_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_630_) );
NOR2X1 NOR2X1_109 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_631_) );
OAI21X1 OAI21X1_88 ( .A(_629_), .B(_631_), .C(_630_), .Y(_40_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_625_) );
NAND3X1 NAND3X1_40 ( .A(_629_), .B(_630_), .C(_625_), .Y(_626_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_627_) );
OAI21X1 OAI21X1_89 ( .A(_631_), .B(_627_), .C(_41__3_), .Y(_628_) );
NAND2X1 NAND2X1_99 ( .A(_628_), .B(_626_), .Y(_0__59_) );
INVX1 INVX1_90 ( .A(_41__1_), .Y(_636_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_637_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_638_) );
OAI21X1 OAI21X1_90 ( .A(_636_), .B(_638_), .C(_637_), .Y(_41__2_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_632_) );
NAND3X1 NAND3X1_41 ( .A(_636_), .B(_637_), .C(_632_), .Y(_633_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_634_) );
OAI21X1 OAI21X1_91 ( .A(_638_), .B(_634_), .C(_41__1_), .Y(_635_) );
NAND2X1 NAND2X1_101 ( .A(_635_), .B(_633_), .Y(_0__57_) );
INVX1 INVX1_91 ( .A(_41__2_), .Y(_643_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_644_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_645_) );
OAI21X1 OAI21X1_92 ( .A(_643_), .B(_645_), .C(_644_), .Y(_41__3_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_639_) );
NAND3X1 NAND3X1_42 ( .A(_643_), .B(_644_), .C(_639_), .Y(_640_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_641_) );
OAI21X1 OAI21X1_93 ( .A(_645_), .B(_641_), .C(_41__2_), .Y(_642_) );
NAND2X1 NAND2X1_103 ( .A(_642_), .B(_640_), .Y(_0__58_) );
INVX1 INVX1_92 ( .A(i_add_term1[56]), .Y(_646_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term2[56]), .B(_646_), .Y(_647_) );
INVX1 INVX1_93 ( .A(i_add_term2[56]), .Y(_648_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term1[56]), .B(_648_), .Y(_649_) );
INVX1 INVX1_94 ( .A(i_add_term1[57]), .Y(_650_) );
NOR2X1 NOR2X1_114 ( .A(i_add_term2[57]), .B(_650_), .Y(_651_) );
INVX1 INVX1_95 ( .A(i_add_term2[57]), .Y(_652_) );
NOR2X1 NOR2X1_115 ( .A(i_add_term1[57]), .B(_652_), .Y(_653_) );
OAI22X1 OAI22X1_11 ( .A(_647_), .B(_649_), .C(_651_), .D(_653_), .Y(_654_) );
NOR2X1 NOR2X1_116 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_655_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_656_) );
NOR2X1 NOR2X1_117 ( .A(_655_), .B(_656_), .Y(_657_) );
XOR2X1 XOR2X1_11 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_658_) );
NAND2X1 NAND2X1_104 ( .A(_657_), .B(_658_), .Y(_659_) );
NOR2X1 NOR2X1_118 ( .A(_654_), .B(_659_), .Y(_42_) );
INVX1 INVX1_96 ( .A(_40_), .Y(_660_) );
NAND2X1 NAND2X1_105 ( .A(1'b0), .B(_42_), .Y(_661_) );
OAI21X1 OAI21X1_94 ( .A(_42_), .B(_660_), .C(_661_), .Y(w_cout_14_) );
INVX1 INVX1_97 ( .A(w_cout_14_), .Y(_666_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_667_) );
NOR2X1 NOR2X1_119 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_668_) );
OAI21X1 OAI21X1_95 ( .A(_666_), .B(_668_), .C(_667_), .Y(_44__1_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_662_) );
NAND3X1 NAND3X1_43 ( .A(_666_), .B(_667_), .C(_662_), .Y(_663_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_664_) );
OAI21X1 OAI21X1_96 ( .A(_668_), .B(_664_), .C(w_cout_14_), .Y(_665_) );
NAND2X1 NAND2X1_107 ( .A(_665_), .B(_663_), .Y(_0__60_) );
INVX1 INVX1_98 ( .A(_44__3_), .Y(_673_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_674_) );
NOR2X1 NOR2X1_120 ( .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_675_) );
OAI21X1 OAI21X1_97 ( .A(_673_), .B(_675_), .C(_674_), .Y(_43_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_669_) );
NAND3X1 NAND3X1_44 ( .A(_673_), .B(_674_), .C(_669_), .Y(_670_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_671_) );
OAI21X1 OAI21X1_98 ( .A(_675_), .B(_671_), .C(_44__3_), .Y(_672_) );
NAND2X1 NAND2X1_109 ( .A(_672_), .B(_670_), .Y(_0__63_) );
INVX1 INVX1_99 ( .A(_44__1_), .Y(_680_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_681_) );
NOR2X1 NOR2X1_121 ( .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_682_) );
OAI21X1 OAI21X1_99 ( .A(_680_), .B(_682_), .C(_681_), .Y(_44__2_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_676_) );
NAND3X1 NAND3X1_45 ( .A(_680_), .B(_681_), .C(_676_), .Y(_677_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_678_) );
OAI21X1 OAI21X1_100 ( .A(_682_), .B(_678_), .C(_44__1_), .Y(_679_) );
NAND2X1 NAND2X1_111 ( .A(_679_), .B(_677_), .Y(_0__61_) );
INVX1 INVX1_100 ( .A(_44__2_), .Y(_687_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_688_) );
NOR2X1 NOR2X1_122 ( .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_689_) );
OAI21X1 OAI21X1_101 ( .A(_687_), .B(_689_), .C(_688_), .Y(_44__3_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_683_) );
NAND3X1 NAND3X1_46 ( .A(_687_), .B(_688_), .C(_683_), .Y(_684_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_685_) );
OAI21X1 OAI21X1_102 ( .A(_689_), .B(_685_), .C(_44__2_), .Y(_686_) );
NAND2X1 NAND2X1_113 ( .A(_686_), .B(_684_), .Y(_0__62_) );
INVX1 INVX1_101 ( .A(i_add_term1[60]), .Y(_690_) );
NOR2X1 NOR2X1_123 ( .A(i_add_term2[60]), .B(_690_), .Y(_691_) );
INVX1 INVX1_102 ( .A(i_add_term2[60]), .Y(_692_) );
NOR2X1 NOR2X1_124 ( .A(i_add_term1[60]), .B(_692_), .Y(_693_) );
INVX1 INVX1_103 ( .A(i_add_term1[61]), .Y(_694_) );
NOR2X1 NOR2X1_125 ( .A(i_add_term2[61]), .B(_694_), .Y(_695_) );
INVX1 INVX1_104 ( .A(i_add_term2[61]), .Y(_696_) );
NOR2X1 NOR2X1_126 ( .A(i_add_term1[61]), .B(_696_), .Y(_697_) );
OAI22X1 OAI22X1_12 ( .A(_691_), .B(_693_), .C(_695_), .D(_697_), .Y(_698_) );
NOR2X1 NOR2X1_127 ( .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_699_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_700_) );
NOR2X1 NOR2X1_128 ( .A(_699_), .B(_700_), .Y(_701_) );
XOR2X1 XOR2X1_12 ( .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_702_) );
NAND2X1 NAND2X1_114 ( .A(_701_), .B(_702_), .Y(_703_) );
NOR2X1 NOR2X1_129 ( .A(_698_), .B(_703_), .Y(_45_) );
INVX1 INVX1_105 ( .A(_43_), .Y(_704_) );
NAND2X1 NAND2X1_115 ( .A(1'b0), .B(_45_), .Y(_705_) );
OAI21X1 OAI21X1_103 ( .A(_45_), .B(_704_), .C(_705_), .Y(w_cout_15_) );
INVX1 INVX1_106 ( .A(1'b0), .Y(_710_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_711_) );
NOR2X1 NOR2X1_130 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_712_) );
OAI21X1 OAI21X1_104 ( .A(_710_), .B(_712_), .C(_711_), .Y(rca_inst_fa0_o_carry) );
OR2X2 OR2X2_46 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_706_) );
NAND3X1 NAND3X1_47 ( .A(_710_), .B(_711_), .C(_706_), .Y(_707_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_708_) );
OAI21X1 OAI21X1_105 ( .A(_712_), .B(_708_), .C(1'b0), .Y(_709_) );
NAND2X1 NAND2X1_117 ( .A(_709_), .B(_707_), .Y(rca_inst_fa0_o_sum) );
INVX1 INVX1_107 ( .A(rca_inst_fa3_i_carry), .Y(_717_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_718_) );
NOR2X1 NOR2X1_131 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_719_) );
OAI21X1 OAI21X1_106 ( .A(_717_), .B(_719_), .C(_718_), .Y(cout0) );
OR2X2 OR2X2_47 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_713_) );
NAND3X1 NAND3X1_48 ( .A(_717_), .B(_718_), .C(_713_), .Y(_714_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_715_) );
OAI21X1 OAI21X1_107 ( .A(_719_), .B(_715_), .C(rca_inst_fa3_i_carry), .Y(_716_) );
NAND2X1 NAND2X1_119 ( .A(_716_), .B(_714_), .Y(rca_inst_fa3_o_sum) );
INVX1 INVX1_108 ( .A(rca_inst_fa0_o_carry), .Y(_724_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_725_) );
NOR2X1 NOR2X1_132 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_726_) );
OAI21X1 OAI21X1_108 ( .A(_724_), .B(_726_), .C(_725_), .Y(rca_inst_fa_1__o_carry) );
OR2X2 OR2X2_48 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_720_) );
NAND3X1 NAND3X1_49 ( .A(_724_), .B(_725_), .C(_720_), .Y(_721_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_722_) );
OAI21X1 OAI21X1_109 ( .A(_726_), .B(_722_), .C(rca_inst_fa0_o_carry), .Y(_723_) );
NAND2X1 NAND2X1_121 ( .A(_723_), .B(_721_), .Y(rca_inst_fa_1__o_sum) );
INVX1 INVX1_109 ( .A(rca_inst_fa_1__o_carry), .Y(_731_) );
NAND2X1 NAND2X1_122 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_732_) );
NOR2X1 NOR2X1_133 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_733_) );
OAI21X1 OAI21X1_110 ( .A(_731_), .B(_733_), .C(_732_), .Y(rca_inst_fa3_i_carry) );
OR2X2 OR2X2_49 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_727_) );
NAND3X1 NAND3X1_50 ( .A(_731_), .B(_732_), .C(_727_), .Y(_728_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_729_) );
OAI21X1 OAI21X1_111 ( .A(_733_), .B(_729_), .C(rca_inst_fa_1__o_carry), .Y(_730_) );
NAND2X1 NAND2X1_123 ( .A(_730_), .B(_728_), .Y(rca_inst_fa_2__o_sum) );
INVX1 INVX1_110 ( .A(i_add_term1[0]), .Y(_734_) );
NOR2X1 NOR2X1_134 ( .A(i_add_term2[0]), .B(_734_), .Y(_735_) );
INVX1 INVX1_111 ( .A(i_add_term2[0]), .Y(_736_) );
NOR2X1 NOR2X1_135 ( .A(i_add_term1[0]), .B(_736_), .Y(_737_) );
INVX1 INVX1_112 ( .A(i_add_term1[1]), .Y(_738_) );
NOR2X1 NOR2X1_136 ( .A(i_add_term2[1]), .B(_738_), .Y(_739_) );
INVX1 INVX1_113 ( .A(i_add_term2[1]), .Y(_740_) );
NOR2X1 NOR2X1_137 ( .A(i_add_term1[1]), .B(_740_), .Y(_741_) );
OAI22X1 OAI22X1_13 ( .A(_735_), .B(_737_), .C(_739_), .D(_741_), .Y(_742_) );
NOR2X1 NOR2X1_138 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_743_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_744_) );
NOR2X1 NOR2X1_139 ( .A(_743_), .B(_744_), .Y(_745_) );
XOR2X1 XOR2X1_13 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_746_) );
NAND2X1 NAND2X1_124 ( .A(_745_), .B(_746_), .Y(_747_) );
NOR2X1 NOR2X1_140 ( .A(_742_), .B(_747_), .Y(skip0_P) );
INVX1 INVX1_114 ( .A(cout0), .Y(_748_) );
NAND2X1 NAND2X1_125 ( .A(1'b0), .B(skip0_P), .Y(_749_) );
OAI21X1 OAI21X1_112 ( .A(skip0_P), .B(_748_), .C(_749_), .Y(skip0_cin_next) );
BUFX2 BUFX2_1 ( .A(w_cout_15_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .A(_0__54_), .Y(sum[54]) );
BUFX2 BUFX2_57 ( .A(_0__55_), .Y(sum[55]) );
BUFX2 BUFX2_58 ( .A(_0__56_), .Y(sum[56]) );
BUFX2 BUFX2_59 ( .A(_0__57_), .Y(sum[57]) );
BUFX2 BUFX2_60 ( .A(_0__58_), .Y(sum[58]) );
BUFX2 BUFX2_61 ( .A(_0__59_), .Y(sum[59]) );
BUFX2 BUFX2_62 ( .A(_0__60_), .Y(sum[60]) );
BUFX2 BUFX2_63 ( .A(_0__61_), .Y(sum[61]) );
BUFX2 BUFX2_64 ( .A(_0__62_), .Y(sum[62]) );
BUFX2 BUFX2_65 ( .A(_0__63_), .Y(sum[63]) );
INVX1 INVX1_115 ( .A(skip0_cin_next), .Y(_50_) );
NAND2X1 NAND2X1_126 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_51_) );
NOR2X1 NOR2X1_141 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_52_) );
OAI21X1 OAI21X1_113 ( .A(_50_), .B(_52_), .C(_51_), .Y(_2__1_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_46_) );
NAND3X1 NAND3X1_51 ( .A(_50_), .B(_51_), .C(_46_), .Y(_47_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_48_) );
OAI21X1 OAI21X1_114 ( .A(_52_), .B(_48_), .C(skip0_cin_next), .Y(_49_) );
NAND2X1 NAND2X1_127 ( .A(_49_), .B(_47_), .Y(_0__4_) );
INVX1 INVX1_116 ( .A(_2__3_), .Y(_57_) );
NAND2X1 NAND2X1_128 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_58_) );
NOR2X1 NOR2X1_142 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_59_) );
OAI21X1 OAI21X1_115 ( .A(_57_), .B(_59_), .C(_58_), .Y(_1_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_53_) );
NAND3X1 NAND3X1_52 ( .A(_57_), .B(_58_), .C(_53_), .Y(_54_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_55_) );
OAI21X1 OAI21X1_116 ( .A(_59_), .B(_55_), .C(_2__3_), .Y(_56_) );
NAND2X1 NAND2X1_129 ( .A(_56_), .B(_54_), .Y(_0__7_) );
INVX1 INVX1_117 ( .A(_2__1_), .Y(_64_) );
NAND2X1 NAND2X1_130 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_65_) );
NOR2X1 NOR2X1_143 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_66_) );
OAI21X1 OAI21X1_117 ( .A(_64_), .B(_66_), .C(_65_), .Y(_2__2_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_60_) );
NAND3X1 NAND3X1_53 ( .A(_64_), .B(_65_), .C(_60_), .Y(_61_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_62_) );
OAI21X1 OAI21X1_118 ( .A(_66_), .B(_62_), .C(_2__1_), .Y(_63_) );
NAND2X1 NAND2X1_131 ( .A(_63_), .B(_61_), .Y(_0__5_) );
INVX1 INVX1_118 ( .A(_2__2_), .Y(_71_) );
NAND2X1 NAND2X1_132 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_72_) );
NOR2X1 NOR2X1_144 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_73_) );
OAI21X1 OAI21X1_119 ( .A(_71_), .B(_73_), .C(_72_), .Y(_2__3_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_67_) );
NAND3X1 NAND3X1_54 ( .A(_71_), .B(_72_), .C(_67_), .Y(_68_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_69_) );
OAI21X1 OAI21X1_120 ( .A(_73_), .B(_69_), .C(_2__2_), .Y(_70_) );
NAND2X1 NAND2X1_133 ( .A(_70_), .B(_68_), .Y(_0__6_) );
INVX1 INVX1_119 ( .A(i_add_term1[4]), .Y(_74_) );
NOR2X1 NOR2X1_145 ( .A(i_add_term2[4]), .B(_74_), .Y(_75_) );
INVX1 INVX1_120 ( .A(i_add_term2[4]), .Y(_76_) );
NOR2X1 NOR2X1_146 ( .A(i_add_term1[4]), .B(_76_), .Y(_77_) );
INVX1 INVX1_121 ( .A(i_add_term1[5]), .Y(_78_) );
NOR2X1 NOR2X1_147 ( .A(i_add_term2[5]), .B(_78_), .Y(_79_) );
INVX1 INVX1_122 ( .A(i_add_term2[5]), .Y(_80_) );
NOR2X1 NOR2X1_148 ( .A(i_add_term1[5]), .B(_80_), .Y(_81_) );
OAI22X1 OAI22X1_14 ( .A(_75_), .B(_77_), .C(_79_), .D(_81_), .Y(_82_) );
NOR2X1 NOR2X1_149 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_83_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_84_) );
NOR2X1 NOR2X1_150 ( .A(_83_), .B(_84_), .Y(_85_) );
XOR2X1 XOR2X1_14 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_86_) );
NAND2X1 NAND2X1_134 ( .A(_85_), .B(_86_), .Y(_87_) );
NOR2X1 NOR2X1_151 ( .A(_82_), .B(_87_), .Y(_3_) );
INVX1 INVX1_123 ( .A(_1_), .Y(_88_) );
NAND2X1 NAND2X1_135 ( .A(1'b0), .B(_3_), .Y(_89_) );
OAI21X1 OAI21X1_121 ( .A(_3_), .B(_88_), .C(_89_), .Y(w_cout_1_) );
INVX1 INVX1_124 ( .A(w_cout_1_), .Y(_94_) );
NAND2X1 NAND2X1_136 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_95_) );
NOR2X1 NOR2X1_152 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_96_) );
OAI21X1 OAI21X1_122 ( .A(_94_), .B(_96_), .C(_95_), .Y(_5__1_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_90_) );
NAND3X1 NAND3X1_55 ( .A(_94_), .B(_95_), .C(_90_), .Y(_91_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_92_) );
OAI21X1 OAI21X1_123 ( .A(_96_), .B(_92_), .C(w_cout_1_), .Y(_93_) );
NAND2X1 NAND2X1_137 ( .A(_93_), .B(_91_), .Y(_0__8_) );
INVX1 INVX1_125 ( .A(_5__3_), .Y(_101_) );
NAND2X1 NAND2X1_138 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_102_) );
NOR2X1 NOR2X1_153 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_103_) );
OAI21X1 OAI21X1_124 ( .A(_101_), .B(_103_), .C(_102_), .Y(_4_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_97_) );
NAND3X1 NAND3X1_56 ( .A(_101_), .B(_102_), .C(_97_), .Y(_98_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_99_) );
OAI21X1 OAI21X1_125 ( .A(_103_), .B(_99_), .C(_5__3_), .Y(_100_) );
NAND2X1 NAND2X1_139 ( .A(_100_), .B(_98_), .Y(_0__11_) );
INVX1 INVX1_126 ( .A(_5__1_), .Y(_108_) );
NAND2X1 NAND2X1_140 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_109_) );
NOR2X1 NOR2X1_154 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_110_) );
OAI21X1 OAI21X1_126 ( .A(_108_), .B(_110_), .C(_109_), .Y(_5__2_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_104_) );
NAND3X1 NAND3X1_57 ( .A(_108_), .B(_109_), .C(_104_), .Y(_105_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_106_) );
OAI21X1 OAI21X1_127 ( .A(_110_), .B(_106_), .C(_5__1_), .Y(_107_) );
NAND2X1 NAND2X1_141 ( .A(_107_), .B(_105_), .Y(_0__9_) );
INVX1 INVX1_127 ( .A(_5__2_), .Y(_115_) );
NAND2X1 NAND2X1_142 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_116_) );
NOR2X1 NOR2X1_155 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_117_) );
OAI21X1 OAI21X1_128 ( .A(_115_), .B(_117_), .C(_116_), .Y(_5__3_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_111_) );
NAND3X1 NAND3X1_58 ( .A(_115_), .B(_116_), .C(_111_), .Y(_112_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_113_) );
OAI21X1 OAI21X1_129 ( .A(_117_), .B(_113_), .C(_5__2_), .Y(_114_) );
NAND2X1 NAND2X1_143 ( .A(_114_), .B(_112_), .Y(_0__10_) );
INVX1 INVX1_128 ( .A(i_add_term1[8]), .Y(_118_) );
NOR2X1 NOR2X1_156 ( .A(i_add_term2[8]), .B(_118_), .Y(_119_) );
INVX1 INVX1_129 ( .A(i_add_term2[8]), .Y(_120_) );
NOR2X1 NOR2X1_157 ( .A(i_add_term1[8]), .B(_120_), .Y(_121_) );
INVX1 INVX1_130 ( .A(i_add_term1[9]), .Y(_122_) );
NOR2X1 NOR2X1_158 ( .A(i_add_term2[9]), .B(_122_), .Y(_123_) );
INVX1 INVX1_131 ( .A(i_add_term2[9]), .Y(_124_) );
NOR2X1 NOR2X1_159 ( .A(i_add_term1[9]), .B(_124_), .Y(_125_) );
OAI22X1 OAI22X1_15 ( .A(_119_), .B(_121_), .C(_123_), .D(_125_), .Y(_126_) );
NOR2X1 NOR2X1_160 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_127_) );
AND2X2 AND2X2_73 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_128_) );
NOR2X1 NOR2X1_161 ( .A(_127_), .B(_128_), .Y(_129_) );
XOR2X1 XOR2X1_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_130_) );
NAND2X1 NAND2X1_144 ( .A(_129_), .B(_130_), .Y(_131_) );
NOR2X1 NOR2X1_162 ( .A(_126_), .B(_131_), .Y(_6_) );
INVX1 INVX1_132 ( .A(_4_), .Y(_132_) );
NAND2X1 NAND2X1_145 ( .A(1'b0), .B(_6_), .Y(_133_) );
OAI21X1 OAI21X1_130 ( .A(_6_), .B(_132_), .C(_133_), .Y(w_cout_2_) );
INVX1 INVX1_133 ( .A(w_cout_2_), .Y(_138_) );
NAND2X1 NAND2X1_146 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_139_) );
NOR2X1 NOR2X1_163 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_140_) );
OAI21X1 OAI21X1_131 ( .A(_138_), .B(_140_), .C(_139_), .Y(_8__1_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_134_) );
NAND3X1 NAND3X1_59 ( .A(_138_), .B(_139_), .C(_134_), .Y(_135_) );
AND2X2 AND2X2_74 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_136_) );
OAI21X1 OAI21X1_132 ( .A(_140_), .B(_136_), .C(w_cout_2_), .Y(_137_) );
NAND2X1 NAND2X1_147 ( .A(_137_), .B(_135_), .Y(_0__12_) );
INVX1 INVX1_134 ( .A(_8__3_), .Y(_145_) );
NAND2X1 NAND2X1_148 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_146_) );
NOR2X1 NOR2X1_164 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_147_) );
OAI21X1 OAI21X1_133 ( .A(_145_), .B(_147_), .C(_146_), .Y(_7_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_141_) );
NAND3X1 NAND3X1_60 ( .A(_145_), .B(_146_), .C(_141_), .Y(_142_) );
AND2X2 AND2X2_75 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_143_) );
OAI21X1 OAI21X1_134 ( .A(_147_), .B(_143_), .C(_8__3_), .Y(_144_) );
NAND2X1 NAND2X1_149 ( .A(_144_), .B(_142_), .Y(_0__15_) );
INVX1 INVX1_135 ( .A(_8__1_), .Y(_152_) );
NAND2X1 NAND2X1_150 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_153_) );
NOR2X1 NOR2X1_165 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_154_) );
OAI21X1 OAI21X1_135 ( .A(_152_), .B(_154_), .C(_153_), .Y(_8__2_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_148_) );
NAND3X1 NAND3X1_61 ( .A(_152_), .B(_153_), .C(_148_), .Y(_149_) );
AND2X2 AND2X2_76 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_150_) );
OAI21X1 OAI21X1_136 ( .A(_154_), .B(_150_), .C(_8__1_), .Y(_151_) );
NAND2X1 NAND2X1_151 ( .A(_151_), .B(_149_), .Y(_0__13_) );
INVX1 INVX1_136 ( .A(_8__2_), .Y(_159_) );
NAND2X1 NAND2X1_152 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_160_) );
NOR2X1 NOR2X1_166 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_161_) );
OAI21X1 OAI21X1_137 ( .A(_159_), .B(_161_), .C(_160_), .Y(_8__3_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_155_) );
NAND3X1 NAND3X1_62 ( .A(_159_), .B(_160_), .C(_155_), .Y(_156_) );
AND2X2 AND2X2_77 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_157_) );
OAI21X1 OAI21X1_138 ( .A(_161_), .B(_157_), .C(_8__2_), .Y(_158_) );
NAND2X1 NAND2X1_153 ( .A(_158_), .B(_156_), .Y(_0__14_) );
INVX1 INVX1_137 ( .A(i_add_term1[12]), .Y(_162_) );
NOR2X1 NOR2X1_167 ( .A(i_add_term2[12]), .B(_162_), .Y(_163_) );
INVX1 INVX1_138 ( .A(i_add_term2[12]), .Y(_164_) );
NOR2X1 NOR2X1_168 ( .A(i_add_term1[12]), .B(_164_), .Y(_165_) );
INVX1 INVX1_139 ( .A(i_add_term1[13]), .Y(_166_) );
NOR2X1 NOR2X1_169 ( .A(i_add_term2[13]), .B(_166_), .Y(_167_) );
INVX1 INVX1_140 ( .A(i_add_term2[13]), .Y(_168_) );
NOR2X1 NOR2X1_170 ( .A(i_add_term1[13]), .B(_168_), .Y(_169_) );
OAI22X1 OAI22X1_16 ( .A(_163_), .B(_165_), .C(_167_), .D(_169_), .Y(_170_) );
NOR2X1 NOR2X1_171 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_171_) );
AND2X2 AND2X2_78 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_172_) );
NOR2X1 NOR2X1_172 ( .A(_171_), .B(_172_), .Y(_173_) );
XOR2X1 XOR2X1_16 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_174_) );
NAND2X1 NAND2X1_154 ( .A(_173_), .B(_174_), .Y(_175_) );
NOR2X1 NOR2X1_173 ( .A(_170_), .B(_175_), .Y(_9_) );
INVX1 INVX1_141 ( .A(_7_), .Y(_176_) );
NAND2X1 NAND2X1_155 ( .A(1'b0), .B(_9_), .Y(_177_) );
OAI21X1 OAI21X1_139 ( .A(_9_), .B(_176_), .C(_177_), .Y(w_cout_3_) );
INVX1 INVX1_142 ( .A(w_cout_3_), .Y(_182_) );
NAND2X1 NAND2X1_156 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_183_) );
NOR2X1 NOR2X1_174 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_184_) );
OAI21X1 OAI21X1_140 ( .A(_182_), .B(_184_), .C(_183_), .Y(_11__1_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_178_) );
NAND3X1 NAND3X1_63 ( .A(_182_), .B(_183_), .C(_178_), .Y(_179_) );
AND2X2 AND2X2_79 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_180_) );
OAI21X1 OAI21X1_141 ( .A(_184_), .B(_180_), .C(w_cout_3_), .Y(_181_) );
NAND2X1 NAND2X1_157 ( .A(_181_), .B(_179_), .Y(_0__16_) );
INVX1 INVX1_143 ( .A(_11__3_), .Y(_189_) );
NAND2X1 NAND2X1_158 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_190_) );
NOR2X1 NOR2X1_175 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_191_) );
OAI21X1 OAI21X1_142 ( .A(_189_), .B(_191_), .C(_190_), .Y(_10_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_185_) );
NAND3X1 NAND3X1_64 ( .A(_189_), .B(_190_), .C(_185_), .Y(_186_) );
AND2X2 AND2X2_80 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_187_) );
OAI21X1 OAI21X1_143 ( .A(_191_), .B(_187_), .C(_11__3_), .Y(_188_) );
NAND2X1 NAND2X1_159 ( .A(_188_), .B(_186_), .Y(_0__19_) );
INVX1 INVX1_144 ( .A(_11__1_), .Y(_196_) );
NAND2X1 NAND2X1_160 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_197_) );
NOR2X1 NOR2X1_176 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_198_) );
OAI21X1 OAI21X1_144 ( .A(_196_), .B(_198_), .C(_197_), .Y(_11__2_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_192_) );
BUFX2 BUFX2_66 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_67 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_68 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_69 ( .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_70 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
