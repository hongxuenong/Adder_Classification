module CSkipA_9bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [8:0] i_add_term1;
input [8:0] i_add_term2;
output [8:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX2 BUFX2_1 ( .A(cskip1_inst_sum), .Y(sum[8]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_5_) );
OAI21X1 OAI21X1_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .C(gnd), .Y(_6_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_7_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_8_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_9_) );
NAND3X1 NAND3X1_1 ( .A(_7_), .B(_8_), .C(_9_), .Y(_10_) );
OAI21X1 OAI21X1_2 ( .A(_6_), .B(_10_), .C(_5_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3_), .Y(_11_) );
OAI21X1 OAI21X1_3 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .C(gnd), .Y(_12_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_13_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_14_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_15_) );
NAND3X1 NAND3X1_2 ( .A(_13_), .B(_14_), .C(_15_), .Y(_16_) );
OAI21X1 OAI21X1_4 ( .A(_12_), .B(_16_), .C(_11_), .Y(cskip1_inst_cin) );
INVX1 INVX1_3 ( .A(gnd), .Y(_20_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_21_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_22_) );
NAND3X1 NAND3X1_3 ( .A(_20_), .B(_22_), .C(_21_), .Y(_23_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_17_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_18_) );
OAI21X1 OAI21X1_5 ( .A(_17_), .B(_18_), .C(gnd), .Y(_19_) );
NAND2X1 NAND2X1_2 ( .A(_19_), .B(_23_), .Y(_0__0_) );
OAI21X1 OAI21X1_6 ( .A(_20_), .B(_17_), .C(_22_), .Y(_2__1_) );
INVX1 INVX1_4 ( .A(_2__1_), .Y(_27_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_28_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_29_) );
NAND3X1 NAND3X1_4 ( .A(_27_), .B(_29_), .C(_28_), .Y(_30_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_24_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_25_) );
OAI21X1 OAI21X1_7 ( .A(_24_), .B(_25_), .C(_2__1_), .Y(_26_) );
NAND2X1 NAND2X1_4 ( .A(_26_), .B(_30_), .Y(_0__1_) );
OAI21X1 OAI21X1_8 ( .A(_27_), .B(_24_), .C(_29_), .Y(_2__2_) );
INVX1 INVX1_5 ( .A(_2__2_), .Y(_34_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_35_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_36_) );
NAND3X1 NAND3X1_5 ( .A(_34_), .B(_36_), .C(_35_), .Y(_37_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_31_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_32_) );
OAI21X1 OAI21X1_9 ( .A(_31_), .B(_32_), .C(_2__2_), .Y(_33_) );
NAND2X1 NAND2X1_6 ( .A(_33_), .B(_37_), .Y(_0__2_) );
OAI21X1 OAI21X1_10 ( .A(_34_), .B(_31_), .C(_36_), .Y(_2__3_) );
INVX1 INVX1_6 ( .A(_2__3_), .Y(_41_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_42_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_43_) );
NAND3X1 NAND3X1_6 ( .A(_41_), .B(_43_), .C(_42_), .Y(_44_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_38_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_39_) );
OAI21X1 OAI21X1_11 ( .A(_38_), .B(_39_), .C(_2__3_), .Y(_40_) );
NAND2X1 NAND2X1_8 ( .A(_40_), .B(_44_), .Y(_0__3_) );
OAI21X1 OAI21X1_12 ( .A(_41_), .B(_38_), .C(_43_), .Y(_1_) );
INVX1 INVX1_7 ( .A(w_cout_1_), .Y(_48_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_49_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_50_) );
NAND3X1 NAND3X1_7 ( .A(_48_), .B(_50_), .C(_49_), .Y(_51_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_45_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_46_) );
OAI21X1 OAI21X1_13 ( .A(_45_), .B(_46_), .C(w_cout_1_), .Y(_47_) );
NAND2X1 NAND2X1_10 ( .A(_47_), .B(_51_), .Y(_0__4_) );
OAI21X1 OAI21X1_14 ( .A(_48_), .B(_45_), .C(_50_), .Y(_4__1_) );
INVX1 INVX1_8 ( .A(_4__1_), .Y(_55_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_56_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_57_) );
NAND3X1 NAND3X1_8 ( .A(_55_), .B(_57_), .C(_56_), .Y(_58_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_52_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_53_) );
OAI21X1 OAI21X1_15 ( .A(_52_), .B(_53_), .C(_4__1_), .Y(_54_) );
NAND2X1 NAND2X1_12 ( .A(_54_), .B(_58_), .Y(_0__5_) );
OAI21X1 OAI21X1_16 ( .A(_55_), .B(_52_), .C(_57_), .Y(_4__2_) );
INVX1 INVX1_9 ( .A(_4__2_), .Y(_62_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_63_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_64_) );
NAND3X1 NAND3X1_9 ( .A(_62_), .B(_64_), .C(_63_), .Y(_65_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_59_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_60_) );
OAI21X1 OAI21X1_17 ( .A(_59_), .B(_60_), .C(_4__2_), .Y(_61_) );
NAND2X1 NAND2X1_14 ( .A(_61_), .B(_65_), .Y(_0__6_) );
OAI21X1 OAI21X1_18 ( .A(_62_), .B(_59_), .C(_64_), .Y(_4__3_) );
INVX1 INVX1_10 ( .A(_4__3_), .Y(_69_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_70_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_71_) );
NAND3X1 NAND3X1_10 ( .A(_69_), .B(_71_), .C(_70_), .Y(_72_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_66_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_67_) );
OAI21X1 OAI21X1_19 ( .A(_66_), .B(_67_), .C(_4__3_), .Y(_68_) );
NAND2X1 NAND2X1_16 ( .A(_68_), .B(_72_), .Y(_0__7_) );
OAI21X1 OAI21X1_20 ( .A(_69_), .B(_66_), .C(_71_), .Y(_3_) );
INVX1 INVX1_11 ( .A(cskip1_inst_cin), .Y(_76_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_77_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_78_) );
NAND3X1 NAND3X1_11 ( .A(_76_), .B(_78_), .C(_77_), .Y(_79_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_73_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_74_) );
OAI21X1 OAI21X1_21 ( .A(_73_), .B(_74_), .C(cskip1_inst_cin), .Y(_75_) );
NAND2X1 NAND2X1_18 ( .A(_75_), .B(_79_), .Y(cskip1_inst_sum) );
OAI21X1 OAI21X1_22 ( .A(_76_), .B(_73_), .C(_78_), .Y(cskip1_inst_rca0_w_CARRY_1_) );
INVX1 INVX1_12 ( .A(cskip1_inst_rca0_w_CARRY_1_), .Y(_81_) );
NAND2X1 NAND2X1_19 ( .A(gnd), .B(gnd), .Y(_82_) );
NOR2X1 NOR2X1_10 ( .A(gnd), .B(gnd), .Y(_80_) );
OAI21X1 OAI21X1_23 ( .A(_81_), .B(_80_), .C(_82_), .Y(cskip1_inst_rca0_w_CARRY_2_) );
INVX1 INVX1_13 ( .A(cskip1_inst_rca0_w_CARRY_2_), .Y(_84_) );
NAND2X1 NAND2X1_20 ( .A(gnd), .B(gnd), .Y(_85_) );
NOR2X1 NOR2X1_11 ( .A(gnd), .B(gnd), .Y(_83_) );
OAI21X1 OAI21X1_24 ( .A(_84_), .B(_83_), .C(_85_), .Y(cskip1_inst_rca0_w_CARRY_3_) );
INVX1 INVX1_14 ( .A(cskip1_inst_rca0_w_CARRY_3_), .Y(_87_) );
NAND2X1 NAND2X1_21 ( .A(gnd), .B(gnd), .Y(_88_) );
NOR2X1 NOR2X1_12 ( .A(gnd), .B(gnd), .Y(_86_) );
OAI21X1 OAI21X1_25 ( .A(_87_), .B(_86_), .C(_88_), .Y(cskip1_inst_cout0) );
INVX1 INVX1_15 ( .A(cskip1_inst_cout0), .Y(_89_) );
OAI21X1 OAI21X1_26 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .C(gnd), .Y(_90_) );
NAND2X1 NAND2X1_22 ( .A(_89_), .B(_90_), .Y(w_cout_3_) );
BUFX2 BUFX2_2 ( .A(w_cout_3_), .Y(cout) );
BUFX2 BUFX2_3 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_4 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_5 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_6 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_7 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_8 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_9 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_10 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_11 ( .A(cskip1_inst_sum), .Y(_0__8_) );
BUFX2 BUFX2_12 ( .A(gnd), .Y(_2__0_) );
BUFX2 BUFX2_13 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_14 ( .A(w_cout_1_), .Y(_4__0_) );
BUFX2 BUFX2_15 ( .A(_3_), .Y(_4__4_) );
BUFX2 BUFX2_16 ( .A(cskip1_inst_cin), .Y(cskip1_inst_rca0_w_CARRY_0_) );
BUFX2 BUFX2_17 ( .A(cskip1_inst_cout0), .Y(cskip1_inst_rca0_w_CARRY_4_) );
BUFX2 BUFX2_18 ( .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_19 ( .A(cskip1_inst_cin), .Y(w_cout_2_) );
endmodule
