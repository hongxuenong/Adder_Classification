module csa_20bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_4_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_25_) );
NAND2X1 NAND2X1_1 ( .A(_2_), .B(rca_inst_cout), .Y(_26_) );
OAI21X1 OAI21X1_1 ( .A(rca_inst_cout), .B(_25_), .C(_26_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3__0_), .Y(_27_) );
NAND2X1 NAND2X1_2 ( .A(_4__0_), .B(rca_inst_cout), .Y(_28_) );
OAI21X1 OAI21X1_2 ( .A(rca_inst_cout), .B(_27_), .C(_28_), .Y(_0__4_) );
INVX1 INVX1_3 ( .A(_3__1_), .Y(_29_) );
NAND2X1 NAND2X1_3 ( .A(rca_inst_cout), .B(_4__1_), .Y(_30_) );
OAI21X1 OAI21X1_3 ( .A(rca_inst_cout), .B(_29_), .C(_30_), .Y(_0__5_) );
INVX1 INVX1_4 ( .A(_3__2_), .Y(_31_) );
NAND2X1 NAND2X1_4 ( .A(rca_inst_cout), .B(_4__2_), .Y(_32_) );
OAI21X1 OAI21X1_4 ( .A(rca_inst_cout), .B(_31_), .C(_32_), .Y(_0__6_) );
INVX1 INVX1_5 ( .A(_3__3_), .Y(_33_) );
NAND2X1 NAND2X1_5 ( .A(rca_inst_cout), .B(_4__3_), .Y(_34_) );
OAI21X1 OAI21X1_5 ( .A(rca_inst_cout), .B(_33_), .C(_34_), .Y(_0__7_) );
INVX1 INVX1_6 ( .A(_7_), .Y(_35_) );
NAND2X1 NAND2X1_6 ( .A(_8_), .B(w_cout_1_), .Y(_36_) );
OAI21X1 OAI21X1_6 ( .A(w_cout_1_), .B(_35_), .C(_36_), .Y(w_cout_2_) );
INVX1 INVX1_7 ( .A(_9__0_), .Y(_37_) );
NAND2X1 NAND2X1_7 ( .A(_10__0_), .B(w_cout_1_), .Y(_38_) );
OAI21X1 OAI21X1_7 ( .A(w_cout_1_), .B(_37_), .C(_38_), .Y(_0__8_) );
INVX1 INVX1_8 ( .A(_9__1_), .Y(_39_) );
NAND2X1 NAND2X1_8 ( .A(w_cout_1_), .B(_10__1_), .Y(_40_) );
OAI21X1 OAI21X1_8 ( .A(w_cout_1_), .B(_39_), .C(_40_), .Y(_0__9_) );
INVX1 INVX1_9 ( .A(_9__2_), .Y(_41_) );
NAND2X1 NAND2X1_9 ( .A(w_cout_1_), .B(_10__2_), .Y(_42_) );
OAI21X1 OAI21X1_9 ( .A(w_cout_1_), .B(_41_), .C(_42_), .Y(_0__10_) );
INVX1 INVX1_10 ( .A(_9__3_), .Y(_43_) );
NAND2X1 NAND2X1_10 ( .A(w_cout_1_), .B(_10__3_), .Y(_44_) );
OAI21X1 OAI21X1_10 ( .A(w_cout_1_), .B(_43_), .C(_44_), .Y(_0__11_) );
INVX1 INVX1_11 ( .A(_13_), .Y(_45_) );
NAND2X1 NAND2X1_11 ( .A(_14_), .B(w_cout_2_), .Y(_46_) );
OAI21X1 OAI21X1_11 ( .A(w_cout_2_), .B(_45_), .C(_46_), .Y(w_cout_3_) );
INVX1 INVX1_12 ( .A(_15__0_), .Y(_47_) );
NAND2X1 NAND2X1_12 ( .A(_16__0_), .B(w_cout_2_), .Y(_48_) );
OAI21X1 OAI21X1_12 ( .A(w_cout_2_), .B(_47_), .C(_48_), .Y(_0__12_) );
INVX1 INVX1_13 ( .A(_15__1_), .Y(_49_) );
NAND2X1 NAND2X1_13 ( .A(w_cout_2_), .B(_16__1_), .Y(_50_) );
OAI21X1 OAI21X1_13 ( .A(w_cout_2_), .B(_49_), .C(_50_), .Y(_0__13_) );
INVX1 INVX1_14 ( .A(_15__2_), .Y(_51_) );
NAND2X1 NAND2X1_14 ( .A(w_cout_2_), .B(_16__2_), .Y(_52_) );
OAI21X1 OAI21X1_14 ( .A(w_cout_2_), .B(_51_), .C(_52_), .Y(_0__14_) );
INVX1 INVX1_15 ( .A(_15__3_), .Y(_53_) );
NAND2X1 NAND2X1_15 ( .A(w_cout_2_), .B(_16__3_), .Y(_54_) );
OAI21X1 OAI21X1_15 ( .A(w_cout_2_), .B(_53_), .C(_54_), .Y(_0__15_) );
INVX1 INVX1_16 ( .A(_19_), .Y(_55_) );
NAND2X1 NAND2X1_16 ( .A(_20_), .B(w_cout_3_), .Y(_56_) );
OAI21X1 OAI21X1_16 ( .A(w_cout_3_), .B(_55_), .C(_56_), .Y(w_cout_4_) );
INVX1 INVX1_17 ( .A(_21__0_), .Y(_57_) );
NAND2X1 NAND2X1_17 ( .A(_22__0_), .B(w_cout_3_), .Y(_58_) );
OAI21X1 OAI21X1_17 ( .A(w_cout_3_), .B(_57_), .C(_58_), .Y(_0__16_) );
INVX1 INVX1_18 ( .A(_21__1_), .Y(_59_) );
NAND2X1 NAND2X1_18 ( .A(w_cout_3_), .B(_22__1_), .Y(_60_) );
OAI21X1 OAI21X1_18 ( .A(w_cout_3_), .B(_59_), .C(_60_), .Y(_0__17_) );
INVX1 INVX1_19 ( .A(_21__2_), .Y(_61_) );
NAND2X1 NAND2X1_19 ( .A(w_cout_3_), .B(_22__2_), .Y(_62_) );
OAI21X1 OAI21X1_19 ( .A(w_cout_3_), .B(_61_), .C(_62_), .Y(_0__18_) );
INVX1 INVX1_20 ( .A(_21__3_), .Y(_63_) );
NAND2X1 NAND2X1_20 ( .A(w_cout_3_), .B(_22__3_), .Y(_64_) );
OAI21X1 OAI21X1_20 ( .A(w_cout_3_), .B(_63_), .C(_64_), .Y(_0__19_) );
INVX1 INVX1_21 ( .A(1'b0), .Y(_68_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_69_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_70_) );
NAND3X1 NAND3X1_1 ( .A(_68_), .B(_70_), .C(_69_), .Y(_71_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_65_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_66_) );
OAI21X1 OAI21X1_21 ( .A(_65_), .B(_66_), .C(1'b0), .Y(_67_) );
NAND2X1 NAND2X1_22 ( .A(_67_), .B(_71_), .Y(_3__0_) );
OAI21X1 OAI21X1_22 ( .A(_68_), .B(_65_), .C(_70_), .Y(_5__1_) );
INVX1 INVX1_22 ( .A(_5__1_), .Y(_75_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_76_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_77_) );
NAND3X1 NAND3X1_2 ( .A(_75_), .B(_77_), .C(_76_), .Y(_78_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_72_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_73_) );
OAI21X1 OAI21X1_23 ( .A(_72_), .B(_73_), .C(_5__1_), .Y(_74_) );
NAND2X1 NAND2X1_24 ( .A(_74_), .B(_78_), .Y(_3__1_) );
OAI21X1 OAI21X1_24 ( .A(_75_), .B(_72_), .C(_77_), .Y(_5__2_) );
INVX1 INVX1_23 ( .A(_5__2_), .Y(_82_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_83_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_84_) );
NAND3X1 NAND3X1_3 ( .A(_82_), .B(_84_), .C(_83_), .Y(_85_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_79_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_80_) );
OAI21X1 OAI21X1_25 ( .A(_79_), .B(_80_), .C(_5__2_), .Y(_81_) );
NAND2X1 NAND2X1_26 ( .A(_81_), .B(_85_), .Y(_3__2_) );
OAI21X1 OAI21X1_26 ( .A(_82_), .B(_79_), .C(_84_), .Y(_5__3_) );
INVX1 INVX1_24 ( .A(_5__3_), .Y(_89_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_90_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_91_) );
NAND3X1 NAND3X1_4 ( .A(_89_), .B(_91_), .C(_90_), .Y(_92_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_86_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_87_) );
OAI21X1 OAI21X1_27 ( .A(_86_), .B(_87_), .C(_5__3_), .Y(_88_) );
NAND2X1 NAND2X1_28 ( .A(_88_), .B(_92_), .Y(_3__3_) );
OAI21X1 OAI21X1_28 ( .A(_89_), .B(_86_), .C(_91_), .Y(_1_) );
INVX1 INVX1_25 ( .A(1'b1), .Y(_96_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_97_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_98_) );
NAND3X1 NAND3X1_5 ( .A(_96_), .B(_98_), .C(_97_), .Y(_99_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_93_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_94_) );
OAI21X1 OAI21X1_29 ( .A(_93_), .B(_94_), .C(1'b1), .Y(_95_) );
NAND2X1 NAND2X1_30 ( .A(_95_), .B(_99_), .Y(_4__0_) );
OAI21X1 OAI21X1_30 ( .A(_96_), .B(_93_), .C(_98_), .Y(_6__1_) );
INVX1 INVX1_26 ( .A(_6__1_), .Y(_103_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_104_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_105_) );
NAND3X1 NAND3X1_6 ( .A(_103_), .B(_105_), .C(_104_), .Y(_106_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_100_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_101_) );
OAI21X1 OAI21X1_31 ( .A(_100_), .B(_101_), .C(_6__1_), .Y(_102_) );
NAND2X1 NAND2X1_32 ( .A(_102_), .B(_106_), .Y(_4__1_) );
OAI21X1 OAI21X1_32 ( .A(_103_), .B(_100_), .C(_105_), .Y(_6__2_) );
INVX1 INVX1_27 ( .A(_6__2_), .Y(_110_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_111_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_112_) );
NAND3X1 NAND3X1_7 ( .A(_110_), .B(_112_), .C(_111_), .Y(_113_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_107_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_108_) );
OAI21X1 OAI21X1_33 ( .A(_107_), .B(_108_), .C(_6__2_), .Y(_109_) );
NAND2X1 NAND2X1_34 ( .A(_109_), .B(_113_), .Y(_4__2_) );
OAI21X1 OAI21X1_34 ( .A(_110_), .B(_107_), .C(_112_), .Y(_6__3_) );
INVX1 INVX1_28 ( .A(_6__3_), .Y(_117_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_118_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_119_) );
NAND3X1 NAND3X1_8 ( .A(_117_), .B(_119_), .C(_118_), .Y(_120_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_114_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_115_) );
OAI21X1 OAI21X1_35 ( .A(_114_), .B(_115_), .C(_6__3_), .Y(_116_) );
NAND2X1 NAND2X1_36 ( .A(_116_), .B(_120_), .Y(_4__3_) );
OAI21X1 OAI21X1_36 ( .A(_117_), .B(_114_), .C(_119_), .Y(_2_) );
INVX1 INVX1_29 ( .A(1'b0), .Y(_124_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_125_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_126_) );
NAND3X1 NAND3X1_9 ( .A(_124_), .B(_126_), .C(_125_), .Y(_127_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_121_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_122_) );
OAI21X1 OAI21X1_37 ( .A(_121_), .B(_122_), .C(1'b0), .Y(_123_) );
NAND2X1 NAND2X1_38 ( .A(_123_), .B(_127_), .Y(_9__0_) );
OAI21X1 OAI21X1_38 ( .A(_124_), .B(_121_), .C(_126_), .Y(_11__1_) );
INVX1 INVX1_30 ( .A(_11__1_), .Y(_131_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_132_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_133_) );
NAND3X1 NAND3X1_10 ( .A(_131_), .B(_133_), .C(_132_), .Y(_134_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_128_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_129_) );
OAI21X1 OAI21X1_39 ( .A(_128_), .B(_129_), .C(_11__1_), .Y(_130_) );
NAND2X1 NAND2X1_40 ( .A(_130_), .B(_134_), .Y(_9__1_) );
OAI21X1 OAI21X1_40 ( .A(_131_), .B(_128_), .C(_133_), .Y(_11__2_) );
INVX1 INVX1_31 ( .A(_11__2_), .Y(_138_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_139_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_140_) );
NAND3X1 NAND3X1_11 ( .A(_138_), .B(_140_), .C(_139_), .Y(_141_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_135_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_136_) );
OAI21X1 OAI21X1_41 ( .A(_135_), .B(_136_), .C(_11__2_), .Y(_137_) );
NAND2X1 NAND2X1_42 ( .A(_137_), .B(_141_), .Y(_9__2_) );
OAI21X1 OAI21X1_42 ( .A(_138_), .B(_135_), .C(_140_), .Y(_11__3_) );
INVX1 INVX1_32 ( .A(_11__3_), .Y(_145_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_146_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_147_) );
NAND3X1 NAND3X1_12 ( .A(_145_), .B(_147_), .C(_146_), .Y(_148_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_142_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_143_) );
OAI21X1 OAI21X1_43 ( .A(_142_), .B(_143_), .C(_11__3_), .Y(_144_) );
NAND2X1 NAND2X1_44 ( .A(_144_), .B(_148_), .Y(_9__3_) );
OAI21X1 OAI21X1_44 ( .A(_145_), .B(_142_), .C(_147_), .Y(_7_) );
INVX1 INVX1_33 ( .A(1'b1), .Y(_152_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_153_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_154_) );
NAND3X1 NAND3X1_13 ( .A(_152_), .B(_154_), .C(_153_), .Y(_155_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_149_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_150_) );
OAI21X1 OAI21X1_45 ( .A(_149_), .B(_150_), .C(1'b1), .Y(_151_) );
NAND2X1 NAND2X1_46 ( .A(_151_), .B(_155_), .Y(_10__0_) );
OAI21X1 OAI21X1_46 ( .A(_152_), .B(_149_), .C(_154_), .Y(_12__1_) );
INVX1 INVX1_34 ( .A(_12__1_), .Y(_159_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_160_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_161_) );
NAND3X1 NAND3X1_14 ( .A(_159_), .B(_161_), .C(_160_), .Y(_162_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_156_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_157_) );
OAI21X1 OAI21X1_47 ( .A(_156_), .B(_157_), .C(_12__1_), .Y(_158_) );
NAND2X1 NAND2X1_48 ( .A(_158_), .B(_162_), .Y(_10__1_) );
OAI21X1 OAI21X1_48 ( .A(_159_), .B(_156_), .C(_161_), .Y(_12__2_) );
INVX1 INVX1_35 ( .A(_12__2_), .Y(_166_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_167_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_168_) );
NAND3X1 NAND3X1_15 ( .A(_166_), .B(_168_), .C(_167_), .Y(_169_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_163_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_164_) );
OAI21X1 OAI21X1_49 ( .A(_163_), .B(_164_), .C(_12__2_), .Y(_165_) );
NAND2X1 NAND2X1_50 ( .A(_165_), .B(_169_), .Y(_10__2_) );
OAI21X1 OAI21X1_50 ( .A(_166_), .B(_163_), .C(_168_), .Y(_12__3_) );
INVX1 INVX1_36 ( .A(_12__3_), .Y(_173_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_174_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_175_) );
NAND3X1 NAND3X1_16 ( .A(_173_), .B(_175_), .C(_174_), .Y(_176_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_170_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_171_) );
OAI21X1 OAI21X1_51 ( .A(_170_), .B(_171_), .C(_12__3_), .Y(_172_) );
NAND2X1 NAND2X1_52 ( .A(_172_), .B(_176_), .Y(_10__3_) );
OAI21X1 OAI21X1_52 ( .A(_173_), .B(_170_), .C(_175_), .Y(_8_) );
INVX1 INVX1_37 ( .A(1'b0), .Y(_180_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_181_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_182_) );
NAND3X1 NAND3X1_17 ( .A(_180_), .B(_182_), .C(_181_), .Y(_183_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_177_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_178_) );
OAI21X1 OAI21X1_53 ( .A(_177_), .B(_178_), .C(1'b0), .Y(_179_) );
NAND2X1 NAND2X1_54 ( .A(_179_), .B(_183_), .Y(_15__0_) );
OAI21X1 OAI21X1_54 ( .A(_180_), .B(_177_), .C(_182_), .Y(_17__1_) );
INVX1 INVX1_38 ( .A(_17__1_), .Y(_187_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_188_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_189_) );
NAND3X1 NAND3X1_18 ( .A(_187_), .B(_189_), .C(_188_), .Y(_190_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_184_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_185_) );
OAI21X1 OAI21X1_55 ( .A(_184_), .B(_185_), .C(_17__1_), .Y(_186_) );
NAND2X1 NAND2X1_56 ( .A(_186_), .B(_190_), .Y(_15__1_) );
OAI21X1 OAI21X1_56 ( .A(_187_), .B(_184_), .C(_189_), .Y(_17__2_) );
INVX1 INVX1_39 ( .A(_17__2_), .Y(_194_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_195_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_196_) );
NAND3X1 NAND3X1_19 ( .A(_194_), .B(_196_), .C(_195_), .Y(_197_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_191_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_192_) );
OAI21X1 OAI21X1_57 ( .A(_191_), .B(_192_), .C(_17__2_), .Y(_193_) );
NAND2X1 NAND2X1_58 ( .A(_193_), .B(_197_), .Y(_15__2_) );
OAI21X1 OAI21X1_58 ( .A(_194_), .B(_191_), .C(_196_), .Y(_17__3_) );
INVX1 INVX1_40 ( .A(_17__3_), .Y(_201_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_202_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_203_) );
NAND3X1 NAND3X1_20 ( .A(_201_), .B(_203_), .C(_202_), .Y(_204_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_198_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_199_) );
OAI21X1 OAI21X1_59 ( .A(_198_), .B(_199_), .C(_17__3_), .Y(_200_) );
NAND2X1 NAND2X1_60 ( .A(_200_), .B(_204_), .Y(_15__3_) );
OAI21X1 OAI21X1_60 ( .A(_201_), .B(_198_), .C(_203_), .Y(_13_) );
INVX1 INVX1_41 ( .A(1'b1), .Y(_208_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_209_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_210_) );
NAND3X1 NAND3X1_21 ( .A(_208_), .B(_210_), .C(_209_), .Y(_211_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_205_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_206_) );
OAI21X1 OAI21X1_61 ( .A(_205_), .B(_206_), .C(1'b1), .Y(_207_) );
NAND2X1 NAND2X1_62 ( .A(_207_), .B(_211_), .Y(_16__0_) );
OAI21X1 OAI21X1_62 ( .A(_208_), .B(_205_), .C(_210_), .Y(_18__1_) );
INVX1 INVX1_42 ( .A(_18__1_), .Y(_215_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_216_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_217_) );
NAND3X1 NAND3X1_22 ( .A(_215_), .B(_217_), .C(_216_), .Y(_218_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_212_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_213_) );
OAI21X1 OAI21X1_63 ( .A(_212_), .B(_213_), .C(_18__1_), .Y(_214_) );
NAND2X1 NAND2X1_64 ( .A(_214_), .B(_218_), .Y(_16__1_) );
OAI21X1 OAI21X1_64 ( .A(_215_), .B(_212_), .C(_217_), .Y(_18__2_) );
INVX1 INVX1_43 ( .A(_18__2_), .Y(_222_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_223_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_224_) );
NAND3X1 NAND3X1_23 ( .A(_222_), .B(_224_), .C(_223_), .Y(_225_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_219_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_220_) );
OAI21X1 OAI21X1_65 ( .A(_219_), .B(_220_), .C(_18__2_), .Y(_221_) );
NAND2X1 NAND2X1_66 ( .A(_221_), .B(_225_), .Y(_16__2_) );
OAI21X1 OAI21X1_66 ( .A(_222_), .B(_219_), .C(_224_), .Y(_18__3_) );
INVX1 INVX1_44 ( .A(_18__3_), .Y(_229_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_230_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_231_) );
NAND3X1 NAND3X1_24 ( .A(_229_), .B(_231_), .C(_230_), .Y(_232_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_226_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_227_) );
OAI21X1 OAI21X1_67 ( .A(_226_), .B(_227_), .C(_18__3_), .Y(_228_) );
NAND2X1 NAND2X1_68 ( .A(_228_), .B(_232_), .Y(_16__3_) );
OAI21X1 OAI21X1_68 ( .A(_229_), .B(_226_), .C(_231_), .Y(_14_) );
INVX1 INVX1_45 ( .A(1'b0), .Y(_236_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_237_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_238_) );
NAND3X1 NAND3X1_25 ( .A(_236_), .B(_238_), .C(_237_), .Y(_239_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_233_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_234_) );
OAI21X1 OAI21X1_69 ( .A(_233_), .B(_234_), .C(1'b0), .Y(_235_) );
NAND2X1 NAND2X1_70 ( .A(_235_), .B(_239_), .Y(_21__0_) );
OAI21X1 OAI21X1_70 ( .A(_236_), .B(_233_), .C(_238_), .Y(_23__1_) );
INVX1 INVX1_46 ( .A(_23__1_), .Y(_243_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_244_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_245_) );
NAND3X1 NAND3X1_26 ( .A(_243_), .B(_245_), .C(_244_), .Y(_246_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_240_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_241_) );
OAI21X1 OAI21X1_71 ( .A(_240_), .B(_241_), .C(_23__1_), .Y(_242_) );
NAND2X1 NAND2X1_72 ( .A(_242_), .B(_246_), .Y(_21__1_) );
OAI21X1 OAI21X1_72 ( .A(_243_), .B(_240_), .C(_245_), .Y(_23__2_) );
INVX1 INVX1_47 ( .A(_23__2_), .Y(_250_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_251_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_252_) );
NAND3X1 NAND3X1_27 ( .A(_250_), .B(_252_), .C(_251_), .Y(_253_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_247_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_248_) );
OAI21X1 OAI21X1_73 ( .A(_247_), .B(_248_), .C(_23__2_), .Y(_249_) );
NAND2X1 NAND2X1_74 ( .A(_249_), .B(_253_), .Y(_21__2_) );
OAI21X1 OAI21X1_74 ( .A(_250_), .B(_247_), .C(_252_), .Y(_23__3_) );
INVX1 INVX1_48 ( .A(_23__3_), .Y(_257_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_258_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_259_) );
NAND3X1 NAND3X1_28 ( .A(_257_), .B(_259_), .C(_258_), .Y(_260_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_254_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_255_) );
OAI21X1 OAI21X1_75 ( .A(_254_), .B(_255_), .C(_23__3_), .Y(_256_) );
NAND2X1 NAND2X1_76 ( .A(_256_), .B(_260_), .Y(_21__3_) );
OAI21X1 OAI21X1_76 ( .A(_257_), .B(_254_), .C(_259_), .Y(_19_) );
INVX1 INVX1_49 ( .A(1'b1), .Y(_264_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_265_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_266_) );
NAND3X1 NAND3X1_29 ( .A(_264_), .B(_266_), .C(_265_), .Y(_267_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_261_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_262_) );
OAI21X1 OAI21X1_77 ( .A(_261_), .B(_262_), .C(1'b1), .Y(_263_) );
NAND2X1 NAND2X1_78 ( .A(_263_), .B(_267_), .Y(_22__0_) );
OAI21X1 OAI21X1_78 ( .A(_264_), .B(_261_), .C(_266_), .Y(_24__1_) );
INVX1 INVX1_50 ( .A(_24__1_), .Y(_271_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_272_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_273_) );
NAND3X1 NAND3X1_30 ( .A(_271_), .B(_273_), .C(_272_), .Y(_274_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_268_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_269_) );
OAI21X1 OAI21X1_79 ( .A(_268_), .B(_269_), .C(_24__1_), .Y(_270_) );
NAND2X1 NAND2X1_80 ( .A(_270_), .B(_274_), .Y(_22__1_) );
OAI21X1 OAI21X1_80 ( .A(_271_), .B(_268_), .C(_273_), .Y(_24__2_) );
INVX1 INVX1_51 ( .A(_24__2_), .Y(_278_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_279_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_280_) );
NAND3X1 NAND3X1_31 ( .A(_278_), .B(_280_), .C(_279_), .Y(_281_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_275_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_276_) );
OAI21X1 OAI21X1_81 ( .A(_275_), .B(_276_), .C(_24__2_), .Y(_277_) );
NAND2X1 NAND2X1_82 ( .A(_277_), .B(_281_), .Y(_22__2_) );
OAI21X1 OAI21X1_82 ( .A(_278_), .B(_275_), .C(_280_), .Y(_24__3_) );
INVX1 INVX1_52 ( .A(_24__3_), .Y(_285_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_286_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_287_) );
NAND3X1 NAND3X1_32 ( .A(_285_), .B(_287_), .C(_286_), .Y(_288_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_282_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_283_) );
OAI21X1 OAI21X1_83 ( .A(_282_), .B(_283_), .C(_24__3_), .Y(_284_) );
NAND2X1 NAND2X1_84 ( .A(_284_), .B(_288_), .Y(_22__3_) );
OAI21X1 OAI21X1_84 ( .A(_285_), .B(_282_), .C(_287_), .Y(_20_) );
INVX1 INVX1_53 ( .A(1'b0), .Y(_292_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_293_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_294_) );
NAND3X1 NAND3X1_33 ( .A(_292_), .B(_294_), .C(_293_), .Y(_295_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_289_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_290_) );
OAI21X1 OAI21X1_85 ( .A(_289_), .B(_290_), .C(1'b0), .Y(_291_) );
NAND2X1 NAND2X1_86 ( .A(_291_), .B(_295_), .Y(_0__0_) );
OAI21X1 OAI21X1_86 ( .A(_292_), .B(_289_), .C(_294_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_54 ( .A(rca_inst_w_CARRY_1_), .Y(_299_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_300_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_301_) );
NAND3X1 NAND3X1_34 ( .A(_299_), .B(_301_), .C(_300_), .Y(_302_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_296_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_297_) );
OAI21X1 OAI21X1_87 ( .A(_296_), .B(_297_), .C(rca_inst_w_CARRY_1_), .Y(_298_) );
NAND2X1 NAND2X1_88 ( .A(_298_), .B(_302_), .Y(_0__1_) );
OAI21X1 OAI21X1_88 ( .A(_299_), .B(_296_), .C(_301_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_55 ( .A(rca_inst_w_CARRY_2_), .Y(_306_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_307_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_308_) );
NAND3X1 NAND3X1_35 ( .A(_306_), .B(_308_), .C(_307_), .Y(_309_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_303_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_304_) );
OAI21X1 OAI21X1_89 ( .A(_303_), .B(_304_), .C(rca_inst_w_CARRY_2_), .Y(_305_) );
NAND2X1 NAND2X1_90 ( .A(_305_), .B(_309_), .Y(_0__2_) );
OAI21X1 OAI21X1_90 ( .A(_306_), .B(_303_), .C(_308_), .Y(rca_inst_w_CARRY_3_) );
INVX1 INVX1_56 ( .A(rca_inst_w_CARRY_3_), .Y(_313_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_314_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_315_) );
NAND3X1 NAND3X1_36 ( .A(_313_), .B(_315_), .C(_314_), .Y(_316_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_310_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_311_) );
OAI21X1 OAI21X1_91 ( .A(_310_), .B(_311_), .C(rca_inst_w_CARRY_3_), .Y(_312_) );
NAND2X1 NAND2X1_92 ( .A(_312_), .B(_316_), .Y(_0__3_) );
OAI21X1 OAI21X1_92 ( .A(_313_), .B(_310_), .C(_315_), .Y(rca_inst_cout) );
BUFX2 BUFX2_22 ( .A(1'b0), .Y(_5__0_) );
BUFX2 BUFX2_23 ( .A(_1_), .Y(_5__4_) );
BUFX2 BUFX2_24 ( .A(1'b1), .Y(_6__0_) );
BUFX2 BUFX2_25 ( .A(_2_), .Y(_6__4_) );
BUFX2 BUFX2_26 ( .A(1'b0), .Y(_11__0_) );
BUFX2 BUFX2_27 ( .A(_7_), .Y(_11__4_) );
BUFX2 BUFX2_28 ( .A(1'b1), .Y(_12__0_) );
BUFX2 BUFX2_29 ( .A(_8_), .Y(_12__4_) );
BUFX2 BUFX2_30 ( .A(1'b0), .Y(_17__0_) );
BUFX2 BUFX2_31 ( .A(_13_), .Y(_17__4_) );
BUFX2 BUFX2_32 ( .A(1'b1), .Y(_18__0_) );
BUFX2 BUFX2_33 ( .A(_14_), .Y(_18__4_) );
BUFX2 BUFX2_34 ( .A(1'b0), .Y(_23__0_) );
BUFX2 BUFX2_35 ( .A(_19_), .Y(_23__4_) );
BUFX2 BUFX2_36 ( .A(1'b1), .Y(_24__0_) );
BUFX2 BUFX2_37 ( .A(_20_), .Y(_24__4_) );
BUFX2 BUFX2_38 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_39 ( .A(rca_inst_cout), .Y(rca_inst_w_CARRY_4_) );
BUFX2 BUFX2_40 ( .A(rca_inst_cout), .Y(w_cout_0_) );
endmodule
