module csa_11bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output cout;

BUFX2 BUFX2_1 ( .A(_0_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_1__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_1__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_1__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_1__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_1__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_1__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_1__10_), .Y(sum[10]) );
INVX1 INVX1_1 ( .A(_2_), .Y(_8_) );
NAND2X1 NAND2X1_1 ( .A(_3_), .B(rca_inst_cout), .Y(_9_) );
OAI21X1 OAI21X1_1 ( .A(rca_inst_cout), .B(_8_), .C(_9_), .Y(csa_inst_cin) );
INVX1 INVX1_2 ( .A(_4__0_), .Y(_10_) );
NAND2X1 NAND2X1_2 ( .A(_5__0_), .B(rca_inst_cout), .Y(_11_) );
OAI21X1 OAI21X1_2 ( .A(rca_inst_cout), .B(_10_), .C(_11_), .Y(_1__4_) );
INVX1 INVX1_3 ( .A(_4__1_), .Y(_12_) );
NAND2X1 NAND2X1_3 ( .A(rca_inst_cout), .B(_5__1_), .Y(_13_) );
OAI21X1 OAI21X1_3 ( .A(rca_inst_cout), .B(_12_), .C(_13_), .Y(_1__5_) );
INVX1 INVX1_4 ( .A(_4__2_), .Y(_14_) );
NAND2X1 NAND2X1_4 ( .A(rca_inst_cout), .B(_5__2_), .Y(_15_) );
OAI21X1 OAI21X1_4 ( .A(rca_inst_cout), .B(_14_), .C(_15_), .Y(_1__6_) );
INVX1 INVX1_5 ( .A(_4__3_), .Y(_16_) );
NAND2X1 NAND2X1_5 ( .A(rca_inst_cout), .B(_5__3_), .Y(_17_) );
OAI21X1 OAI21X1_5 ( .A(rca_inst_cout), .B(_16_), .C(_17_), .Y(_1__7_) );
INVX1 INVX1_6 ( .A(1'b0), .Y(_21_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_22_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_23_) );
NAND3X1 NAND3X1_1 ( .A(_21_), .B(_23_), .C(_22_), .Y(_24_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_18_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_19_) );
OAI21X1 OAI21X1_6 ( .A(_18_), .B(_19_), .C(1'b0), .Y(_20_) );
NAND2X1 NAND2X1_7 ( .A(_20_), .B(_24_), .Y(_4__0_) );
OAI21X1 OAI21X1_7 ( .A(_21_), .B(_18_), .C(_23_), .Y(_6__1_) );
INVX1 INVX1_7 ( .A(_6__3_), .Y(_28_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_29_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_30_) );
NAND3X1 NAND3X1_2 ( .A(_28_), .B(_30_), .C(_29_), .Y(_31_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_25_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_26_) );
OAI21X1 OAI21X1_8 ( .A(_25_), .B(_26_), .C(_6__3_), .Y(_27_) );
NAND2X1 NAND2X1_9 ( .A(_27_), .B(_31_), .Y(_4__3_) );
OAI21X1 OAI21X1_9 ( .A(_28_), .B(_25_), .C(_30_), .Y(_2_) );
INVX1 INVX1_8 ( .A(_6__1_), .Y(_35_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_36_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_37_) );
NAND3X1 NAND3X1_3 ( .A(_35_), .B(_37_), .C(_36_), .Y(_38_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_32_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_33_) );
OAI21X1 OAI21X1_10 ( .A(_32_), .B(_33_), .C(_6__1_), .Y(_34_) );
NAND2X1 NAND2X1_11 ( .A(_34_), .B(_38_), .Y(_4__1_) );
OAI21X1 OAI21X1_11 ( .A(_35_), .B(_32_), .C(_37_), .Y(_6__2_) );
INVX1 INVX1_9 ( .A(_6__2_), .Y(_42_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_43_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_44_) );
NAND3X1 NAND3X1_4 ( .A(_42_), .B(_44_), .C(_43_), .Y(_45_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_39_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_40_) );
OAI21X1 OAI21X1_12 ( .A(_39_), .B(_40_), .C(_6__2_), .Y(_41_) );
NAND2X1 NAND2X1_13 ( .A(_41_), .B(_45_), .Y(_4__2_) );
OAI21X1 OAI21X1_13 ( .A(_42_), .B(_39_), .C(_44_), .Y(_6__3_) );
INVX1 INVX1_10 ( .A(1'b1), .Y(_49_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_50_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_51_) );
NAND3X1 NAND3X1_5 ( .A(_49_), .B(_51_), .C(_50_), .Y(_52_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_46_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_47_) );
OAI21X1 OAI21X1_14 ( .A(_46_), .B(_47_), .C(1'b1), .Y(_48_) );
NAND2X1 NAND2X1_15 ( .A(_48_), .B(_52_), .Y(_5__0_) );
OAI21X1 OAI21X1_15 ( .A(_49_), .B(_46_), .C(_51_), .Y(_7__1_) );
INVX1 INVX1_11 ( .A(_7__3_), .Y(_56_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_57_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_58_) );
NAND3X1 NAND3X1_6 ( .A(_56_), .B(_58_), .C(_57_), .Y(_59_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_53_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_54_) );
OAI21X1 OAI21X1_16 ( .A(_53_), .B(_54_), .C(_7__3_), .Y(_55_) );
NAND2X1 NAND2X1_17 ( .A(_55_), .B(_59_), .Y(_5__3_) );
OAI21X1 OAI21X1_17 ( .A(_56_), .B(_53_), .C(_58_), .Y(_3_) );
INVX1 INVX1_12 ( .A(_7__1_), .Y(_63_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_64_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_65_) );
NAND3X1 NAND3X1_7 ( .A(_63_), .B(_65_), .C(_64_), .Y(_66_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_60_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_61_) );
OAI21X1 OAI21X1_18 ( .A(_60_), .B(_61_), .C(_7__1_), .Y(_62_) );
NAND2X1 NAND2X1_19 ( .A(_62_), .B(_66_), .Y(_5__1_) );
OAI21X1 OAI21X1_19 ( .A(_63_), .B(_60_), .C(_65_), .Y(_7__2_) );
INVX1 INVX1_13 ( .A(_7__2_), .Y(_70_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_71_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_72_) );
NAND3X1 NAND3X1_8 ( .A(_70_), .B(_72_), .C(_71_), .Y(_73_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_67_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_68_) );
OAI21X1 OAI21X1_20 ( .A(_67_), .B(_68_), .C(_7__2_), .Y(_69_) );
NAND2X1 NAND2X1_21 ( .A(_69_), .B(_73_), .Y(_5__2_) );
OAI21X1 OAI21X1_21 ( .A(_70_), .B(_67_), .C(_72_), .Y(_7__3_) );
INVX1 INVX1_14 ( .A(csa_inst_cout0_0), .Y(_74_) );
NAND2X1 NAND2X1_22 ( .A(csa_inst_cout0_1), .B(csa_inst_cin), .Y(_75_) );
OAI21X1 OAI21X1_22 ( .A(csa_inst_cin), .B(_74_), .C(_75_), .Y(_0_) );
INVX1 INVX1_15 ( .A(csa_inst_rca0_0_fa0_o_sum), .Y(_76_) );
NAND2X1 NAND2X1_23 ( .A(csa_inst_rca0_1_fa0_o_sum), .B(csa_inst_cin), .Y(_77_) );
OAI21X1 OAI21X1_23 ( .A(csa_inst_cin), .B(_76_), .C(_77_), .Y(_1__8_) );
INVX1 INVX1_16 ( .A(csa_inst_rca0_0_fa1_o_sum), .Y(_78_) );
NAND2X1 NAND2X1_24 ( .A(csa_inst_cin), .B(csa_inst_rca0_1_fa1_o_sum), .Y(_79_) );
OAI21X1 OAI21X1_24 ( .A(csa_inst_cin), .B(_78_), .C(_79_), .Y(_1__9_) );
INVX1 INVX1_17 ( .A(csa_inst_rca0_0_fa2_o_sum), .Y(_80_) );
NAND2X1 NAND2X1_25 ( .A(csa_inst_cin), .B(csa_inst_rca0_1_fa2_o_sum), .Y(_81_) );
OAI21X1 OAI21X1_25 ( .A(csa_inst_cin), .B(_80_), .C(_81_), .Y(_1__10_) );
INVX1 INVX1_18 ( .A(1'b0), .Y(_85_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_86_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_87_) );
NAND3X1 NAND3X1_9 ( .A(_85_), .B(_87_), .C(_86_), .Y(_88_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_82_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_83_) );
OAI21X1 OAI21X1_26 ( .A(_82_), .B(_83_), .C(1'b0), .Y(_84_) );
NAND2X1 NAND2X1_27 ( .A(_84_), .B(_88_), .Y(csa_inst_rca0_0_fa0_o_sum) );
OAI21X1 OAI21X1_27 ( .A(_85_), .B(_82_), .C(_87_), .Y(csa_inst_rca0_0_fa0_o_carry) );
INVX1 INVX1_19 ( .A(csa_inst_rca0_0_fa0_o_carry), .Y(_92_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_93_) );
NAND2X1 NAND2X1_28 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_94_) );
NAND3X1 NAND3X1_10 ( .A(_92_), .B(_94_), .C(_93_), .Y(_95_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_89_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_90_) );
OAI21X1 OAI21X1_28 ( .A(_89_), .B(_90_), .C(csa_inst_rca0_0_fa0_o_carry), .Y(_91_) );
NAND2X1 NAND2X1_29 ( .A(_91_), .B(_95_), .Y(csa_inst_rca0_0_fa1_o_sum) );
OAI21X1 OAI21X1_29 ( .A(_92_), .B(_89_), .C(_94_), .Y(csa_inst_rca0_0_fa1_o_carry) );
INVX1 INVX1_20 ( .A(csa_inst_rca0_0_fa1_o_carry), .Y(_99_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_100_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_101_) );
NAND3X1 NAND3X1_11 ( .A(_99_), .B(_101_), .C(_100_), .Y(_102_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_96_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_97_) );
OAI21X1 OAI21X1_30 ( .A(_96_), .B(_97_), .C(csa_inst_rca0_0_fa1_o_carry), .Y(_98_) );
NAND2X1 NAND2X1_31 ( .A(_98_), .B(_102_), .Y(csa_inst_rca0_0_fa2_o_sum) );
OAI21X1 OAI21X1_31 ( .A(_99_), .B(_96_), .C(_101_), .Y(csa_inst_cout0_0) );
INVX1 INVX1_21 ( .A(1'b1), .Y(_106_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_107_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_108_) );
NAND3X1 NAND3X1_12 ( .A(_106_), .B(_108_), .C(_107_), .Y(_109_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_103_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_104_) );
OAI21X1 OAI21X1_32 ( .A(_103_), .B(_104_), .C(1'b1), .Y(_105_) );
NAND2X1 NAND2X1_33 ( .A(_105_), .B(_109_), .Y(csa_inst_rca0_1_fa0_o_sum) );
OAI21X1 OAI21X1_33 ( .A(_106_), .B(_103_), .C(_108_), .Y(csa_inst_rca0_1_fa0_o_carry) );
INVX1 INVX1_22 ( .A(csa_inst_rca0_1_fa0_o_carry), .Y(_113_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_114_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_115_) );
NAND3X1 NAND3X1_13 ( .A(_113_), .B(_115_), .C(_114_), .Y(_116_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_110_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_111_) );
OAI21X1 OAI21X1_34 ( .A(_110_), .B(_111_), .C(csa_inst_rca0_1_fa0_o_carry), .Y(_112_) );
NAND2X1 NAND2X1_35 ( .A(_112_), .B(_116_), .Y(csa_inst_rca0_1_fa1_o_sum) );
OAI21X1 OAI21X1_35 ( .A(_113_), .B(_110_), .C(_115_), .Y(csa_inst_rca0_1_fa1_o_carry) );
INVX1 INVX1_23 ( .A(csa_inst_rca0_1_fa1_o_carry), .Y(_120_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_121_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_122_) );
NAND3X1 NAND3X1_14 ( .A(_120_), .B(_122_), .C(_121_), .Y(_123_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_117_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_118_) );
OAI21X1 OAI21X1_36 ( .A(_117_), .B(_118_), .C(csa_inst_rca0_1_fa1_o_carry), .Y(_119_) );
NAND2X1 NAND2X1_37 ( .A(_119_), .B(_123_), .Y(csa_inst_rca0_1_fa2_o_sum) );
OAI21X1 OAI21X1_37 ( .A(_120_), .B(_117_), .C(_122_), .Y(csa_inst_cout0_1) );
INVX1 INVX1_24 ( .A(1'b0), .Y(_127_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_128_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_129_) );
NAND3X1 NAND3X1_15 ( .A(_127_), .B(_129_), .C(_128_), .Y(_130_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_124_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_125_) );
OAI21X1 OAI21X1_38 ( .A(_124_), .B(_125_), .C(1'b0), .Y(_126_) );
NAND2X1 NAND2X1_39 ( .A(_126_), .B(_130_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_39 ( .A(_127_), .B(_124_), .C(_129_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_25 ( .A(rca_inst_fa3_i_carry), .Y(_134_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_135_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_136_) );
NAND3X1 NAND3X1_16 ( .A(_134_), .B(_136_), .C(_135_), .Y(_137_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_131_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_132_) );
OAI21X1 OAI21X1_40 ( .A(_131_), .B(_132_), .C(rca_inst_fa3_i_carry), .Y(_133_) );
NAND2X1 NAND2X1_41 ( .A(_133_), .B(_137_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_41 ( .A(_134_), .B(_131_), .C(_136_), .Y(rca_inst_cout) );
INVX1 INVX1_26 ( .A(rca_inst_fa0_o_carry), .Y(_141_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_142_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_143_) );
NAND3X1 NAND3X1_17 ( .A(_141_), .B(_143_), .C(_142_), .Y(_144_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_138_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_139_) );
OAI21X1 OAI21X1_42 ( .A(_138_), .B(_139_), .C(rca_inst_fa0_o_carry), .Y(_140_) );
NAND2X1 NAND2X1_43 ( .A(_140_), .B(_144_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_43 ( .A(_141_), .B(_138_), .C(_143_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_27 ( .A(rca_inst_fa_1__o_carry), .Y(_148_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_149_) );
NAND2X1 NAND2X1_44 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_150_) );
NAND3X1 NAND3X1_18 ( .A(_148_), .B(_150_), .C(_149_), .Y(_151_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_145_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_146_) );
OAI21X1 OAI21X1_44 ( .A(_145_), .B(_146_), .C(rca_inst_fa_1__o_carry), .Y(_147_) );
NAND2X1 NAND2X1_45 ( .A(_147_), .B(_151_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_45 ( .A(_148_), .B(_145_), .C(_150_), .Y(rca_inst_fa3_i_carry) );
BUFX2 BUFX2_13 ( .A(rca_inst_fa0_o_sum), .Y(_1__0_) );
BUFX2 BUFX2_14 ( .A(rca_inst_fa_1__o_sum), .Y(_1__1_) );
BUFX2 BUFX2_15 ( .A(rca_inst_fa_2__o_sum), .Y(_1__2_) );
BUFX2 BUFX2_16 ( .A(rca_inst_fa3_o_sum), .Y(_1__3_) );
endmodule
