module CSkipA_29bit ( gnd, vdd, i_add_term1, i_add_term2, sum, cout);

input gnd, vdd;
output cout;
input [28:0] i_add_term1;
input [28:0] i_add_term2;
output [28:0] sum;

BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .Y(cout) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_sum), .Y(sum[28]) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .Y(_22_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(_22_), .Y(_23_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .Y(_24_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .B(_24_), .Y(_25_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .Y(_26_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(_26_), .Y(_27_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .Y(_28_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .B(_28_), .Y(_29_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_25_), .C(_27_), .D(_29_), .Y(_30_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_31_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_32_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_32_), .Y(_33_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_34_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_34_), .Y(_35_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_35_), .Y(_3_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_36_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_3_), .Y(_37_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_36_), .C(_37_), .Y(w_cout_1_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[4]), .Y(_38_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(_38_), .Y(_39_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .Y(_40_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[4]), .B(_40_), .Y(_41_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[5]), .Y(_42_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(_42_), .Y(_43_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .Y(_44_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[5]), .B(_44_), .Y(_45_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_41_), .C(_43_), .D(_45_), .Y(_46_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_47_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_48_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_48_), .Y(_49_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_50_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_50_), .Y(_51_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_51_), .Y(_6_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(_52_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_6_), .Y(_53_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_52_), .C(_53_), .Y(w_cout_2_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[8]), .Y(_54_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(_54_), .Y(_55_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .Y(_56_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[8]), .B(_56_), .Y(_57_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[9]), .Y(_58_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(_58_), .Y(_59_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .Y(_60_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[9]), .B(_60_), .Y(_61_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_57_), .C(_59_), .D(_61_), .Y(_62_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_63_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_64_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_64_), .Y(_65_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_66_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_66_), .Y(_67_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_67_), .Y(_9_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_68_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_9_), .Y(_69_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_68_), .C(_69_), .Y(w_cout_3_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[12]), .Y(_70_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(_70_), .Y(_71_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .Y(_72_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[12]), .B(_72_), .Y(_73_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[13]), .Y(_74_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(_74_), .Y(_75_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .Y(_76_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[13]), .B(_76_), .Y(_77_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_73_), .C(_75_), .D(_77_), .Y(_78_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_79_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_80_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_80_), .Y(_81_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_82_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_82_), .Y(_83_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_83_), .Y(_12_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(_84_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_12_), .Y(_85_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_84_), .C(_85_), .Y(w_cout_4_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[16]), .Y(_86_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(_86_), .Y(_87_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .Y(_88_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[16]), .B(_88_), .Y(_89_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[17]), .Y(_90_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(_90_), .Y(_91_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .Y(_92_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[17]), .B(_92_), .Y(_93_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_89_), .C(_91_), .D(_93_), .Y(_94_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_95_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_96_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_96_), .Y(_97_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_98_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_98_), .Y(_99_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_99_), .Y(_15_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_100_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_15_), .Y(_101_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_100_), .C(_101_), .Y(w_cout_5_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[20]), .Y(_102_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(_102_), .Y(_103_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .Y(_104_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[20]), .B(_104_), .Y(_105_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[21]), .Y(_106_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(_106_), .Y(_107_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .Y(_108_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[21]), .B(_108_), .Y(_109_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_105_), .C(_107_), .D(_109_), .Y(_110_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_111_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_112_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_112_), .Y(_113_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_114_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_114_), .Y(_115_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_115_), .Y(_18_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_116_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_18_), .Y(_117_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_116_), .C(_117_), .Y(w_cout_6_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[24]), .Y(_118_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(_118_), .Y(_119_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .Y(_120_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[24]), .B(_120_), .Y(_121_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[25]), .Y(_122_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(_122_), .Y(_123_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .Y(_124_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[25]), .B(_124_), .Y(_125_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_121_), .C(_123_), .D(_125_), .Y(_126_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_127_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_128_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_128_), .Y(_129_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_130_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_129_), .B(_130_), .Y(_131_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_131_), .Y(_21_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_132_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_21_), .Y(_133_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_132_), .C(_133_), .Y(cskip1_inst_cin) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_137_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_138_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_139_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(_139_), .C(_138_), .Y(_140_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_134_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_135_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_135_), .C(gnd), .Y(_136_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_140_), .Y(_0__0_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(_134_), .C(_139_), .Y(_2__1_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_2__1_), .Y(_144_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_145_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_146_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_146_), .C(_145_), .Y(_147_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_141_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_142_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_142_), .C(_2__1_), .Y(_143_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_147_), .Y(_0__1_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_141_), .C(_146_), .Y(_2__2_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_2__2_), .Y(_151_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_152_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_153_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_153_), .C(_152_), .Y(_154_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_148_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_149_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_149_), .C(_2__2_), .Y(_150_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_154_), .Y(_0__2_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_148_), .C(_153_), .Y(_2__3_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_2__3_), .Y(_158_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_159_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_160_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_160_), .C(_159_), .Y(_161_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_155_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_156_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_156_), .C(_2__3_), .Y(_157_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_161_), .Y(_0__3_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_155_), .C(_160_), .Y(_1_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .Y(_165_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_166_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_167_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_167_), .C(_166_), .Y(_168_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_162_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_163_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_163_), .C(w_cout_1_), .Y(_164_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_168_), .Y(_0__4_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_162_), .C(_167_), .Y(_5__1_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_5__1_), .Y(_172_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_173_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_174_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_174_), .C(_173_), .Y(_175_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_169_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_170_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_170_), .C(_5__1_), .Y(_171_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_175_), .Y(_0__5_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_169_), .C(_174_), .Y(_5__2_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_5__2_), .Y(_179_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_180_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_181_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_181_), .C(_180_), .Y(_182_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_176_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_177_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_177_), .C(_5__2_), .Y(_178_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_182_), .Y(_0__6_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_176_), .C(_181_), .Y(_5__3_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_5__3_), .Y(_186_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_187_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_188_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_188_), .C(_187_), .Y(_189_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_183_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_184_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_184_), .C(_5__3_), .Y(_185_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_189_), .Y(_0__7_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_183_), .C(_188_), .Y(_4_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .Y(_193_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_194_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_195_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_195_), .C(_194_), .Y(_196_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_190_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_191_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_191_), .C(w_cout_2_), .Y(_192_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(_196_), .Y(_0__8_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_190_), .C(_195_), .Y(_8__1_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_8__1_), .Y(_200_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_201_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_202_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_202_), .C(_201_), .Y(_203_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_197_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_198_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_198_), .C(_8__1_), .Y(_199_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_203_), .Y(_0__9_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_197_), .C(_202_), .Y(_8__2_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_8__2_), .Y(_207_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_208_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_209_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_209_), .C(_208_), .Y(_210_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_204_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_205_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_205_), .C(_8__2_), .Y(_206_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_210_), .Y(_0__10_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_204_), .C(_209_), .Y(_8__3_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_8__3_), .Y(_214_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_215_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_216_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_216_), .C(_215_), .Y(_217_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_211_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_212_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_212_), .C(_8__3_), .Y(_213_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_217_), .Y(_0__11_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_211_), .C(_216_), .Y(_7_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .Y(_221_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_222_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_223_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_223_), .C(_222_), .Y(_224_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_218_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_219_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(_219_), .C(w_cout_3_), .Y(_220_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_224_), .Y(_0__12_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_218_), .C(_223_), .Y(_11__1_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_11__1_), .Y(_228_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_229_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_230_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_230_), .C(_229_), .Y(_231_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_225_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_226_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_226_), .C(_11__1_), .Y(_227_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_231_), .Y(_0__13_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_225_), .C(_230_), .Y(_11__2_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_11__2_), .Y(_235_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_236_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_237_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_237_), .C(_236_), .Y(_238_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_232_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_233_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_233_), .C(_11__2_), .Y(_234_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_238_), .Y(_0__14_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_232_), .C(_237_), .Y(_11__3_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_11__3_), .Y(_242_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_243_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_244_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_244_), .C(_243_), .Y(_245_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_239_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_240_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_240_), .C(_11__3_), .Y(_241_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_245_), .Y(_0__15_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_239_), .C(_244_), .Y(_10_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .Y(_249_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_250_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_251_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_251_), .C(_250_), .Y(_252_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_246_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_247_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_247_), .C(w_cout_4_), .Y(_248_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_252_), .Y(_0__16_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_246_), .C(_251_), .Y(_14__1_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_14__1_), .Y(_256_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_257_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_258_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_258_), .C(_257_), .Y(_259_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_253_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_254_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_253_), .B(_254_), .C(_14__1_), .Y(_255_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_259_), .Y(_0__17_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_253_), .C(_258_), .Y(_14__2_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_14__2_), .Y(_263_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_264_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_265_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_265_), .C(_264_), .Y(_266_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_260_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_261_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_261_), .C(_14__2_), .Y(_262_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_266_), .Y(_0__18_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_260_), .C(_265_), .Y(_14__3_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_14__3_), .Y(_270_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_271_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_272_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_272_), .C(_271_), .Y(_273_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_267_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_268_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_268_), .C(_14__3_), .Y(_269_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_273_), .Y(_0__19_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_267_), .C(_272_), .Y(_13_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .Y(_277_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_278_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_279_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_279_), .C(_278_), .Y(_280_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_274_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_275_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_275_), .C(w_cout_5_), .Y(_276_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_280_), .Y(_0__20_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_274_), .C(_279_), .Y(_17__1_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_17__1_), .Y(_284_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_285_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_286_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_286_), .C(_285_), .Y(_287_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_281_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_282_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_282_), .C(_17__1_), .Y(_283_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_283_), .B(_287_), .Y(_0__21_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_281_), .C(_286_), .Y(_17__2_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_17__2_), .Y(_291_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_292_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_293_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_293_), .C(_292_), .Y(_294_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_288_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_289_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_289_), .C(_17__2_), .Y(_290_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_294_), .Y(_0__22_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_288_), .C(_293_), .Y(_17__3_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_17__3_), .Y(_298_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_299_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_300_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_300_), .C(_299_), .Y(_301_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_295_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_296_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_296_), .C(_17__3_), .Y(_297_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_301_), .Y(_0__23_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_295_), .C(_300_), .Y(_16_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .Y(_305_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_306_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_307_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_307_), .C(_306_), .Y(_308_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_302_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_303_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_303_), .C(w_cout_6_), .Y(_304_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_308_), .Y(_0__24_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_302_), .C(_307_), .Y(_20__1_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_20__1_), .Y(_312_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_313_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_314_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_314_), .C(_313_), .Y(_315_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_309_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_310_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_310_), .C(_20__1_), .Y(_311_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_315_), .Y(_0__25_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_309_), .C(_314_), .Y(_20__2_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_20__2_), .Y(_319_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_320_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_321_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_321_), .C(_320_), .Y(_322_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_316_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_317_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_316_), .B(_317_), .C(_20__2_), .Y(_318_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_322_), .Y(_0__26_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_316_), .C(_321_), .Y(_20__3_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_20__3_), .Y(_326_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_327_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_328_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_328_), .C(_327_), .Y(_329_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_323_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_324_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_324_), .C(_20__3_), .Y(_325_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_329_), .Y(_0__27_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_323_), .C(_328_), .Y(_19_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_cin), .Y(_333_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_334_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_335_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_335_), .C(_334_), .Y(_336_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_330_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_331_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_331_), .C(cskip1_inst_cin), .Y(_332_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_336_), .Y(cskip1_inst_sum) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_330_), .C(_335_), .Y(cskip1_inst_rca0_w_CARRY_1_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_rca0_w_CARRY_1_), .Y(_338_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_339_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_337_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_337_), .C(_339_), .Y(cskip1_inst_rca0_w_CARRY_2_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_rca0_w_CARRY_2_), .Y(_341_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_342_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_340_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_340_), .C(_342_), .Y(cskip1_inst_rca0_w_CARRY_3_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_rca0_w_CARRY_3_), .Y(_344_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_345_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_343_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_343_), .C(_345_), .Y(cskip1_inst_cout0) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_346_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_347_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_347_), .Y(cskip1_inst_skip0_P) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_cout0), .Y(_348_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(cskip1_inst_skip0_P), .Y(_349_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_skip0_P), .B(_348_), .C(_349_), .Y(w_cout_8_) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_sum), .Y(_0__28_) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_2__0_) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .Y(_5__0_) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(_5__4_) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .Y(_8__0_) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .Y(_11__0_) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(_11__4_) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .Y(_14__0_) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .Y(_17__0_) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_17__4_) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .Y(_20__0_) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_20__4_) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_cin), .Y(cskip1_inst_rca0_w_CARRY_0_) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_cout0), .Y(cskip1_inst_rca0_w_CARRY_4_) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_cin), .Y(w_cout_7_) );
endmodule
