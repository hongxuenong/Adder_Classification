module cla_55bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add1[19], i_add1[20], i_add1[21], i_add1[22], i_add1[23], i_add1[24], i_add1[25], i_add1[26], i_add1[27], i_add1[28], i_add1[29], i_add1[30], i_add1[31], i_add1[32], i_add1[33], i_add1[34], i_add1[35], i_add1[36], i_add1[37], i_add1[38], i_add1[39], i_add1[40], i_add1[41], i_add1[42], i_add1[43], i_add1[44], i_add1[45], i_add1[46], i_add1[47], i_add1[48], i_add1[49], i_add1[50], i_add1[51], i_add1[52], i_add1[53], i_add1[54], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], i_add2[19], i_add2[20], i_add2[21], i_add2[22], i_add2[23], i_add2[24], i_add2[25], i_add2[26], i_add2[27], i_add2[28], i_add2[29], i_add2[30], i_add2[31], i_add2[32], i_add2[33], i_add2[34], i_add2[35], i_add2[36], i_add2[37], i_add2[38], i_add2[39], i_add2[40], i_add2[41], i_add2[42], i_add2[43], i_add2[44], i_add2[45], i_add2[46], i_add2[47], i_add2[48], i_add2[49], i_add2[50], i_add2[51], i_add2[52], i_add2[53], i_add2[54], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21], o_result[22], o_result[23], o_result[24], o_result[25], o_result[26], o_result[27], o_result[28], o_result[29], o_result[30], o_result[31], o_result[32], o_result[33], o_result[34], o_result[35], o_result[36], o_result[37], o_result[38], o_result[39], o_result[40], o_result[41], o_result[42], o_result[43], o_result[44], o_result[45], o_result[46], o_result[47], o_result[48], o_result[49], o_result[50], o_result[51], o_result[52], o_result[53], o_result[54], o_result[55]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add1[19];
input i_add1[20];
input i_add1[21];
input i_add1[22];
input i_add1[23];
input i_add1[24];
input i_add1[25];
input i_add1[26];
input i_add1[27];
input i_add1[28];
input i_add1[29];
input i_add1[30];
input i_add1[31];
input i_add1[32];
input i_add1[33];
input i_add1[34];
input i_add1[35];
input i_add1[36];
input i_add1[37];
input i_add1[38];
input i_add1[39];
input i_add1[40];
input i_add1[41];
input i_add1[42];
input i_add1[43];
input i_add1[44];
input i_add1[45];
input i_add1[46];
input i_add1[47];
input i_add1[48];
input i_add1[49];
input i_add1[50];
input i_add1[51];
input i_add1[52];
input i_add1[53];
input i_add1[54];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
input i_add2[19];
input i_add2[20];
input i_add2[21];
input i_add2[22];
input i_add2[23];
input i_add2[24];
input i_add2[25];
input i_add2[26];
input i_add2[27];
input i_add2[28];
input i_add2[29];
input i_add2[30];
input i_add2[31];
input i_add2[32];
input i_add2[33];
input i_add2[34];
input i_add2[35];
input i_add2[36];
input i_add2[37];
input i_add2[38];
input i_add2[39];
input i_add2[40];
input i_add2[41];
input i_add2[42];
input i_add2[43];
input i_add2[44];
input i_add2[45];
input i_add2[46];
input i_add2[47];
input i_add2[48];
input i_add2[49];
input i_add2[50];
input i_add2[51];
input i_add2[52];
input i_add2[53];
input i_add2[54];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];
output o_result[22];
output o_result[23];
output o_result[24];
output o_result[25];
output o_result[26];
output o_result[27];
output o_result[28];
output o_result[29];
output o_result[30];
output o_result[31];
output o_result[32];
output o_result[33];
output o_result[34];
output o_result[35];
output o_result[36];
output o_result[37];
output o_result[38];
output o_result[39];
output o_result[40];
output o_result[41];
output o_result[42];
output o_result[43];
output o_result[44];
output o_result[45];
output o_result[46];
output o_result[47];
output o_result[48];
output o_result[49];
output o_result[50];
output o_result[51];
output o_result[52];
output o_result[53];
output o_result[54];
output o_result[55];

NOR2X1 NOR2X1_1 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_36_) );
INVX1 INVX1_1 ( .A(_36_), .Y(_37_) );
NAND3X1 NAND3X1_1 ( .A(_35_), .B(_37_), .C(_30_), .Y(_38_) );
OAI21X1 OAI21X1_1 ( .A(_32_), .B(_33_), .C(_38_), .Y(w_C_9_) );
NOR2X1 NOR2X1_2 ( .A(_32_), .B(_33_), .Y(_39_) );
INVX1 INVX1_2 ( .A(_39_), .Y(_40_) );
AND2X2 AND2X2_1 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_41_) );
INVX1 INVX1_3 ( .A(_41_), .Y(_42_) );
NAND3X1 NAND3X1_2 ( .A(_40_), .B(_42_), .C(_38_), .Y(_43_) );
OAI21X1 OAI21X1_2 ( .A(i_add2[9]), .B(i_add1[9]), .C(_43_), .Y(_44_) );
INVX1 INVX1_4 ( .A(_44_), .Y(w_C_10_) );
INVX1 INVX1_5 ( .A(i_add2[10]), .Y(_45_) );
INVX1 INVX1_6 ( .A(i_add1[10]), .Y(_46_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_47_) );
INVX1 INVX1_7 ( .A(_47_), .Y(_48_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_49_) );
INVX1 INVX1_8 ( .A(_49_), .Y(_50_) );
NAND3X1 NAND3X1_3 ( .A(_48_), .B(_50_), .C(_43_), .Y(_51_) );
OAI21X1 OAI21X1_3 ( .A(_45_), .B(_46_), .C(_51_), .Y(w_C_11_) );
NOR2X1 NOR2X1_5 ( .A(_45_), .B(_46_), .Y(_52_) );
INVX1 INVX1_9 ( .A(_52_), .Y(_53_) );
AND2X2 AND2X2_2 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_54_) );
INVX1 INVX1_10 ( .A(_54_), .Y(_55_) );
NAND3X1 NAND3X1_4 ( .A(_53_), .B(_55_), .C(_51_), .Y(_56_) );
OAI21X1 OAI21X1_4 ( .A(i_add2[11]), .B(i_add1[11]), .C(_56_), .Y(_57_) );
INVX1 INVX1_11 ( .A(_57_), .Y(w_C_12_) );
INVX1 INVX1_12 ( .A(i_add2[12]), .Y(_58_) );
INVX1 INVX1_13 ( .A(i_add1[12]), .Y(_59_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_60_) );
INVX1 INVX1_14 ( .A(_60_), .Y(_61_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_62_) );
INVX1 INVX1_15 ( .A(_62_), .Y(_63_) );
NAND3X1 NAND3X1_5 ( .A(_61_), .B(_63_), .C(_56_), .Y(_64_) );
OAI21X1 OAI21X1_5 ( .A(_58_), .B(_59_), .C(_64_), .Y(w_C_13_) );
NOR2X1 NOR2X1_8 ( .A(_58_), .B(_59_), .Y(_65_) );
INVX1 INVX1_16 ( .A(_65_), .Y(_66_) );
AND2X2 AND2X2_3 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_67_) );
INVX1 INVX1_17 ( .A(_67_), .Y(_68_) );
NAND3X1 NAND3X1_6 ( .A(_66_), .B(_68_), .C(_64_), .Y(_69_) );
OAI21X1 OAI21X1_6 ( .A(i_add2[13]), .B(i_add1[13]), .C(_69_), .Y(_70_) );
INVX1 INVX1_18 ( .A(_70_), .Y(w_C_14_) );
INVX1 INVX1_19 ( .A(i_add2[14]), .Y(_71_) );
INVX1 INVX1_20 ( .A(i_add1[14]), .Y(_72_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_73_) );
INVX1 INVX1_21 ( .A(_73_), .Y(_74_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_75_) );
INVX1 INVX1_22 ( .A(_75_), .Y(_76_) );
NAND3X1 NAND3X1_7 ( .A(_74_), .B(_76_), .C(_69_), .Y(_77_) );
OAI21X1 OAI21X1_7 ( .A(_71_), .B(_72_), .C(_77_), .Y(w_C_15_) );
NOR2X1 NOR2X1_11 ( .A(_71_), .B(_72_), .Y(_78_) );
INVX1 INVX1_23 ( .A(_78_), .Y(_79_) );
AND2X2 AND2X2_4 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_80_) );
INVX1 INVX1_24 ( .A(_80_), .Y(_81_) );
NAND3X1 NAND3X1_8 ( .A(_79_), .B(_81_), .C(_77_), .Y(_82_) );
OAI21X1 OAI21X1_8 ( .A(i_add2[15]), .B(i_add1[15]), .C(_82_), .Y(_83_) );
INVX1 INVX1_25 ( .A(_83_), .Y(w_C_16_) );
INVX1 INVX1_26 ( .A(i_add2[16]), .Y(_84_) );
INVX1 INVX1_27 ( .A(i_add1[16]), .Y(_85_) );
NOR2X1 NOR2X1_12 ( .A(_84_), .B(_85_), .Y(_86_) );
INVX1 INVX1_28 ( .A(_86_), .Y(_87_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_88_) );
INVX1 INVX1_29 ( .A(_88_), .Y(_89_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_90_) );
INVX1 INVX1_30 ( .A(_90_), .Y(_91_) );
NAND3X1 NAND3X1_9 ( .A(_89_), .B(_91_), .C(_82_), .Y(_92_) );
AND2X2 AND2X2_5 ( .A(_92_), .B(_87_), .Y(_93_) );
INVX1 INVX1_31 ( .A(_93_), .Y(w_C_17_) );
AND2X2 AND2X2_6 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_94_) );
INVX1 INVX1_32 ( .A(_94_), .Y(_95_) );
NAND3X1 NAND3X1_10 ( .A(_87_), .B(_95_), .C(_92_), .Y(_96_) );
OAI21X1 OAI21X1_9 ( .A(i_add2[17]), .B(i_add1[17]), .C(_96_), .Y(_97_) );
INVX1 INVX1_33 ( .A(_97_), .Y(w_C_18_) );
INVX1 INVX1_34 ( .A(i_add2[18]), .Y(_98_) );
INVX1 INVX1_35 ( .A(i_add1[18]), .Y(_99_) );
NOR2X1 NOR2X1_15 ( .A(_98_), .B(_99_), .Y(_100_) );
INVX1 INVX1_36 ( .A(_100_), .Y(_101_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_102_) );
INVX1 INVX1_37 ( .A(_102_), .Y(_103_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_104_) );
INVX1 INVX1_38 ( .A(_104_), .Y(_105_) );
NAND3X1 NAND3X1_11 ( .A(_103_), .B(_105_), .C(_96_), .Y(_106_) );
AND2X2 AND2X2_7 ( .A(_106_), .B(_101_), .Y(_107_) );
INVX1 INVX1_39 ( .A(_107_), .Y(w_C_19_) );
AND2X2 AND2X2_8 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_108_) );
INVX1 INVX1_40 ( .A(_108_), .Y(_109_) );
NAND3X1 NAND3X1_12 ( .A(_101_), .B(_109_), .C(_106_), .Y(_110_) );
OAI21X1 OAI21X1_10 ( .A(i_add2[19]), .B(i_add1[19]), .C(_110_), .Y(_111_) );
INVX1 INVX1_41 ( .A(_111_), .Y(w_C_20_) );
INVX1 INVX1_42 ( .A(i_add2[20]), .Y(_112_) );
INVX1 INVX1_43 ( .A(i_add1[20]), .Y(_113_) );
NOR2X1 NOR2X1_18 ( .A(_112_), .B(_113_), .Y(_114_) );
INVX1 INVX1_44 ( .A(_114_), .Y(_115_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_116_) );
INVX1 INVX1_45 ( .A(_116_), .Y(_117_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_118_) );
INVX1 INVX1_46 ( .A(_118_), .Y(_119_) );
NAND3X1 NAND3X1_13 ( .A(_117_), .B(_119_), .C(_110_), .Y(_120_) );
AND2X2 AND2X2_9 ( .A(_120_), .B(_115_), .Y(_121_) );
INVX1 INVX1_47 ( .A(_121_), .Y(w_C_21_) );
AND2X2 AND2X2_10 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_122_) );
INVX1 INVX1_48 ( .A(_122_), .Y(_123_) );
NAND3X1 NAND3X1_14 ( .A(_115_), .B(_123_), .C(_120_), .Y(_124_) );
OAI21X1 OAI21X1_11 ( .A(i_add2[21]), .B(i_add1[21]), .C(_124_), .Y(_125_) );
INVX1 INVX1_49 ( .A(_125_), .Y(w_C_22_) );
INVX1 INVX1_50 ( .A(i_add2[22]), .Y(_126_) );
INVX1 INVX1_51 ( .A(i_add1[22]), .Y(_127_) );
NOR2X1 NOR2X1_21 ( .A(_126_), .B(_127_), .Y(_128_) );
BUFX2 BUFX2_1 ( .A(_333__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_333__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_333__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_333__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_333__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_333__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_333__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_333__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_333__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_333__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_333__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_333__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_333__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_333__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_333__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_333__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_333__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_333__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_333__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_333__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_333__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_333__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_333__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_333__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_333__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_333__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_333__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_333__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_333__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_333__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_333__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_333__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_333__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_333__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_333__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_333__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_333__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(_333__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .A(_333__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .A(_333__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .A(_333__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .A(_333__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .A(_333__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .A(_333__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .A(_333__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .A(_333__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .A(_333__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .A(_333__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .A(_333__48_), .Y(o_result[48]) );
BUFX2 BUFX2_50 ( .A(_333__49_), .Y(o_result[49]) );
BUFX2 BUFX2_51 ( .A(_333__50_), .Y(o_result[50]) );
BUFX2 BUFX2_52 ( .A(_333__51_), .Y(o_result[51]) );
BUFX2 BUFX2_53 ( .A(_333__52_), .Y(o_result[52]) );
BUFX2 BUFX2_54 ( .A(_333__53_), .Y(o_result[53]) );
BUFX2 BUFX2_55 ( .A(_333__54_), .Y(o_result[54]) );
BUFX2 BUFX2_56 ( .A(w_C_55_), .Y(o_result[55]) );
INVX1 INVX1_52 ( .A(w_C_4_), .Y(_337_) );
OR2X2 OR2X2_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_338_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_339_) );
NAND3X1 NAND3X1_15 ( .A(_337_), .B(_339_), .C(_338_), .Y(_340_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_334_) );
AND2X2 AND2X2_11 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_335_) );
OAI21X1 OAI21X1_12 ( .A(_334_), .B(_335_), .C(w_C_4_), .Y(_336_) );
NAND2X1 NAND2X1_2 ( .A(_336_), .B(_340_), .Y(_333__4_) );
INVX1 INVX1_53 ( .A(w_C_5_), .Y(_344_) );
OR2X2 OR2X2_2 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_345_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_346_) );
NAND3X1 NAND3X1_16 ( .A(_344_), .B(_346_), .C(_345_), .Y(_347_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_341_) );
AND2X2 AND2X2_12 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_342_) );
OAI21X1 OAI21X1_13 ( .A(_341_), .B(_342_), .C(w_C_5_), .Y(_343_) );
NAND2X1 NAND2X1_4 ( .A(_343_), .B(_347_), .Y(_333__5_) );
INVX1 INVX1_54 ( .A(w_C_6_), .Y(_351_) );
OR2X2 OR2X2_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_352_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_353_) );
NAND3X1 NAND3X1_17 ( .A(_351_), .B(_353_), .C(_352_), .Y(_354_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_348_) );
AND2X2 AND2X2_13 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_349_) );
OAI21X1 OAI21X1_14 ( .A(_348_), .B(_349_), .C(w_C_6_), .Y(_350_) );
NAND2X1 NAND2X1_6 ( .A(_350_), .B(_354_), .Y(_333__6_) );
INVX1 INVX1_55 ( .A(w_C_7_), .Y(_358_) );
OR2X2 OR2X2_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_359_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_360_) );
NAND3X1 NAND3X1_18 ( .A(_358_), .B(_360_), .C(_359_), .Y(_361_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_355_) );
AND2X2 AND2X2_14 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_356_) );
OAI21X1 OAI21X1_15 ( .A(_355_), .B(_356_), .C(w_C_7_), .Y(_357_) );
NAND2X1 NAND2X1_8 ( .A(_357_), .B(_361_), .Y(_333__7_) );
INVX1 INVX1_56 ( .A(w_C_8_), .Y(_365_) );
OR2X2 OR2X2_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_366_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_367_) );
NAND3X1 NAND3X1_19 ( .A(_365_), .B(_367_), .C(_366_), .Y(_368_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_362_) );
AND2X2 AND2X2_15 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_363_) );
OAI21X1 OAI21X1_16 ( .A(_362_), .B(_363_), .C(w_C_8_), .Y(_364_) );
NAND2X1 NAND2X1_10 ( .A(_364_), .B(_368_), .Y(_333__8_) );
INVX1 INVX1_57 ( .A(w_C_9_), .Y(_372_) );
OR2X2 OR2X2_6 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_373_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_374_) );
NAND3X1 NAND3X1_20 ( .A(_372_), .B(_374_), .C(_373_), .Y(_375_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_369_) );
AND2X2 AND2X2_16 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_370_) );
OAI21X1 OAI21X1_17 ( .A(_369_), .B(_370_), .C(w_C_9_), .Y(_371_) );
NAND2X1 NAND2X1_12 ( .A(_371_), .B(_375_), .Y(_333__9_) );
INVX1 INVX1_58 ( .A(w_C_10_), .Y(_379_) );
OR2X2 OR2X2_7 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_380_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_381_) );
NAND3X1 NAND3X1_21 ( .A(_379_), .B(_381_), .C(_380_), .Y(_382_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_376_) );
AND2X2 AND2X2_17 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_377_) );
OAI21X1 OAI21X1_18 ( .A(_376_), .B(_377_), .C(w_C_10_), .Y(_378_) );
NAND2X1 NAND2X1_14 ( .A(_378_), .B(_382_), .Y(_333__10_) );
INVX1 INVX1_59 ( .A(w_C_11_), .Y(_386_) );
OR2X2 OR2X2_8 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_387_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_388_) );
NAND3X1 NAND3X1_22 ( .A(_386_), .B(_388_), .C(_387_), .Y(_389_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_383_) );
AND2X2 AND2X2_18 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_384_) );
OAI21X1 OAI21X1_19 ( .A(_383_), .B(_384_), .C(w_C_11_), .Y(_385_) );
NAND2X1 NAND2X1_16 ( .A(_385_), .B(_389_), .Y(_333__11_) );
INVX1 INVX1_60 ( .A(w_C_12_), .Y(_393_) );
OR2X2 OR2X2_9 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_394_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_395_) );
NAND3X1 NAND3X1_23 ( .A(_393_), .B(_395_), .C(_394_), .Y(_396_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_390_) );
AND2X2 AND2X2_19 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_391_) );
OAI21X1 OAI21X1_20 ( .A(_390_), .B(_391_), .C(w_C_12_), .Y(_392_) );
NAND2X1 NAND2X1_18 ( .A(_392_), .B(_396_), .Y(_333__12_) );
INVX1 INVX1_61 ( .A(w_C_13_), .Y(_400_) );
OR2X2 OR2X2_10 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_401_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_402_) );
NAND3X1 NAND3X1_24 ( .A(_400_), .B(_402_), .C(_401_), .Y(_403_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_397_) );
AND2X2 AND2X2_20 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_398_) );
OAI21X1 OAI21X1_21 ( .A(_397_), .B(_398_), .C(w_C_13_), .Y(_399_) );
NAND2X1 NAND2X1_20 ( .A(_399_), .B(_403_), .Y(_333__13_) );
INVX1 INVX1_62 ( .A(w_C_14_), .Y(_407_) );
OR2X2 OR2X2_11 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_408_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_409_) );
NAND3X1 NAND3X1_25 ( .A(_407_), .B(_409_), .C(_408_), .Y(_410_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_404_) );
AND2X2 AND2X2_21 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_405_) );
OAI21X1 OAI21X1_22 ( .A(_404_), .B(_405_), .C(w_C_14_), .Y(_406_) );
NAND2X1 NAND2X1_22 ( .A(_406_), .B(_410_), .Y(_333__14_) );
INVX1 INVX1_63 ( .A(w_C_15_), .Y(_414_) );
OR2X2 OR2X2_12 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_415_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_416_) );
NAND3X1 NAND3X1_26 ( .A(_414_), .B(_416_), .C(_415_), .Y(_417_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_411_) );
AND2X2 AND2X2_22 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_412_) );
OAI21X1 OAI21X1_23 ( .A(_411_), .B(_412_), .C(w_C_15_), .Y(_413_) );
NAND2X1 NAND2X1_24 ( .A(_413_), .B(_417_), .Y(_333__15_) );
INVX1 INVX1_64 ( .A(w_C_16_), .Y(_421_) );
OR2X2 OR2X2_13 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_422_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_423_) );
NAND3X1 NAND3X1_27 ( .A(_421_), .B(_423_), .C(_422_), .Y(_424_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_418_) );
AND2X2 AND2X2_23 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_419_) );
OAI21X1 OAI21X1_24 ( .A(_418_), .B(_419_), .C(w_C_16_), .Y(_420_) );
NAND2X1 NAND2X1_26 ( .A(_420_), .B(_424_), .Y(_333__16_) );
INVX1 INVX1_65 ( .A(w_C_17_), .Y(_428_) );
OR2X2 OR2X2_14 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_429_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_430_) );
NAND3X1 NAND3X1_28 ( .A(_428_), .B(_430_), .C(_429_), .Y(_431_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_425_) );
AND2X2 AND2X2_24 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_426_) );
OAI21X1 OAI21X1_25 ( .A(_425_), .B(_426_), .C(w_C_17_), .Y(_427_) );
NAND2X1 NAND2X1_28 ( .A(_427_), .B(_431_), .Y(_333__17_) );
INVX1 INVX1_66 ( .A(w_C_18_), .Y(_435_) );
OR2X2 OR2X2_15 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_436_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_437_) );
NAND3X1 NAND3X1_29 ( .A(_435_), .B(_437_), .C(_436_), .Y(_438_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_432_) );
AND2X2 AND2X2_25 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_433_) );
OAI21X1 OAI21X1_26 ( .A(_432_), .B(_433_), .C(w_C_18_), .Y(_434_) );
NAND2X1 NAND2X1_30 ( .A(_434_), .B(_438_), .Y(_333__18_) );
INVX1 INVX1_67 ( .A(w_C_19_), .Y(_442_) );
OR2X2 OR2X2_16 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_443_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_444_) );
NAND3X1 NAND3X1_30 ( .A(_442_), .B(_444_), .C(_443_), .Y(_445_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_439_) );
AND2X2 AND2X2_26 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_440_) );
OAI21X1 OAI21X1_27 ( .A(_439_), .B(_440_), .C(w_C_19_), .Y(_441_) );
NAND2X1 NAND2X1_32 ( .A(_441_), .B(_445_), .Y(_333__19_) );
INVX1 INVX1_68 ( .A(w_C_20_), .Y(_449_) );
OR2X2 OR2X2_17 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_450_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_451_) );
NAND3X1 NAND3X1_31 ( .A(_449_), .B(_451_), .C(_450_), .Y(_452_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_446_) );
AND2X2 AND2X2_27 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_447_) );
OAI21X1 OAI21X1_28 ( .A(_446_), .B(_447_), .C(w_C_20_), .Y(_448_) );
NAND2X1 NAND2X1_34 ( .A(_448_), .B(_452_), .Y(_333__20_) );
INVX1 INVX1_69 ( .A(w_C_21_), .Y(_456_) );
OR2X2 OR2X2_18 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_457_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_458_) );
NAND3X1 NAND3X1_32 ( .A(_456_), .B(_458_), .C(_457_), .Y(_459_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_453_) );
AND2X2 AND2X2_28 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_454_) );
OAI21X1 OAI21X1_29 ( .A(_453_), .B(_454_), .C(w_C_21_), .Y(_455_) );
NAND2X1 NAND2X1_36 ( .A(_455_), .B(_459_), .Y(_333__21_) );
INVX1 INVX1_70 ( .A(w_C_22_), .Y(_463_) );
OR2X2 OR2X2_19 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_464_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_465_) );
NAND3X1 NAND3X1_33 ( .A(_463_), .B(_465_), .C(_464_), .Y(_466_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_460_) );
AND2X2 AND2X2_29 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_461_) );
OAI21X1 OAI21X1_30 ( .A(_460_), .B(_461_), .C(w_C_22_), .Y(_462_) );
NAND2X1 NAND2X1_38 ( .A(_462_), .B(_466_), .Y(_333__22_) );
INVX1 INVX1_71 ( .A(w_C_23_), .Y(_470_) );
OR2X2 OR2X2_20 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_471_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_472_) );
NAND3X1 NAND3X1_34 ( .A(_470_), .B(_472_), .C(_471_), .Y(_473_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_467_) );
AND2X2 AND2X2_30 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_468_) );
OAI21X1 OAI21X1_31 ( .A(_467_), .B(_468_), .C(w_C_23_), .Y(_469_) );
NAND2X1 NAND2X1_40 ( .A(_469_), .B(_473_), .Y(_333__23_) );
INVX1 INVX1_72 ( .A(w_C_24_), .Y(_477_) );
OR2X2 OR2X2_21 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_478_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_479_) );
NAND3X1 NAND3X1_35 ( .A(_477_), .B(_479_), .C(_478_), .Y(_480_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_474_) );
AND2X2 AND2X2_31 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_475_) );
OAI21X1 OAI21X1_32 ( .A(_474_), .B(_475_), .C(w_C_24_), .Y(_476_) );
NAND2X1 NAND2X1_42 ( .A(_476_), .B(_480_), .Y(_333__24_) );
INVX1 INVX1_73 ( .A(w_C_25_), .Y(_484_) );
OR2X2 OR2X2_22 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_485_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_486_) );
NAND3X1 NAND3X1_36 ( .A(_484_), .B(_486_), .C(_485_), .Y(_487_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_481_) );
AND2X2 AND2X2_32 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_482_) );
OAI21X1 OAI21X1_33 ( .A(_481_), .B(_482_), .C(w_C_25_), .Y(_483_) );
NAND2X1 NAND2X1_44 ( .A(_483_), .B(_487_), .Y(_333__25_) );
INVX1 INVX1_74 ( .A(w_C_26_), .Y(_491_) );
OR2X2 OR2X2_23 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_492_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_493_) );
NAND3X1 NAND3X1_37 ( .A(_491_), .B(_493_), .C(_492_), .Y(_494_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_488_) );
AND2X2 AND2X2_33 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_489_) );
OAI21X1 OAI21X1_34 ( .A(_488_), .B(_489_), .C(w_C_26_), .Y(_490_) );
NAND2X1 NAND2X1_46 ( .A(_490_), .B(_494_), .Y(_333__26_) );
INVX1 INVX1_75 ( .A(w_C_27_), .Y(_498_) );
OR2X2 OR2X2_24 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_499_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_500_) );
NAND3X1 NAND3X1_38 ( .A(_498_), .B(_500_), .C(_499_), .Y(_501_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_495_) );
AND2X2 AND2X2_34 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_496_) );
OAI21X1 OAI21X1_35 ( .A(_495_), .B(_496_), .C(w_C_27_), .Y(_497_) );
NAND2X1 NAND2X1_48 ( .A(_497_), .B(_501_), .Y(_333__27_) );
INVX1 INVX1_76 ( .A(w_C_28_), .Y(_505_) );
OR2X2 OR2X2_25 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_506_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_507_) );
NAND3X1 NAND3X1_39 ( .A(_505_), .B(_507_), .C(_506_), .Y(_508_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_502_) );
AND2X2 AND2X2_35 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_503_) );
OAI21X1 OAI21X1_36 ( .A(_502_), .B(_503_), .C(w_C_28_), .Y(_504_) );
NAND2X1 NAND2X1_50 ( .A(_504_), .B(_508_), .Y(_333__28_) );
INVX1 INVX1_77 ( .A(w_C_29_), .Y(_512_) );
OR2X2 OR2X2_26 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_513_) );
NAND2X1 NAND2X1_51 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_514_) );
NAND3X1 NAND3X1_40 ( .A(_512_), .B(_514_), .C(_513_), .Y(_515_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_509_) );
AND2X2 AND2X2_36 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_510_) );
OAI21X1 OAI21X1_37 ( .A(_509_), .B(_510_), .C(w_C_29_), .Y(_511_) );
NAND2X1 NAND2X1_52 ( .A(_511_), .B(_515_), .Y(_333__29_) );
INVX1 INVX1_78 ( .A(w_C_30_), .Y(_519_) );
OR2X2 OR2X2_27 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_520_) );
NAND2X1 NAND2X1_53 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_521_) );
NAND3X1 NAND3X1_41 ( .A(_519_), .B(_521_), .C(_520_), .Y(_522_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_516_) );
AND2X2 AND2X2_37 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_517_) );
OAI21X1 OAI21X1_38 ( .A(_516_), .B(_517_), .C(w_C_30_), .Y(_518_) );
NAND2X1 NAND2X1_54 ( .A(_518_), .B(_522_), .Y(_333__30_) );
INVX1 INVX1_79 ( .A(w_C_31_), .Y(_526_) );
OR2X2 OR2X2_28 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_527_) );
NAND2X1 NAND2X1_55 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_528_) );
NAND3X1 NAND3X1_42 ( .A(_526_), .B(_528_), .C(_527_), .Y(_529_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_523_) );
AND2X2 AND2X2_38 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_524_) );
OAI21X1 OAI21X1_39 ( .A(_523_), .B(_524_), .C(w_C_31_), .Y(_525_) );
NAND2X1 NAND2X1_56 ( .A(_525_), .B(_529_), .Y(_333__31_) );
INVX1 INVX1_80 ( .A(w_C_32_), .Y(_533_) );
OR2X2 OR2X2_29 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_534_) );
NAND2X1 NAND2X1_57 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_535_) );
NAND3X1 NAND3X1_43 ( .A(_533_), .B(_535_), .C(_534_), .Y(_536_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_530_) );
AND2X2 AND2X2_39 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_531_) );
OAI21X1 OAI21X1_40 ( .A(_530_), .B(_531_), .C(w_C_32_), .Y(_532_) );
NAND2X1 NAND2X1_58 ( .A(_532_), .B(_536_), .Y(_333__32_) );
INVX1 INVX1_81 ( .A(w_C_33_), .Y(_540_) );
OR2X2 OR2X2_30 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_541_) );
NAND2X1 NAND2X1_59 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_542_) );
NAND3X1 NAND3X1_44 ( .A(_540_), .B(_542_), .C(_541_), .Y(_543_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_537_) );
AND2X2 AND2X2_40 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_538_) );
OAI21X1 OAI21X1_41 ( .A(_537_), .B(_538_), .C(w_C_33_), .Y(_539_) );
NAND2X1 NAND2X1_60 ( .A(_539_), .B(_543_), .Y(_333__33_) );
INVX1 INVX1_82 ( .A(w_C_34_), .Y(_547_) );
OR2X2 OR2X2_31 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_548_) );
NAND2X1 NAND2X1_61 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_549_) );
NAND3X1 NAND3X1_45 ( .A(_547_), .B(_549_), .C(_548_), .Y(_550_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_544_) );
AND2X2 AND2X2_41 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_545_) );
OAI21X1 OAI21X1_42 ( .A(_544_), .B(_545_), .C(w_C_34_), .Y(_546_) );
NAND2X1 NAND2X1_62 ( .A(_546_), .B(_550_), .Y(_333__34_) );
INVX1 INVX1_83 ( .A(w_C_35_), .Y(_554_) );
OR2X2 OR2X2_32 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_555_) );
NAND2X1 NAND2X1_63 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_556_) );
NAND3X1 NAND3X1_46 ( .A(_554_), .B(_556_), .C(_555_), .Y(_557_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_551_) );
AND2X2 AND2X2_42 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_552_) );
OAI21X1 OAI21X1_43 ( .A(_551_), .B(_552_), .C(w_C_35_), .Y(_553_) );
NAND2X1 NAND2X1_64 ( .A(_553_), .B(_557_), .Y(_333__35_) );
INVX1 INVX1_84 ( .A(w_C_36_), .Y(_561_) );
OR2X2 OR2X2_33 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_562_) );
NAND2X1 NAND2X1_65 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_563_) );
NAND3X1 NAND3X1_47 ( .A(_561_), .B(_563_), .C(_562_), .Y(_564_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_558_) );
AND2X2 AND2X2_43 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_559_) );
OAI21X1 OAI21X1_44 ( .A(_558_), .B(_559_), .C(w_C_36_), .Y(_560_) );
NAND2X1 NAND2X1_66 ( .A(_560_), .B(_564_), .Y(_333__36_) );
INVX1 INVX1_85 ( .A(w_C_37_), .Y(_568_) );
OR2X2 OR2X2_34 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_569_) );
NAND2X1 NAND2X1_67 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_570_) );
NAND3X1 NAND3X1_48 ( .A(_568_), .B(_570_), .C(_569_), .Y(_571_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_565_) );
AND2X2 AND2X2_44 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_566_) );
OAI21X1 OAI21X1_45 ( .A(_565_), .B(_566_), .C(w_C_37_), .Y(_567_) );
NAND2X1 NAND2X1_68 ( .A(_567_), .B(_571_), .Y(_333__37_) );
INVX1 INVX1_86 ( .A(w_C_38_), .Y(_575_) );
OR2X2 OR2X2_35 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_576_) );
NAND2X1 NAND2X1_69 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_577_) );
NAND3X1 NAND3X1_49 ( .A(_575_), .B(_577_), .C(_576_), .Y(_578_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_572_) );
AND2X2 AND2X2_45 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_573_) );
OAI21X1 OAI21X1_46 ( .A(_572_), .B(_573_), .C(w_C_38_), .Y(_574_) );
NAND2X1 NAND2X1_70 ( .A(_574_), .B(_578_), .Y(_333__38_) );
INVX1 INVX1_87 ( .A(w_C_39_), .Y(_582_) );
OR2X2 OR2X2_36 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_583_) );
NAND2X1 NAND2X1_71 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_584_) );
NAND3X1 NAND3X1_50 ( .A(_582_), .B(_584_), .C(_583_), .Y(_585_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_579_) );
AND2X2 AND2X2_46 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_580_) );
OAI21X1 OAI21X1_47 ( .A(_579_), .B(_580_), .C(w_C_39_), .Y(_581_) );
NAND2X1 NAND2X1_72 ( .A(_581_), .B(_585_), .Y(_333__39_) );
INVX1 INVX1_88 ( .A(w_C_40_), .Y(_589_) );
OR2X2 OR2X2_37 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_590_) );
NAND2X1 NAND2X1_73 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_591_) );
NAND3X1 NAND3X1_51 ( .A(_589_), .B(_591_), .C(_590_), .Y(_592_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_586_) );
AND2X2 AND2X2_47 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_587_) );
OAI21X1 OAI21X1_48 ( .A(_586_), .B(_587_), .C(w_C_40_), .Y(_588_) );
NAND2X1 NAND2X1_74 ( .A(_588_), .B(_592_), .Y(_333__40_) );
INVX1 INVX1_89 ( .A(w_C_41_), .Y(_596_) );
OR2X2 OR2X2_38 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_597_) );
NAND2X1 NAND2X1_75 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_598_) );
NAND3X1 NAND3X1_52 ( .A(_596_), .B(_598_), .C(_597_), .Y(_599_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_593_) );
AND2X2 AND2X2_48 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_594_) );
OAI21X1 OAI21X1_49 ( .A(_593_), .B(_594_), .C(w_C_41_), .Y(_595_) );
NAND2X1 NAND2X1_76 ( .A(_595_), .B(_599_), .Y(_333__41_) );
INVX1 INVX1_90 ( .A(w_C_42_), .Y(_603_) );
OR2X2 OR2X2_39 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_604_) );
NAND2X1 NAND2X1_77 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_605_) );
NAND3X1 NAND3X1_53 ( .A(_603_), .B(_605_), .C(_604_), .Y(_606_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_600_) );
AND2X2 AND2X2_49 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_601_) );
OAI21X1 OAI21X1_50 ( .A(_600_), .B(_601_), .C(w_C_42_), .Y(_602_) );
NAND2X1 NAND2X1_78 ( .A(_602_), .B(_606_), .Y(_333__42_) );
INVX1 INVX1_91 ( .A(w_C_43_), .Y(_610_) );
OR2X2 OR2X2_40 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_611_) );
NAND2X1 NAND2X1_79 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_612_) );
NAND3X1 NAND3X1_54 ( .A(_610_), .B(_612_), .C(_611_), .Y(_613_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_607_) );
AND2X2 AND2X2_50 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_608_) );
OAI21X1 OAI21X1_51 ( .A(_607_), .B(_608_), .C(w_C_43_), .Y(_609_) );
NAND2X1 NAND2X1_80 ( .A(_609_), .B(_613_), .Y(_333__43_) );
INVX1 INVX1_92 ( .A(w_C_44_), .Y(_617_) );
OR2X2 OR2X2_41 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_618_) );
NAND2X1 NAND2X1_81 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_619_) );
NAND3X1 NAND3X1_55 ( .A(_617_), .B(_619_), .C(_618_), .Y(_620_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_614_) );
AND2X2 AND2X2_51 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_615_) );
OAI21X1 OAI21X1_52 ( .A(_614_), .B(_615_), .C(w_C_44_), .Y(_616_) );
NAND2X1 NAND2X1_82 ( .A(_616_), .B(_620_), .Y(_333__44_) );
INVX1 INVX1_93 ( .A(w_C_45_), .Y(_624_) );
OR2X2 OR2X2_42 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_625_) );
NAND2X1 NAND2X1_83 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_626_) );
NAND3X1 NAND3X1_56 ( .A(_624_), .B(_626_), .C(_625_), .Y(_627_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_621_) );
AND2X2 AND2X2_52 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_622_) );
OAI21X1 OAI21X1_53 ( .A(_621_), .B(_622_), .C(w_C_45_), .Y(_623_) );
NAND2X1 NAND2X1_84 ( .A(_623_), .B(_627_), .Y(_333__45_) );
INVX1 INVX1_94 ( .A(w_C_46_), .Y(_631_) );
OR2X2 OR2X2_43 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_632_) );
NAND2X1 NAND2X1_85 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_633_) );
NAND3X1 NAND3X1_57 ( .A(_631_), .B(_633_), .C(_632_), .Y(_634_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_628_) );
AND2X2 AND2X2_53 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_629_) );
OAI21X1 OAI21X1_54 ( .A(_628_), .B(_629_), .C(w_C_46_), .Y(_630_) );
NAND2X1 NAND2X1_86 ( .A(_630_), .B(_634_), .Y(_333__46_) );
INVX1 INVX1_95 ( .A(w_C_47_), .Y(_638_) );
OR2X2 OR2X2_44 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_639_) );
NAND2X1 NAND2X1_87 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_640_) );
NAND3X1 NAND3X1_58 ( .A(_638_), .B(_640_), .C(_639_), .Y(_641_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_635_) );
AND2X2 AND2X2_54 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_636_) );
OAI21X1 OAI21X1_55 ( .A(_635_), .B(_636_), .C(w_C_47_), .Y(_637_) );
NAND2X1 NAND2X1_88 ( .A(_637_), .B(_641_), .Y(_333__47_) );
INVX1 INVX1_96 ( .A(w_C_48_), .Y(_645_) );
OR2X2 OR2X2_45 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_646_) );
NAND2X1 NAND2X1_89 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_647_) );
NAND3X1 NAND3X1_59 ( .A(_645_), .B(_647_), .C(_646_), .Y(_648_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_642_) );
AND2X2 AND2X2_55 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_643_) );
OAI21X1 OAI21X1_56 ( .A(_642_), .B(_643_), .C(w_C_48_), .Y(_644_) );
NAND2X1 NAND2X1_90 ( .A(_644_), .B(_648_), .Y(_333__48_) );
INVX1 INVX1_97 ( .A(w_C_49_), .Y(_652_) );
OR2X2 OR2X2_46 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_653_) );
NAND2X1 NAND2X1_91 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_654_) );
NAND3X1 NAND3X1_60 ( .A(_652_), .B(_654_), .C(_653_), .Y(_655_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_649_) );
AND2X2 AND2X2_56 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_650_) );
OAI21X1 OAI21X1_57 ( .A(_649_), .B(_650_), .C(w_C_49_), .Y(_651_) );
NAND2X1 NAND2X1_92 ( .A(_651_), .B(_655_), .Y(_333__49_) );
INVX1 INVX1_98 ( .A(w_C_50_), .Y(_659_) );
OR2X2 OR2X2_47 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_660_) );
NAND2X1 NAND2X1_93 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_661_) );
NAND3X1 NAND3X1_61 ( .A(_659_), .B(_661_), .C(_660_), .Y(_662_) );
NOR2X1 NOR2X1_68 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_656_) );
AND2X2 AND2X2_57 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_657_) );
OAI21X1 OAI21X1_58 ( .A(_656_), .B(_657_), .C(w_C_50_), .Y(_658_) );
NAND2X1 NAND2X1_94 ( .A(_658_), .B(_662_), .Y(_333__50_) );
INVX1 INVX1_99 ( .A(w_C_51_), .Y(_666_) );
OR2X2 OR2X2_48 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_667_) );
NAND2X1 NAND2X1_95 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_668_) );
NAND3X1 NAND3X1_62 ( .A(_666_), .B(_668_), .C(_667_), .Y(_669_) );
NOR2X1 NOR2X1_69 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_663_) );
AND2X2 AND2X2_58 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_664_) );
OAI21X1 OAI21X1_59 ( .A(_663_), .B(_664_), .C(w_C_51_), .Y(_665_) );
NAND2X1 NAND2X1_96 ( .A(_665_), .B(_669_), .Y(_333__51_) );
INVX1 INVX1_100 ( .A(w_C_52_), .Y(_673_) );
OR2X2 OR2X2_49 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_674_) );
NAND2X1 NAND2X1_97 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_675_) );
NAND3X1 NAND3X1_63 ( .A(_673_), .B(_675_), .C(_674_), .Y(_676_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_670_) );
AND2X2 AND2X2_59 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_671_) );
OAI21X1 OAI21X1_60 ( .A(_670_), .B(_671_), .C(w_C_52_), .Y(_672_) );
NAND2X1 NAND2X1_98 ( .A(_672_), .B(_676_), .Y(_333__52_) );
INVX1 INVX1_101 ( .A(w_C_53_), .Y(_680_) );
OR2X2 OR2X2_50 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_681_) );
NAND2X1 NAND2X1_99 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_682_) );
NAND3X1 NAND3X1_64 ( .A(_680_), .B(_682_), .C(_681_), .Y(_683_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_677_) );
AND2X2 AND2X2_60 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_678_) );
OAI21X1 OAI21X1_61 ( .A(_677_), .B(_678_), .C(w_C_53_), .Y(_679_) );
NAND2X1 NAND2X1_100 ( .A(_679_), .B(_683_), .Y(_333__53_) );
INVX1 INVX1_102 ( .A(w_C_54_), .Y(_687_) );
OR2X2 OR2X2_51 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_688_) );
NAND2X1 NAND2X1_101 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_689_) );
NAND3X1 NAND3X1_65 ( .A(_687_), .B(_689_), .C(_688_), .Y(_690_) );
NOR2X1 NOR2X1_72 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_684_) );
AND2X2 AND2X2_61 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_685_) );
OAI21X1 OAI21X1_62 ( .A(_684_), .B(_685_), .C(w_C_54_), .Y(_686_) );
NAND2X1 NAND2X1_102 ( .A(_686_), .B(_690_), .Y(_333__54_) );
INVX1 INVX1_103 ( .A(1'b0), .Y(_694_) );
OR2X2 OR2X2_52 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_695_) );
NAND2X1 NAND2X1_103 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_696_) );
NAND3X1 NAND3X1_66 ( .A(_694_), .B(_696_), .C(_695_), .Y(_697_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_691_) );
AND2X2 AND2X2_62 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_692_) );
OAI21X1 OAI21X1_63 ( .A(_691_), .B(_692_), .C(1'b0), .Y(_693_) );
NAND2X1 NAND2X1_104 ( .A(_693_), .B(_697_), .Y(_333__0_) );
INVX1 INVX1_104 ( .A(w_C_1_), .Y(_701_) );
OR2X2 OR2X2_53 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_702_) );
NAND2X1 NAND2X1_105 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_703_) );
NAND3X1 NAND3X1_67 ( .A(_701_), .B(_703_), .C(_702_), .Y(_704_) );
NOR2X1 NOR2X1_74 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_698_) );
AND2X2 AND2X2_63 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_699_) );
OAI21X1 OAI21X1_64 ( .A(_698_), .B(_699_), .C(w_C_1_), .Y(_700_) );
NAND2X1 NAND2X1_106 ( .A(_700_), .B(_704_), .Y(_333__1_) );
INVX1 INVX1_105 ( .A(w_C_2_), .Y(_708_) );
OR2X2 OR2X2_54 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_709_) );
NAND2X1 NAND2X1_107 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_710_) );
NAND3X1 NAND3X1_68 ( .A(_708_), .B(_710_), .C(_709_), .Y(_711_) );
NOR2X1 NOR2X1_75 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_705_) );
AND2X2 AND2X2_64 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_706_) );
OAI21X1 OAI21X1_65 ( .A(_705_), .B(_706_), .C(w_C_2_), .Y(_707_) );
NAND2X1 NAND2X1_108 ( .A(_707_), .B(_711_), .Y(_333__2_) );
INVX1 INVX1_106 ( .A(w_C_3_), .Y(_715_) );
OR2X2 OR2X2_55 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_716_) );
NAND2X1 NAND2X1_109 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_717_) );
NAND3X1 NAND3X1_69 ( .A(_715_), .B(_717_), .C(_716_), .Y(_718_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_712_) );
AND2X2 AND2X2_65 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_713_) );
OAI21X1 OAI21X1_66 ( .A(_712_), .B(_713_), .C(w_C_3_), .Y(_714_) );
NAND2X1 NAND2X1_110 ( .A(_714_), .B(_718_), .Y(_333__3_) );
INVX1 INVX1_107 ( .A(_128_), .Y(_129_) );
NOR2X1 NOR2X1_77 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_130_) );
INVX1 INVX1_108 ( .A(_130_), .Y(_131_) );
NOR2X1 NOR2X1_78 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_132_) );
INVX1 INVX1_109 ( .A(_132_), .Y(_133_) );
NAND3X1 NAND3X1_70 ( .A(_131_), .B(_133_), .C(_124_), .Y(_134_) );
AND2X2 AND2X2_66 ( .A(_134_), .B(_129_), .Y(_135_) );
INVX1 INVX1_110 ( .A(_135_), .Y(w_C_23_) );
AND2X2 AND2X2_67 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_136_) );
INVX1 INVX1_111 ( .A(_136_), .Y(_137_) );
NAND3X1 NAND3X1_71 ( .A(_129_), .B(_137_), .C(_134_), .Y(_138_) );
OAI21X1 OAI21X1_67 ( .A(i_add2[23]), .B(i_add1[23]), .C(_138_), .Y(_139_) );
INVX1 INVX1_112 ( .A(_139_), .Y(w_C_24_) );
INVX1 INVX1_113 ( .A(i_add2[24]), .Y(_140_) );
INVX1 INVX1_114 ( .A(i_add1[24]), .Y(_141_) );
NOR2X1 NOR2X1_79 ( .A(_140_), .B(_141_), .Y(_142_) );
INVX1 INVX1_115 ( .A(_142_), .Y(_143_) );
NOR2X1 NOR2X1_80 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_144_) );
INVX1 INVX1_116 ( .A(_144_), .Y(_145_) );
NOR2X1 NOR2X1_81 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_146_) );
INVX1 INVX1_117 ( .A(_146_), .Y(_147_) );
NAND3X1 NAND3X1_72 ( .A(_145_), .B(_147_), .C(_138_), .Y(_148_) );
AND2X2 AND2X2_68 ( .A(_148_), .B(_143_), .Y(_149_) );
INVX1 INVX1_118 ( .A(_149_), .Y(w_C_25_) );
AND2X2 AND2X2_69 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_150_) );
INVX1 INVX1_119 ( .A(_150_), .Y(_151_) );
NAND3X1 NAND3X1_73 ( .A(_143_), .B(_151_), .C(_148_), .Y(_152_) );
OAI21X1 OAI21X1_68 ( .A(i_add2[25]), .B(i_add1[25]), .C(_152_), .Y(_153_) );
INVX1 INVX1_120 ( .A(_153_), .Y(w_C_26_) );
INVX1 INVX1_121 ( .A(i_add2[26]), .Y(_154_) );
INVX1 INVX1_122 ( .A(i_add1[26]), .Y(_155_) );
NOR2X1 NOR2X1_82 ( .A(_154_), .B(_155_), .Y(_156_) );
INVX1 INVX1_123 ( .A(_156_), .Y(_157_) );
NOR2X1 NOR2X1_83 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_158_) );
INVX1 INVX1_124 ( .A(_158_), .Y(_159_) );
NOR2X1 NOR2X1_84 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_160_) );
INVX1 INVX1_125 ( .A(_160_), .Y(_161_) );
NAND3X1 NAND3X1_74 ( .A(_159_), .B(_161_), .C(_152_), .Y(_162_) );
AND2X2 AND2X2_70 ( .A(_162_), .B(_157_), .Y(_163_) );
INVX1 INVX1_126 ( .A(_163_), .Y(w_C_27_) );
AND2X2 AND2X2_71 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_164_) );
INVX1 INVX1_127 ( .A(_164_), .Y(_165_) );
NAND3X1 NAND3X1_75 ( .A(_157_), .B(_165_), .C(_162_), .Y(_166_) );
OAI21X1 OAI21X1_69 ( .A(i_add2[27]), .B(i_add1[27]), .C(_166_), .Y(_167_) );
INVX1 INVX1_128 ( .A(_167_), .Y(w_C_28_) );
INVX1 INVX1_129 ( .A(i_add2[28]), .Y(_168_) );
INVX1 INVX1_130 ( .A(i_add1[28]), .Y(_169_) );
NOR2X1 NOR2X1_85 ( .A(_168_), .B(_169_), .Y(_170_) );
INVX1 INVX1_131 ( .A(_170_), .Y(_171_) );
NOR2X1 NOR2X1_86 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_172_) );
INVX1 INVX1_132 ( .A(_172_), .Y(_173_) );
NOR2X1 NOR2X1_87 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_174_) );
INVX1 INVX1_133 ( .A(_174_), .Y(_175_) );
NAND3X1 NAND3X1_76 ( .A(_173_), .B(_175_), .C(_166_), .Y(_176_) );
AND2X2 AND2X2_72 ( .A(_176_), .B(_171_), .Y(_177_) );
INVX1 INVX1_134 ( .A(_177_), .Y(w_C_29_) );
AND2X2 AND2X2_73 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_178_) );
INVX1 INVX1_135 ( .A(_178_), .Y(_179_) );
NAND3X1 NAND3X1_77 ( .A(_171_), .B(_179_), .C(_176_), .Y(_180_) );
OAI21X1 OAI21X1_70 ( .A(i_add2[29]), .B(i_add1[29]), .C(_180_), .Y(_181_) );
INVX1 INVX1_136 ( .A(_181_), .Y(w_C_30_) );
INVX1 INVX1_137 ( .A(i_add2[30]), .Y(_182_) );
INVX1 INVX1_138 ( .A(i_add1[30]), .Y(_183_) );
NOR2X1 NOR2X1_88 ( .A(_182_), .B(_183_), .Y(_184_) );
INVX1 INVX1_139 ( .A(_184_), .Y(_185_) );
NOR2X1 NOR2X1_89 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_186_) );
INVX1 INVX1_140 ( .A(_186_), .Y(_187_) );
NOR2X1 NOR2X1_90 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_188_) );
INVX1 INVX1_141 ( .A(_188_), .Y(_189_) );
NAND3X1 NAND3X1_78 ( .A(_187_), .B(_189_), .C(_180_), .Y(_190_) );
AND2X2 AND2X2_74 ( .A(_190_), .B(_185_), .Y(_191_) );
INVX1 INVX1_142 ( .A(_191_), .Y(w_C_31_) );
AND2X2 AND2X2_75 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_192_) );
INVX1 INVX1_143 ( .A(_192_), .Y(_193_) );
NAND3X1 NAND3X1_79 ( .A(_185_), .B(_193_), .C(_190_), .Y(_194_) );
OAI21X1 OAI21X1_71 ( .A(i_add2[31]), .B(i_add1[31]), .C(_194_), .Y(_195_) );
INVX1 INVX1_144 ( .A(_195_), .Y(w_C_32_) );
INVX1 INVX1_145 ( .A(i_add2[32]), .Y(_196_) );
INVX1 INVX1_146 ( .A(i_add1[32]), .Y(_197_) );
NOR2X1 NOR2X1_91 ( .A(_196_), .B(_197_), .Y(_198_) );
INVX1 INVX1_147 ( .A(_198_), .Y(_199_) );
NOR2X1 NOR2X1_92 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_200_) );
INVX1 INVX1_148 ( .A(_200_), .Y(_201_) );
NOR2X1 NOR2X1_93 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_202_) );
INVX1 INVX1_149 ( .A(_202_), .Y(_203_) );
NAND3X1 NAND3X1_80 ( .A(_201_), .B(_203_), .C(_194_), .Y(_204_) );
AND2X2 AND2X2_76 ( .A(_204_), .B(_199_), .Y(_205_) );
INVX1 INVX1_150 ( .A(_205_), .Y(w_C_33_) );
AND2X2 AND2X2_77 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_206_) );
INVX1 INVX1_151 ( .A(_206_), .Y(_207_) );
NAND3X1 NAND3X1_81 ( .A(_199_), .B(_207_), .C(_204_), .Y(_208_) );
OAI21X1 OAI21X1_72 ( .A(i_add2[33]), .B(i_add1[33]), .C(_208_), .Y(_209_) );
INVX1 INVX1_152 ( .A(_209_), .Y(w_C_34_) );
INVX1 INVX1_153 ( .A(i_add2[34]), .Y(_210_) );
INVX1 INVX1_154 ( .A(i_add1[34]), .Y(_211_) );
NOR2X1 NOR2X1_94 ( .A(_210_), .B(_211_), .Y(_212_) );
INVX1 INVX1_155 ( .A(_212_), .Y(_213_) );
NOR2X1 NOR2X1_95 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_214_) );
INVX1 INVX1_156 ( .A(_214_), .Y(_215_) );
NOR2X1 NOR2X1_96 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_216_) );
INVX1 INVX1_157 ( .A(_216_), .Y(_217_) );
NAND3X1 NAND3X1_82 ( .A(_215_), .B(_217_), .C(_208_), .Y(_218_) );
AND2X2 AND2X2_78 ( .A(_218_), .B(_213_), .Y(_219_) );
INVX1 INVX1_158 ( .A(_219_), .Y(w_C_35_) );
AND2X2 AND2X2_79 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_220_) );
INVX1 INVX1_159 ( .A(_220_), .Y(_221_) );
NAND3X1 NAND3X1_83 ( .A(_213_), .B(_221_), .C(_218_), .Y(_222_) );
OAI21X1 OAI21X1_73 ( .A(i_add2[35]), .B(i_add1[35]), .C(_222_), .Y(_223_) );
INVX1 INVX1_160 ( .A(_223_), .Y(w_C_36_) );
INVX1 INVX1_161 ( .A(i_add2[36]), .Y(_224_) );
INVX1 INVX1_162 ( .A(i_add1[36]), .Y(_225_) );
NOR2X1 NOR2X1_97 ( .A(_224_), .B(_225_), .Y(_226_) );
INVX1 INVX1_163 ( .A(_226_), .Y(_227_) );
NOR2X1 NOR2X1_98 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_228_) );
INVX1 INVX1_164 ( .A(_228_), .Y(_229_) );
NOR2X1 NOR2X1_99 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_230_) );
INVX1 INVX1_165 ( .A(_230_), .Y(_231_) );
NAND3X1 NAND3X1_84 ( .A(_229_), .B(_231_), .C(_222_), .Y(_232_) );
AND2X2 AND2X2_80 ( .A(_232_), .B(_227_), .Y(_233_) );
INVX1 INVX1_166 ( .A(_233_), .Y(w_C_37_) );
AND2X2 AND2X2_81 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_234_) );
INVX1 INVX1_167 ( .A(_234_), .Y(_235_) );
NAND3X1 NAND3X1_85 ( .A(_227_), .B(_235_), .C(_232_), .Y(_236_) );
OAI21X1 OAI21X1_74 ( .A(i_add2[37]), .B(i_add1[37]), .C(_236_), .Y(_237_) );
INVX1 INVX1_168 ( .A(_237_), .Y(w_C_38_) );
INVX1 INVX1_169 ( .A(i_add2[38]), .Y(_238_) );
INVX1 INVX1_170 ( .A(i_add1[38]), .Y(_239_) );
NOR2X1 NOR2X1_100 ( .A(_238_), .B(_239_), .Y(_240_) );
INVX1 INVX1_171 ( .A(_240_), .Y(_241_) );
NOR2X1 NOR2X1_101 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_242_) );
INVX1 INVX1_172 ( .A(_242_), .Y(_243_) );
NOR2X1 NOR2X1_102 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_244_) );
INVX1 INVX1_173 ( .A(_244_), .Y(_245_) );
NAND3X1 NAND3X1_86 ( .A(_243_), .B(_245_), .C(_236_), .Y(_246_) );
AND2X2 AND2X2_82 ( .A(_246_), .B(_241_), .Y(_247_) );
INVX1 INVX1_174 ( .A(_247_), .Y(w_C_39_) );
AND2X2 AND2X2_83 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_248_) );
INVX1 INVX1_175 ( .A(_248_), .Y(_249_) );
NAND3X1 NAND3X1_87 ( .A(_241_), .B(_249_), .C(_246_), .Y(_250_) );
OAI21X1 OAI21X1_75 ( .A(i_add2[39]), .B(i_add1[39]), .C(_250_), .Y(_251_) );
INVX1 INVX1_176 ( .A(_251_), .Y(w_C_40_) );
INVX1 INVX1_177 ( .A(i_add2[40]), .Y(_252_) );
INVX1 INVX1_178 ( .A(i_add1[40]), .Y(_253_) );
NOR2X1 NOR2X1_103 ( .A(_252_), .B(_253_), .Y(_254_) );
INVX1 INVX1_179 ( .A(_254_), .Y(_255_) );
NOR2X1 NOR2X1_104 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_256_) );
INVX1 INVX1_180 ( .A(_256_), .Y(_257_) );
NOR2X1 NOR2X1_105 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_258_) );
INVX1 INVX1_181 ( .A(_258_), .Y(_259_) );
NAND3X1 NAND3X1_88 ( .A(_257_), .B(_259_), .C(_250_), .Y(_260_) );
AND2X2 AND2X2_84 ( .A(_260_), .B(_255_), .Y(_261_) );
INVX1 INVX1_182 ( .A(_261_), .Y(w_C_41_) );
AND2X2 AND2X2_85 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_262_) );
INVX1 INVX1_183 ( .A(_262_), .Y(_263_) );
NAND3X1 NAND3X1_89 ( .A(_255_), .B(_263_), .C(_260_), .Y(_264_) );
OAI21X1 OAI21X1_76 ( .A(i_add2[41]), .B(i_add1[41]), .C(_264_), .Y(_265_) );
INVX1 INVX1_184 ( .A(_265_), .Y(w_C_42_) );
INVX1 INVX1_185 ( .A(i_add2[42]), .Y(_266_) );
INVX1 INVX1_186 ( .A(i_add1[42]), .Y(_267_) );
NOR2X1 NOR2X1_106 ( .A(_266_), .B(_267_), .Y(_268_) );
INVX1 INVX1_187 ( .A(_268_), .Y(_269_) );
NOR2X1 NOR2X1_107 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_270_) );
INVX1 INVX1_188 ( .A(_270_), .Y(_271_) );
NOR2X1 NOR2X1_108 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_272_) );
INVX1 INVX1_189 ( .A(_272_), .Y(_273_) );
NAND3X1 NAND3X1_90 ( .A(_271_), .B(_273_), .C(_264_), .Y(_274_) );
AND2X2 AND2X2_86 ( .A(_274_), .B(_269_), .Y(_275_) );
INVX1 INVX1_190 ( .A(_275_), .Y(w_C_43_) );
AND2X2 AND2X2_87 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_276_) );
INVX1 INVX1_191 ( .A(_276_), .Y(_277_) );
NAND3X1 NAND3X1_91 ( .A(_269_), .B(_277_), .C(_274_), .Y(_278_) );
OAI21X1 OAI21X1_77 ( .A(i_add2[43]), .B(i_add1[43]), .C(_278_), .Y(_279_) );
INVX1 INVX1_192 ( .A(_279_), .Y(w_C_44_) );
NAND2X1 NAND2X1_111 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_280_) );
NOR2X1 NOR2X1_109 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_281_) );
OAI21X1 OAI21X1_78 ( .A(_281_), .B(_279_), .C(_280_), .Y(w_C_45_) );
OR2X2 OR2X2_56 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_282_) );
NOR2X1 NOR2X1_110 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_283_) );
INVX1 INVX1_193 ( .A(_283_), .Y(_284_) );
INVX1 INVX1_194 ( .A(_281_), .Y(_285_) );
NAND3X1 NAND3X1_92 ( .A(_284_), .B(_285_), .C(_278_), .Y(_286_) );
NAND2X1 NAND2X1_112 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_287_) );
NAND3X1 NAND3X1_93 ( .A(_280_), .B(_287_), .C(_286_), .Y(_288_) );
AND2X2 AND2X2_88 ( .A(_288_), .B(_282_), .Y(w_C_46_) );
INVX1 INVX1_195 ( .A(i_add2[46]), .Y(_289_) );
INVX1 INVX1_196 ( .A(i_add1[46]), .Y(_290_) );
NAND2X1 NAND2X1_113 ( .A(_289_), .B(_290_), .Y(_291_) );
NAND3X1 NAND3X1_94 ( .A(_282_), .B(_291_), .C(_288_), .Y(_292_) );
OAI21X1 OAI21X1_79 ( .A(_289_), .B(_290_), .C(_292_), .Y(w_C_47_) );
INVX1 INVX1_197 ( .A(i_add2[47]), .Y(_293_) );
INVX1 INVX1_198 ( .A(i_add1[47]), .Y(_294_) );
NAND2X1 NAND2X1_114 ( .A(_293_), .B(_294_), .Y(_295_) );
NAND2X1 NAND2X1_115 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_296_) );
NAND2X1 NAND2X1_116 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_297_) );
NAND3X1 NAND3X1_95 ( .A(_296_), .B(_297_), .C(_292_), .Y(_298_) );
AND2X2 AND2X2_89 ( .A(_298_), .B(_295_), .Y(w_C_48_) );
INVX1 INVX1_199 ( .A(i_add2[48]), .Y(_299_) );
INVX1 INVX1_200 ( .A(i_add1[48]), .Y(_300_) );
NAND2X1 NAND2X1_117 ( .A(_299_), .B(_300_), .Y(_301_) );
NAND3X1 NAND3X1_96 ( .A(_295_), .B(_301_), .C(_298_), .Y(_302_) );
OAI21X1 OAI21X1_80 ( .A(_299_), .B(_300_), .C(_302_), .Y(w_C_49_) );
INVX1 INVX1_201 ( .A(i_add2[49]), .Y(_303_) );
INVX1 INVX1_202 ( .A(i_add1[49]), .Y(_304_) );
OAI21X1 OAI21X1_81 ( .A(i_add2[49]), .B(i_add1[49]), .C(w_C_49_), .Y(_305_) );
OAI21X1 OAI21X1_82 ( .A(_303_), .B(_304_), .C(_305_), .Y(w_C_50_) );
NOR2X1 NOR2X1_111 ( .A(_303_), .B(_304_), .Y(_306_) );
INVX1 INVX1_203 ( .A(_306_), .Y(_307_) );
AND2X2 AND2X2_90 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_308_) );
INVX1 INVX1_204 ( .A(_308_), .Y(_309_) );
NAND3X1 NAND3X1_97 ( .A(_307_), .B(_309_), .C(_305_), .Y(_310_) );
OAI21X1 OAI21X1_83 ( .A(i_add2[50]), .B(i_add1[50]), .C(_310_), .Y(_311_) );
INVX1 INVX1_205 ( .A(_311_), .Y(w_C_51_) );
NAND2X1 NAND2X1_118 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_312_) );
NOR2X1 NOR2X1_112 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_313_) );
OAI21X1 OAI21X1_84 ( .A(_313_), .B(_311_), .C(_312_), .Y(w_C_52_) );
NAND2X1 NAND2X1_119 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_314_) );
INVX1 INVX1_206 ( .A(_313_), .Y(_315_) );
NOR2X1 NOR2X1_113 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_316_) );
INVX1 INVX1_207 ( .A(_316_), .Y(_317_) );
NOR2X1 NOR2X1_114 ( .A(_299_), .B(_300_), .Y(_318_) );
INVX1 INVX1_208 ( .A(_318_), .Y(_319_) );
NAND3X1 NAND3X1_98 ( .A(_319_), .B(_307_), .C(_302_), .Y(_320_) );
NOR2X1 NOR2X1_115 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_321_) );
INVX1 INVX1_209 ( .A(_321_), .Y(_322_) );
NAND3X1 NAND3X1_99 ( .A(_317_), .B(_322_), .C(_320_), .Y(_323_) );
NAND3X1 NAND3X1_100 ( .A(_309_), .B(_312_), .C(_323_), .Y(_324_) );
OR2X2 OR2X2_57 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_325_) );
NAND3X1 NAND3X1_101 ( .A(_315_), .B(_325_), .C(_324_), .Y(_326_) );
NAND2X1 NAND2X1_120 ( .A(_314_), .B(_326_), .Y(w_C_53_) );
OR2X2 OR2X2_58 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_327_) );
NAND2X1 NAND2X1_121 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_328_) );
NAND3X1 NAND3X1_102 ( .A(_314_), .B(_328_), .C(_326_), .Y(_329_) );
AND2X2 AND2X2_91 ( .A(_329_), .B(_327_), .Y(w_C_54_) );
NAND2X1 NAND2X1_122 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_330_) );
OR2X2 OR2X2_59 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_331_) );
NAND3X1 NAND3X1_103 ( .A(_327_), .B(_331_), .C(_329_), .Y(_332_) );
NAND2X1 NAND2X1_123 ( .A(_330_), .B(_332_), .Y(w_C_55_) );
NAND2X1 NAND2X1_124 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_210 ( .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_125 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_126 ( .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_85 ( .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_211 ( .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_127 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_60 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_61 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_104 ( .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_128 ( .A(_4_), .B(_7_), .Y(w_C_3_) );
INVX1 INVX1_212 ( .A(i_add2[3]), .Y(_8_) );
INVX1 INVX1_213 ( .A(i_add1[3]), .Y(_9_) );
NAND2X1 NAND2X1_129 ( .A(_8_), .B(_9_), .Y(_10_) );
NAND2X1 NAND2X1_130 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_11_) );
NAND3X1 NAND3X1_105 ( .A(_4_), .B(_11_), .C(_7_), .Y(_12_) );
AND2X2 AND2X2_92 ( .A(_12_), .B(_10_), .Y(w_C_4_) );
NAND2X1 NAND2X1_131 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
OR2X2 OR2X2_62 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_14_) );
NAND3X1 NAND3X1_106 ( .A(_10_), .B(_14_), .C(_12_), .Y(_15_) );
NAND2X1 NAND2X1_132 ( .A(_13_), .B(_15_), .Y(w_C_5_) );
NAND2X1 NAND2X1_133 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_16_) );
NAND3X1 NAND3X1_107 ( .A(_13_), .B(_16_), .C(_15_), .Y(_17_) );
OAI21X1 OAI21X1_86 ( .A(i_add2[5]), .B(i_add1[5]), .C(_17_), .Y(_18_) );
INVX1 INVX1_214 ( .A(_18_), .Y(w_C_6_) );
INVX1 INVX1_215 ( .A(i_add2[6]), .Y(_19_) );
INVX1 INVX1_216 ( .A(i_add1[6]), .Y(_20_) );
NOR2X1 NOR2X1_116 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_21_) );
INVX1 INVX1_217 ( .A(_21_), .Y(_22_) );
NOR2X1 NOR2X1_117 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_23_) );
INVX1 INVX1_218 ( .A(_23_), .Y(_24_) );
NAND3X1 NAND3X1_108 ( .A(_22_), .B(_24_), .C(_17_), .Y(_25_) );
OAI21X1 OAI21X1_87 ( .A(_19_), .B(_20_), .C(_25_), .Y(w_C_7_) );
NOR2X1 NOR2X1_118 ( .A(_19_), .B(_20_), .Y(_26_) );
INVX1 INVX1_219 ( .A(_26_), .Y(_27_) );
AND2X2 AND2X2_93 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_28_) );
INVX1 INVX1_220 ( .A(_28_), .Y(_29_) );
NAND3X1 NAND3X1_109 ( .A(_27_), .B(_29_), .C(_25_), .Y(_30_) );
OAI21X1 OAI21X1_88 ( .A(i_add2[7]), .B(i_add1[7]), .C(_30_), .Y(_31_) );
INVX1 INVX1_221 ( .A(_31_), .Y(w_C_8_) );
INVX1 INVX1_222 ( .A(i_add2[8]), .Y(_32_) );
INVX1 INVX1_223 ( .A(i_add1[8]), .Y(_33_) );
NOR2X1 NOR2X1_119 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_34_) );
INVX1 INVX1_224 ( .A(_34_), .Y(_35_) );
BUFX2 BUFX2_57 ( .A(w_C_55_), .Y(_333__55_) );
BUFX2 BUFX2_58 ( .A(1'b0), .Y(w_C_0_) );
endmodule
