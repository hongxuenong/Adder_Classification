module cla_38bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [37:0] i_add1;
input [37:0] i_add2;
output [38:0] o_result;

OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_414_), .C(w_C_33_), .Y(_415_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_415_), .B(_419_), .Y(_209__33_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(w_C_34_), .Y(_423_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_424_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_425_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_425_), .C(_424_), .Y(_426_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_420_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_421_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_420_), .B(_421_), .C(w_C_34_), .Y(_422_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_422_), .B(_426_), .Y(_209__34_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(w_C_35_), .Y(_430_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_431_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_432_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_432_), .C(_431_), .Y(_433_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_427_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_428_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_427_), .B(_428_), .C(w_C_35_), .Y(_429_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(_433_), .Y(_209__35_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(w_C_36_), .Y(_437_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_438_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_439_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_439_), .C(_438_), .Y(_440_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_434_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_435_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_435_), .C(w_C_36_), .Y(_436_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_440_), .Y(_209__36_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(w_C_37_), .Y(_444_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_445_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_446_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_446_), .C(_445_), .Y(_447_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_441_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_442_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_442_), .C(w_C_37_), .Y(_443_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_447_), .Y(_209__37_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_451_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_452_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_453_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_453_), .C(_452_), .Y(_454_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_448_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_449_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_448_), .B(_449_), .C(gnd), .Y(_450_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_454_), .Y(_209__0_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_458_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_459_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_460_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_460_), .C(_459_), .Y(_461_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_455_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_456_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_456_), .C(w_C_1_), .Y(_457_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_461_), .Y(_209__1_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_465_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_466_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_467_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_467_), .C(_466_), .Y(_468_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_462_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_463_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_462_), .B(_463_), .C(w_C_2_), .Y(_464_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_468_), .Y(_209__2_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_472_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_473_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_474_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_474_), .C(_473_), .Y(_475_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_469_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_470_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_470_), .C(w_C_3_), .Y(_471_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_475_), .Y(_209__3_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_2_), .Y(w_C_2_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .Y(_3_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add1[2]), .Y(_4_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_2_), .C(_6_), .Y(_7_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_9_), .C(_7_), .Y(_10_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_10_), .Y(w_C_4_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(_12_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_13_), .C(_10_), .Y(_14_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_12_), .Y(w_C_5_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .Y(_15_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add1[5]), .Y(_16_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_17_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_17_), .Y(_18_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_18_), .C(_14_), .Y(_19_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_16_), .C(_19_), .Y(w_C_6_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_20_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_20_), .Y(_21_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_16_), .Y(_22_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_23_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_24_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_24_), .Y(_25_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_25_), .C(_19_), .Y(_26_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_21_), .Y(w_C_7_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_27_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(_28_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_29_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_29_), .Y(_30_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_30_), .C(_26_), .Y(_31_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_28_), .Y(_32_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_32_), .Y(w_C_8_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_33_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_33_), .Y(_34_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_35_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_32_), .C(_34_), .Y(w_C_9_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_36_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_36_), .Y(_37_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_35_), .Y(_38_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_34_), .C(_31_), .Y(_39_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_40_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_40_), .Y(_41_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_41_), .C(_39_), .Y(_42_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_37_), .Y(_43_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(w_C_10_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_44_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_44_), .Y(_45_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_46_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_43_), .C(_45_), .Y(w_C_11_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .Y(_47_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add1[11]), .Y(_48_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_46_), .Y(_49_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_45_), .C(_42_), .Y(_50_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_51_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_51_), .Y(_52_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_52_), .C(_50_), .Y(_53_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_48_), .C(_53_), .Y(w_C_12_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_48_), .Y(_54_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_54_), .Y(_55_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_56_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_56_), .Y(_57_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_57_), .C(_53_), .Y(_58_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .C(_58_), .Y(_59_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_59_), .Y(w_C_13_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .Y(_60_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add1[13]), .Y(_61_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_62_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_62_), .Y(_63_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_64_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_64_), .Y(_65_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_65_), .C(_58_), .Y(_66_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_61_), .C(_66_), .Y(w_C_14_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_61_), .Y(_67_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_67_), .Y(_68_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_69_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(_70_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_70_), .C(_66_), .Y(_71_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .C(_71_), .Y(_72_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_72_), .Y(w_C_15_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .Y(_73_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add1[15]), .Y(_74_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_75_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_75_), .Y(_76_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_77_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(_78_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_78_), .C(_71_), .Y(_79_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_74_), .C(_79_), .Y(w_C_16_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_74_), .Y(_80_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_80_), .Y(_81_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_82_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_82_), .Y(_83_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_83_), .C(_79_), .Y(_84_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .C(_84_), .Y(_85_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_85_), .Y(w_C_17_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .Y(_86_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add1[17]), .Y(_87_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_88_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_88_), .Y(_89_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_90_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_90_), .Y(_91_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_91_), .C(_84_), .Y(_92_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_87_), .C(_92_), .Y(w_C_18_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_87_), .Y(_93_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_93_), .Y(_94_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_95_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_95_), .Y(_96_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_96_), .C(_92_), .Y(_97_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .C(_97_), .Y(_98_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_98_), .Y(w_C_19_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .Y(_99_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add1[19]), .Y(_100_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_101_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_101_), .Y(_102_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_103_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_103_), .Y(_104_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_104_), .C(_97_), .Y(_105_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_100_), .C(_105_), .Y(w_C_20_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_100_), .Y(_106_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_106_), .Y(_107_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_108_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_108_), .Y(_109_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_109_), .C(_105_), .Y(_110_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .C(_110_), .Y(_111_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_111_), .Y(w_C_21_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .Y(_112_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add1[21]), .Y(_113_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_114_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_114_), .Y(_115_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_116_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_116_), .Y(_117_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_117_), .C(_110_), .Y(_118_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_113_), .C(_118_), .Y(w_C_22_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_113_), .Y(_119_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_119_), .Y(_120_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_121_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_121_), .Y(_122_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_122_), .C(_118_), .Y(_123_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .C(_123_), .Y(_124_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_124_), .Y(w_C_23_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .Y(_125_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add1[23]), .Y(_126_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_127_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_127_), .Y(_128_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_129_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(_129_), .Y(_130_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_130_), .C(_123_), .Y(_131_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_126_), .C(_131_), .Y(w_C_24_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_126_), .Y(_132_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_132_), .Y(_133_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_134_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_134_), .Y(_135_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_135_), .C(_131_), .Y(_136_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .C(_136_), .Y(_137_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_137_), .Y(w_C_25_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .Y(_138_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add1[25]), .Y(_139_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_140_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(_140_), .Y(_141_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_142_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_142_), .Y(_143_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_143_), .C(_136_), .Y(_144_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_139_), .C(_144_), .Y(w_C_26_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_139_), .Y(_145_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_145_), .Y(_146_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_147_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_147_), .Y(_148_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_148_), .C(_144_), .Y(_149_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .C(_149_), .Y(_150_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_150_), .Y(w_C_27_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .Y(_151_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add1[27]), .Y(_152_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_153_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_153_), .Y(_154_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_155_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(_156_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_156_), .C(_149_), .Y(_157_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_152_), .C(_157_), .Y(w_C_28_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_152_), .Y(_158_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(_158_), .Y(_159_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_160_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(_160_), .Y(_161_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_159_), .B(_161_), .C(_157_), .Y(_162_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .C(_162_), .Y(_163_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_163_), .Y(w_C_29_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .Y(_164_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add1[29]), .Y(_165_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_166_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(_166_), .Y(_167_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_168_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_168_), .Y(_169_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_169_), .C(_162_), .Y(_170_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_165_), .C(_170_), .Y(w_C_30_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_171_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_171_), .Y(_172_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_165_), .Y(_173_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(_173_), .Y(_174_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_175_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_175_), .C(_170_), .Y(_176_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_172_), .Y(w_C_31_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .Y(_177_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add1[31]), .Y(_178_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_178_), .Y(_179_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_179_), .C(_176_), .Y(_180_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_178_), .C(_180_), .Y(w_C_32_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .Y(_181_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add1[32]), .Y(_182_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_182_), .Y(_183_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_184_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_185_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_185_), .C(_180_), .Y(_186_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_183_), .Y(w_C_33_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .Y(_187_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add1[33]), .Y(_188_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(_188_), .Y(_189_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_189_), .C(_186_), .Y(_190_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(_188_), .C(_190_), .Y(w_C_34_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(_188_), .Y(_191_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_191_), .Y(_192_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_193_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(_193_), .Y(_194_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(_194_), .C(_190_), .Y(_195_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .C(_195_), .Y(_196_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_196_), .Y(w_C_35_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_197_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_198_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_196_), .C(_197_), .Y(w_C_36_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_199_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_200_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_200_), .Y(_201_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_198_), .Y(_202_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_202_), .C(_195_), .Y(_203_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_204_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_204_), .C(_203_), .Y(_205_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_199_), .Y(w_C_37_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_206_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_207_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_207_), .C(_205_), .Y(_208_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_208_), .Y(w_C_38_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_209__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_209__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_209__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_209__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_209__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_209__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_209__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_209__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_209__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_209__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_209__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_209__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_209__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_209__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_209__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_209__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_209__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_209__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_209__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_209__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_209__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_209__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_209__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_209__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_209__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_209__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_209__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_209__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_209__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_209__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_209__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_209__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_209__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_209__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_209__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_209__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_209__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_209__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(w_C_38_), .Y(o_result[38]) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_213_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_214_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_215_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_215_), .C(_214_), .Y(_216_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_210_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_211_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_210_), .B(_211_), .C(w_C_4_), .Y(_212_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_216_), .Y(_209__4_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_220_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_221_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_222_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_222_), .C(_221_), .Y(_223_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_217_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_218_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_218_), .C(w_C_5_), .Y(_219_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_223_), .Y(_209__5_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_227_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_228_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_229_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_229_), .C(_228_), .Y(_230_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_224_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_225_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_225_), .C(w_C_6_), .Y(_226_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_230_), .Y(_209__6_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_234_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_235_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_236_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_236_), .C(_235_), .Y(_237_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_231_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_232_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_232_), .C(w_C_7_), .Y(_233_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_237_), .Y(_209__7_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_241_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_242_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_243_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_243_), .C(_242_), .Y(_244_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_238_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_239_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_238_), .B(_239_), .C(w_C_8_), .Y(_240_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_244_), .Y(_209__8_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_248_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_249_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_250_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_250_), .C(_249_), .Y(_251_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_245_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_246_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_246_), .C(w_C_9_), .Y(_247_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_251_), .Y(_209__9_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_255_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_256_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_257_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_257_), .C(_256_), .Y(_258_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_252_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_253_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_253_), .C(w_C_10_), .Y(_254_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_258_), .Y(_209__10_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_262_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_263_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_264_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_264_), .C(_263_), .Y(_265_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_259_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_260_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_260_), .C(w_C_11_), .Y(_261_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_265_), .Y(_209__11_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(w_C_12_), .Y(_269_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_270_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_271_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_271_), .C(_270_), .Y(_272_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_266_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_267_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_267_), .C(w_C_12_), .Y(_268_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_272_), .Y(_209__12_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(w_C_13_), .Y(_276_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_277_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_278_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_278_), .C(_277_), .Y(_279_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_273_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_274_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_274_), .C(w_C_13_), .Y(_275_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_279_), .Y(_209__13_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(w_C_14_), .Y(_283_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_284_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_285_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_283_), .B(_285_), .C(_284_), .Y(_286_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_280_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_281_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_281_), .C(w_C_14_), .Y(_282_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_286_), .Y(_209__14_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(_290_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_291_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_292_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_292_), .C(_291_), .Y(_293_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_287_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_288_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_287_), .B(_288_), .C(w_C_15_), .Y(_289_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_293_), .Y(_209__15_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(w_C_16_), .Y(_297_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_298_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_299_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_299_), .C(_298_), .Y(_300_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_294_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_295_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_295_), .C(w_C_16_), .Y(_296_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_300_), .Y(_209__16_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(w_C_17_), .Y(_304_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_305_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_306_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_306_), .C(_305_), .Y(_307_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_301_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_302_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_302_), .C(w_C_17_), .Y(_303_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_307_), .Y(_209__17_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(w_C_18_), .Y(_311_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_312_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_313_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_313_), .C(_312_), .Y(_314_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_308_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_309_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_309_), .C(w_C_18_), .Y(_310_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_314_), .Y(_209__18_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(w_C_19_), .Y(_318_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_319_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_320_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_320_), .C(_319_), .Y(_321_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_315_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_316_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_316_), .C(w_C_19_), .Y(_317_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_321_), .Y(_209__19_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(w_C_20_), .Y(_325_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_326_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_327_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_327_), .C(_326_), .Y(_328_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_322_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_323_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_323_), .C(w_C_20_), .Y(_324_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_328_), .Y(_209__20_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(w_C_21_), .Y(_332_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_333_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_334_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_334_), .C(_333_), .Y(_335_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_329_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_330_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_330_), .C(w_C_21_), .Y(_331_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_335_), .Y(_209__21_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(w_C_22_), .Y(_339_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_340_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_341_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_341_), .C(_340_), .Y(_342_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_336_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_337_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_337_), .C(w_C_22_), .Y(_338_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_342_), .Y(_209__22_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(w_C_23_), .Y(_346_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_347_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_348_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_348_), .C(_347_), .Y(_349_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_343_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_344_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_344_), .C(w_C_23_), .Y(_345_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_349_), .Y(_209__23_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(w_C_24_), .Y(_353_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_354_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_355_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_355_), .C(_354_), .Y(_356_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_350_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_351_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_351_), .C(w_C_24_), .Y(_352_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_356_), .Y(_209__24_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(w_C_25_), .Y(_360_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_361_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_362_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_362_), .C(_361_), .Y(_363_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_357_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_358_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_358_), .C(w_C_25_), .Y(_359_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_363_), .Y(_209__25_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(w_C_26_), .Y(_367_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_368_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_369_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_369_), .C(_368_), .Y(_370_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_364_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_365_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_365_), .C(w_C_26_), .Y(_366_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_370_), .Y(_209__26_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(w_C_27_), .Y(_374_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_375_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_376_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_376_), .C(_375_), .Y(_377_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_371_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_372_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_372_), .C(w_C_27_), .Y(_373_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_373_), .B(_377_), .Y(_209__27_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(w_C_28_), .Y(_381_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_382_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_383_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_383_), .C(_382_), .Y(_384_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_378_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_379_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_379_), .C(w_C_28_), .Y(_380_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_384_), .Y(_209__28_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(w_C_29_), .Y(_388_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_389_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_390_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(_390_), .C(_389_), .Y(_391_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_385_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_386_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_385_), .B(_386_), .C(w_C_29_), .Y(_387_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_391_), .Y(_209__29_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(w_C_30_), .Y(_395_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_396_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_397_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_397_), .C(_396_), .Y(_398_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_392_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_393_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_392_), .B(_393_), .C(w_C_30_), .Y(_394_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_398_), .Y(_209__30_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(w_C_31_), .Y(_402_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_403_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_404_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_404_), .C(_403_), .Y(_405_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_399_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_400_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_400_), .C(w_C_31_), .Y(_401_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_405_), .Y(_209__31_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(w_C_32_), .Y(_409_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_410_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_411_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_411_), .C(_410_), .Y(_412_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_406_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_407_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_406_), .B(_407_), .C(w_C_32_), .Y(_408_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_412_), .Y(_209__32_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(w_C_33_), .Y(_416_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_417_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_418_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_418_), .C(_417_), .Y(_419_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_413_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_414_) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(w_C_38_), .Y(_209__38_) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
