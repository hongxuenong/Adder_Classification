module CSkipA_44bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output cout;

OAI21X1 OAI21X1_1 ( .A(_390_), .B(_387_), .C(_392_), .Y(_23__1_) );
INVX1 INVX1_1 ( .A(_23__1_), .Y(_397_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_398_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_399_) );
NAND3X1 NAND3X1_1 ( .A(_397_), .B(_399_), .C(_398_), .Y(_400_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_394_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_395_) );
OAI21X1 OAI21X1_2 ( .A(_394_), .B(_395_), .C(_23__1_), .Y(_396_) );
NAND2X1 NAND2X1_2 ( .A(_396_), .B(_400_), .Y(_0__33_) );
OAI21X1 OAI21X1_3 ( .A(_397_), .B(_394_), .C(_399_), .Y(_23__2_) );
INVX1 INVX1_2 ( .A(_23__2_), .Y(_404_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_405_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_406_) );
NAND3X1 NAND3X1_2 ( .A(_404_), .B(_406_), .C(_405_), .Y(_407_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_401_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_402_) );
OAI21X1 OAI21X1_4 ( .A(_401_), .B(_402_), .C(_23__2_), .Y(_403_) );
NAND2X1 NAND2X1_4 ( .A(_403_), .B(_407_), .Y(_0__34_) );
OAI21X1 OAI21X1_5 ( .A(_404_), .B(_401_), .C(_406_), .Y(_23__3_) );
INVX1 INVX1_3 ( .A(_23__3_), .Y(_411_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_412_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_413_) );
NAND3X1 NAND3X1_3 ( .A(_411_), .B(_413_), .C(_412_), .Y(_414_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_408_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_409_) );
OAI21X1 OAI21X1_6 ( .A(_408_), .B(_409_), .C(_23__3_), .Y(_410_) );
NAND2X1 NAND2X1_6 ( .A(_410_), .B(_414_), .Y(_0__35_) );
OAI21X1 OAI21X1_7 ( .A(_411_), .B(_408_), .C(_413_), .Y(_22_) );
INVX1 INVX1_4 ( .A(w_cout_8_), .Y(_418_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_419_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_420_) );
NAND3X1 NAND3X1_4 ( .A(_418_), .B(_420_), .C(_419_), .Y(_421_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_415_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_416_) );
OAI21X1 OAI21X1_8 ( .A(_415_), .B(_416_), .C(w_cout_8_), .Y(_417_) );
NAND2X1 NAND2X1_8 ( .A(_417_), .B(_421_), .Y(_0__36_) );
OAI21X1 OAI21X1_9 ( .A(_418_), .B(_415_), .C(_420_), .Y(_26__1_) );
INVX1 INVX1_5 ( .A(_26__1_), .Y(_425_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_426_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_427_) );
NAND3X1 NAND3X1_5 ( .A(_425_), .B(_427_), .C(_426_), .Y(_428_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_422_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_423_) );
OAI21X1 OAI21X1_10 ( .A(_422_), .B(_423_), .C(_26__1_), .Y(_424_) );
NAND2X1 NAND2X1_10 ( .A(_424_), .B(_428_), .Y(_0__37_) );
OAI21X1 OAI21X1_11 ( .A(_425_), .B(_422_), .C(_427_), .Y(_26__2_) );
INVX1 INVX1_6 ( .A(_26__2_), .Y(_432_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_433_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_434_) );
NAND3X1 NAND3X1_6 ( .A(_432_), .B(_434_), .C(_433_), .Y(_435_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_429_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_430_) );
OAI21X1 OAI21X1_12 ( .A(_429_), .B(_430_), .C(_26__2_), .Y(_431_) );
NAND2X1 NAND2X1_12 ( .A(_431_), .B(_435_), .Y(_0__38_) );
OAI21X1 OAI21X1_13 ( .A(_432_), .B(_429_), .C(_434_), .Y(_26__3_) );
INVX1 INVX1_7 ( .A(_26__3_), .Y(_439_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_440_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_441_) );
NAND3X1 NAND3X1_7 ( .A(_439_), .B(_441_), .C(_440_), .Y(_442_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_436_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_437_) );
OAI21X1 OAI21X1_14 ( .A(_436_), .B(_437_), .C(_26__3_), .Y(_438_) );
NAND2X1 NAND2X1_14 ( .A(_438_), .B(_442_), .Y(_0__39_) );
OAI21X1 OAI21X1_15 ( .A(_439_), .B(_436_), .C(_441_), .Y(_25_) );
INVX1 INVX1_8 ( .A(w_cout_9_), .Y(_446_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_447_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_448_) );
NAND3X1 NAND3X1_8 ( .A(_446_), .B(_448_), .C(_447_), .Y(_449_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_443_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_444_) );
OAI21X1 OAI21X1_16 ( .A(_443_), .B(_444_), .C(w_cout_9_), .Y(_445_) );
NAND2X1 NAND2X1_16 ( .A(_445_), .B(_449_), .Y(_0__40_) );
OAI21X1 OAI21X1_17 ( .A(_446_), .B(_443_), .C(_448_), .Y(_29__1_) );
INVX1 INVX1_9 ( .A(_29__1_), .Y(_453_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_454_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_455_) );
NAND3X1 NAND3X1_9 ( .A(_453_), .B(_455_), .C(_454_), .Y(_456_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_450_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_451_) );
OAI21X1 OAI21X1_18 ( .A(_450_), .B(_451_), .C(_29__1_), .Y(_452_) );
NAND2X1 NAND2X1_18 ( .A(_452_), .B(_456_), .Y(_0__41_) );
OAI21X1 OAI21X1_19 ( .A(_453_), .B(_450_), .C(_455_), .Y(_29__2_) );
INVX1 INVX1_10 ( .A(_29__2_), .Y(_460_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_461_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_462_) );
NAND3X1 NAND3X1_10 ( .A(_460_), .B(_462_), .C(_461_), .Y(_463_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_457_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_458_) );
OAI21X1 OAI21X1_20 ( .A(_457_), .B(_458_), .C(_29__2_), .Y(_459_) );
NAND2X1 NAND2X1_20 ( .A(_459_), .B(_463_), .Y(_0__42_) );
OAI21X1 OAI21X1_21 ( .A(_460_), .B(_457_), .C(_462_), .Y(_29__3_) );
INVX1 INVX1_11 ( .A(_29__3_), .Y(_467_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_468_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_469_) );
NAND3X1 NAND3X1_11 ( .A(_467_), .B(_469_), .C(_468_), .Y(_470_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_464_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_465_) );
OAI21X1 OAI21X1_22 ( .A(_464_), .B(_465_), .C(_29__3_), .Y(_466_) );
NAND2X1 NAND2X1_22 ( .A(_466_), .B(_470_), .Y(_0__43_) );
OAI21X1 OAI21X1_23 ( .A(_467_), .B(_464_), .C(_469_), .Y(_28_) );
INVX1 INVX1_12 ( .A(1'b0), .Y(_474_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_475_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_476_) );
NAND3X1 NAND3X1_12 ( .A(_474_), .B(_476_), .C(_475_), .Y(_477_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_471_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_472_) );
OAI21X1 OAI21X1_24 ( .A(_471_), .B(_472_), .C(1'b0), .Y(_473_) );
NAND2X1 NAND2X1_24 ( .A(_473_), .B(_477_), .Y(_0__0_) );
OAI21X1 OAI21X1_25 ( .A(_474_), .B(_471_), .C(_476_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_13 ( .A(rca_inst_w_CARRY_1_), .Y(_481_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_482_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_483_) );
NAND3X1 NAND3X1_13 ( .A(_481_), .B(_483_), .C(_482_), .Y(_484_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_478_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_479_) );
OAI21X1 OAI21X1_26 ( .A(_478_), .B(_479_), .C(rca_inst_w_CARRY_1_), .Y(_480_) );
NAND2X1 NAND2X1_26 ( .A(_480_), .B(_484_), .Y(_0__1_) );
OAI21X1 OAI21X1_27 ( .A(_481_), .B(_478_), .C(_483_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_14 ( .A(rca_inst_w_CARRY_2_), .Y(_488_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_489_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_490_) );
NAND3X1 NAND3X1_14 ( .A(_488_), .B(_490_), .C(_489_), .Y(_491_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_485_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_486_) );
OAI21X1 OAI21X1_28 ( .A(_485_), .B(_486_), .C(rca_inst_w_CARRY_2_), .Y(_487_) );
NAND2X1 NAND2X1_28 ( .A(_487_), .B(_491_), .Y(_0__2_) );
OAI21X1 OAI21X1_29 ( .A(_488_), .B(_485_), .C(_490_), .Y(rca_inst_w_CARRY_3_) );
INVX1 INVX1_15 ( .A(rca_inst_w_CARRY_3_), .Y(_495_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_496_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_497_) );
NAND3X1 NAND3X1_15 ( .A(_495_), .B(_497_), .C(_496_), .Y(_498_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_492_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_493_) );
OAI21X1 OAI21X1_30 ( .A(_492_), .B(_493_), .C(rca_inst_w_CARRY_3_), .Y(_494_) );
NAND2X1 NAND2X1_30 ( .A(_494_), .B(_498_), .Y(_0__3_) );
OAI21X1 OAI21X1_31 ( .A(_495_), .B(_492_), .C(_497_), .Y(cout0) );
INVX1 INVX1_16 ( .A(i_add_term1[0]), .Y(_499_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[0]), .B(_499_), .Y(_500_) );
INVX1 INVX1_17 ( .A(i_add_term2[0]), .Y(_501_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term1[0]), .B(_501_), .Y(_502_) );
INVX1 INVX1_18 ( .A(i_add_term1[1]), .Y(_503_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[1]), .B(_503_), .Y(_504_) );
INVX1 INVX1_19 ( .A(i_add_term2[1]), .Y(_505_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term1[1]), .B(_505_), .Y(_506_) );
OAI22X1 OAI22X1_1 ( .A(_500_), .B(_502_), .C(_504_), .D(_506_), .Y(_507_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_508_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_509_) );
NOR2X1 NOR2X1_21 ( .A(_508_), .B(_509_), .Y(_510_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_511_) );
NAND2X1 NAND2X1_31 ( .A(_510_), .B(_511_), .Y(_512_) );
NOR2X1 NOR2X1_22 ( .A(_507_), .B(_512_), .Y(skip0_P) );
INVX1 INVX1_20 ( .A(cout0), .Y(_513_) );
NAND2X1 NAND2X1_32 ( .A(1'b0), .B(skip0_P), .Y(_514_) );
OAI21X1 OAI21X1_32 ( .A(skip0_P), .B(_513_), .C(_514_), .Y(skip0_cin_next) );
BUFX2 BUFX2_1 ( .A(w_cout_10_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
INVX1 INVX1_21 ( .A(i_add_term1[4]), .Y(_31_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[4]), .B(_31_), .Y(_32_) );
INVX1 INVX1_22 ( .A(i_add_term2[4]), .Y(_33_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term1[4]), .B(_33_), .Y(_34_) );
INVX1 INVX1_23 ( .A(i_add_term1[5]), .Y(_35_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[5]), .B(_35_), .Y(_36_) );
INVX1 INVX1_24 ( .A(i_add_term2[5]), .Y(_37_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term1[5]), .B(_37_), .Y(_38_) );
OAI22X1 OAI22X1_2 ( .A(_32_), .B(_34_), .C(_36_), .D(_38_), .Y(_39_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_40_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_41_) );
NOR2X1 NOR2X1_28 ( .A(_40_), .B(_41_), .Y(_42_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_43_) );
NAND2X1 NAND2X1_33 ( .A(_42_), .B(_43_), .Y(_44_) );
NOR2X1 NOR2X1_29 ( .A(_39_), .B(_44_), .Y(_3_) );
INVX1 INVX1_25 ( .A(_1_), .Y(_45_) );
NAND2X1 NAND2X1_34 ( .A(1'b0), .B(_3_), .Y(_46_) );
OAI21X1 OAI21X1_33 ( .A(_3_), .B(_45_), .C(_46_), .Y(w_cout_1_) );
INVX1 INVX1_26 ( .A(i_add_term1[8]), .Y(_47_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[8]), .B(_47_), .Y(_48_) );
INVX1 INVX1_27 ( .A(i_add_term2[8]), .Y(_49_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term1[8]), .B(_49_), .Y(_50_) );
INVX1 INVX1_28 ( .A(i_add_term1[9]), .Y(_51_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[9]), .B(_51_), .Y(_52_) );
INVX1 INVX1_29 ( .A(i_add_term2[9]), .Y(_53_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term1[9]), .B(_53_), .Y(_54_) );
OAI22X1 OAI22X1_3 ( .A(_48_), .B(_50_), .C(_52_), .D(_54_), .Y(_55_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_56_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_57_) );
NOR2X1 NOR2X1_35 ( .A(_56_), .B(_57_), .Y(_58_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_59_) );
NAND2X1 NAND2X1_35 ( .A(_58_), .B(_59_), .Y(_60_) );
NOR2X1 NOR2X1_36 ( .A(_55_), .B(_60_), .Y(_6_) );
INVX1 INVX1_30 ( .A(_4_), .Y(_61_) );
NAND2X1 NAND2X1_36 ( .A(1'b0), .B(_6_), .Y(_62_) );
OAI21X1 OAI21X1_34 ( .A(_6_), .B(_61_), .C(_62_), .Y(w_cout_2_) );
INVX1 INVX1_31 ( .A(i_add_term1[12]), .Y(_63_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[12]), .B(_63_), .Y(_64_) );
INVX1 INVX1_32 ( .A(i_add_term2[12]), .Y(_65_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term1[12]), .B(_65_), .Y(_66_) );
INVX1 INVX1_33 ( .A(i_add_term1[13]), .Y(_67_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[13]), .B(_67_), .Y(_68_) );
INVX1 INVX1_34 ( .A(i_add_term2[13]), .Y(_69_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term1[13]), .B(_69_), .Y(_70_) );
OAI22X1 OAI22X1_4 ( .A(_64_), .B(_66_), .C(_68_), .D(_70_), .Y(_71_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_72_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_73_) );
NOR2X1 NOR2X1_42 ( .A(_72_), .B(_73_), .Y(_74_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_75_) );
NAND2X1 NAND2X1_37 ( .A(_74_), .B(_75_), .Y(_76_) );
NOR2X1 NOR2X1_43 ( .A(_71_), .B(_76_), .Y(_9_) );
INVX1 INVX1_35 ( .A(_7_), .Y(_77_) );
NAND2X1 NAND2X1_38 ( .A(1'b0), .B(_9_), .Y(_78_) );
OAI21X1 OAI21X1_35 ( .A(_9_), .B(_77_), .C(_78_), .Y(w_cout_3_) );
INVX1 INVX1_36 ( .A(i_add_term1[16]), .Y(_79_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[16]), .B(_79_), .Y(_80_) );
INVX1 INVX1_37 ( .A(i_add_term2[16]), .Y(_81_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term1[16]), .B(_81_), .Y(_82_) );
INVX1 INVX1_38 ( .A(i_add_term1[17]), .Y(_83_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[17]), .B(_83_), .Y(_84_) );
INVX1 INVX1_39 ( .A(i_add_term2[17]), .Y(_85_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term1[17]), .B(_85_), .Y(_86_) );
OAI22X1 OAI22X1_5 ( .A(_80_), .B(_82_), .C(_84_), .D(_86_), .Y(_87_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_88_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_89_) );
NOR2X1 NOR2X1_49 ( .A(_88_), .B(_89_), .Y(_90_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_91_) );
NAND2X1 NAND2X1_39 ( .A(_90_), .B(_91_), .Y(_92_) );
NOR2X1 NOR2X1_50 ( .A(_87_), .B(_92_), .Y(_12_) );
INVX1 INVX1_40 ( .A(_10_), .Y(_93_) );
NAND2X1 NAND2X1_40 ( .A(1'b0), .B(_12_), .Y(_94_) );
OAI21X1 OAI21X1_36 ( .A(_12_), .B(_93_), .C(_94_), .Y(w_cout_4_) );
INVX1 INVX1_41 ( .A(i_add_term1[20]), .Y(_95_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[20]), .B(_95_), .Y(_96_) );
INVX1 INVX1_42 ( .A(i_add_term2[20]), .Y(_97_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term1[20]), .B(_97_), .Y(_98_) );
INVX1 INVX1_43 ( .A(i_add_term1[21]), .Y(_99_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[21]), .B(_99_), .Y(_100_) );
INVX1 INVX1_44 ( .A(i_add_term2[21]), .Y(_101_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term1[21]), .B(_101_), .Y(_102_) );
OAI22X1 OAI22X1_6 ( .A(_96_), .B(_98_), .C(_100_), .D(_102_), .Y(_103_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_104_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_105_) );
NOR2X1 NOR2X1_56 ( .A(_104_), .B(_105_), .Y(_106_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_107_) );
NAND2X1 NAND2X1_41 ( .A(_106_), .B(_107_), .Y(_108_) );
NOR2X1 NOR2X1_57 ( .A(_103_), .B(_108_), .Y(_15_) );
INVX1 INVX1_45 ( .A(_13_), .Y(_109_) );
NAND2X1 NAND2X1_42 ( .A(1'b0), .B(_15_), .Y(_110_) );
OAI21X1 OAI21X1_37 ( .A(_15_), .B(_109_), .C(_110_), .Y(w_cout_5_) );
INVX1 INVX1_46 ( .A(i_add_term1[24]), .Y(_111_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[24]), .B(_111_), .Y(_112_) );
INVX1 INVX1_47 ( .A(i_add_term2[24]), .Y(_113_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term1[24]), .B(_113_), .Y(_114_) );
INVX1 INVX1_48 ( .A(i_add_term1[25]), .Y(_115_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[25]), .B(_115_), .Y(_116_) );
INVX1 INVX1_49 ( .A(i_add_term2[25]), .Y(_117_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term1[25]), .B(_117_), .Y(_118_) );
OAI22X1 OAI22X1_7 ( .A(_112_), .B(_114_), .C(_116_), .D(_118_), .Y(_119_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_120_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_121_) );
NOR2X1 NOR2X1_63 ( .A(_120_), .B(_121_), .Y(_122_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_123_) );
NAND2X1 NAND2X1_43 ( .A(_122_), .B(_123_), .Y(_124_) );
NOR2X1 NOR2X1_64 ( .A(_119_), .B(_124_), .Y(_18_) );
INVX1 INVX1_50 ( .A(_16_), .Y(_125_) );
NAND2X1 NAND2X1_44 ( .A(1'b0), .B(_18_), .Y(_126_) );
OAI21X1 OAI21X1_38 ( .A(_18_), .B(_125_), .C(_126_), .Y(w_cout_6_) );
INVX1 INVX1_51 ( .A(i_add_term1[28]), .Y(_127_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[28]), .B(_127_), .Y(_128_) );
INVX1 INVX1_52 ( .A(i_add_term2[28]), .Y(_129_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term1[28]), .B(_129_), .Y(_130_) );
INVX1 INVX1_53 ( .A(i_add_term1[29]), .Y(_131_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[29]), .B(_131_), .Y(_132_) );
INVX1 INVX1_54 ( .A(i_add_term2[29]), .Y(_133_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term1[29]), .B(_133_), .Y(_134_) );
OAI22X1 OAI22X1_8 ( .A(_128_), .B(_130_), .C(_132_), .D(_134_), .Y(_135_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_136_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_137_) );
NOR2X1 NOR2X1_70 ( .A(_136_), .B(_137_), .Y(_138_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_139_) );
NAND2X1 NAND2X1_45 ( .A(_138_), .B(_139_), .Y(_140_) );
NOR2X1 NOR2X1_71 ( .A(_135_), .B(_140_), .Y(_21_) );
INVX1 INVX1_55 ( .A(_19_), .Y(_141_) );
NAND2X1 NAND2X1_46 ( .A(1'b0), .B(_21_), .Y(_142_) );
OAI21X1 OAI21X1_39 ( .A(_21_), .B(_141_), .C(_142_), .Y(w_cout_7_) );
INVX1 INVX1_56 ( .A(i_add_term1[32]), .Y(_143_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[32]), .B(_143_), .Y(_144_) );
INVX1 INVX1_57 ( .A(i_add_term2[32]), .Y(_145_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term1[32]), .B(_145_), .Y(_146_) );
INVX1 INVX1_58 ( .A(i_add_term1[33]), .Y(_147_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[33]), .B(_147_), .Y(_148_) );
INVX1 INVX1_59 ( .A(i_add_term2[33]), .Y(_149_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term1[33]), .B(_149_), .Y(_150_) );
OAI22X1 OAI22X1_9 ( .A(_144_), .B(_146_), .C(_148_), .D(_150_), .Y(_151_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_152_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_153_) );
NOR2X1 NOR2X1_77 ( .A(_152_), .B(_153_), .Y(_154_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_155_) );
NAND2X1 NAND2X1_47 ( .A(_154_), .B(_155_), .Y(_156_) );
NOR2X1 NOR2X1_78 ( .A(_151_), .B(_156_), .Y(_24_) );
INVX1 INVX1_60 ( .A(_22_), .Y(_157_) );
NAND2X1 NAND2X1_48 ( .A(1'b0), .B(_24_), .Y(_158_) );
OAI21X1 OAI21X1_40 ( .A(_24_), .B(_157_), .C(_158_), .Y(w_cout_8_) );
INVX1 INVX1_61 ( .A(i_add_term1[36]), .Y(_159_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[36]), .B(_159_), .Y(_160_) );
INVX1 INVX1_62 ( .A(i_add_term2[36]), .Y(_161_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term1[36]), .B(_161_), .Y(_162_) );
INVX1 INVX1_63 ( .A(i_add_term1[37]), .Y(_163_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[37]), .B(_163_), .Y(_164_) );
INVX1 INVX1_64 ( .A(i_add_term2[37]), .Y(_165_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term1[37]), .B(_165_), .Y(_166_) );
OAI22X1 OAI22X1_10 ( .A(_160_), .B(_162_), .C(_164_), .D(_166_), .Y(_167_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_168_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_169_) );
NOR2X1 NOR2X1_84 ( .A(_168_), .B(_169_), .Y(_170_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_171_) );
NAND2X1 NAND2X1_49 ( .A(_170_), .B(_171_), .Y(_172_) );
NOR2X1 NOR2X1_85 ( .A(_167_), .B(_172_), .Y(_27_) );
INVX1 INVX1_65 ( .A(_25_), .Y(_173_) );
NAND2X1 NAND2X1_50 ( .A(1'b0), .B(_27_), .Y(_174_) );
OAI21X1 OAI21X1_41 ( .A(_27_), .B(_173_), .C(_174_), .Y(w_cout_9_) );
INVX1 INVX1_66 ( .A(i_add_term1[40]), .Y(_175_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[40]), .B(_175_), .Y(_176_) );
INVX1 INVX1_67 ( .A(i_add_term2[40]), .Y(_177_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term1[40]), .B(_177_), .Y(_178_) );
INVX1 INVX1_68 ( .A(i_add_term1[41]), .Y(_179_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[41]), .B(_179_), .Y(_180_) );
INVX1 INVX1_69 ( .A(i_add_term2[41]), .Y(_181_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term1[41]), .B(_181_), .Y(_182_) );
OAI22X1 OAI22X1_11 ( .A(_176_), .B(_178_), .C(_180_), .D(_182_), .Y(_183_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_184_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_185_) );
NOR2X1 NOR2X1_91 ( .A(_184_), .B(_185_), .Y(_186_) );
XOR2X1 XOR2X1_11 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_187_) );
NAND2X1 NAND2X1_51 ( .A(_186_), .B(_187_), .Y(_188_) );
NOR2X1 NOR2X1_92 ( .A(_183_), .B(_188_), .Y(_30_) );
INVX1 INVX1_70 ( .A(_28_), .Y(_189_) );
NAND2X1 NAND2X1_52 ( .A(1'b0), .B(_30_), .Y(_190_) );
OAI21X1 OAI21X1_42 ( .A(_30_), .B(_189_), .C(_190_), .Y(w_cout_10_) );
INVX1 INVX1_71 ( .A(skip0_cin_next), .Y(_194_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_195_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_196_) );
NAND3X1 NAND3X1_16 ( .A(_194_), .B(_196_), .C(_195_), .Y(_197_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_191_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_192_) );
OAI21X1 OAI21X1_43 ( .A(_191_), .B(_192_), .C(skip0_cin_next), .Y(_193_) );
NAND2X1 NAND2X1_54 ( .A(_193_), .B(_197_), .Y(_0__4_) );
OAI21X1 OAI21X1_44 ( .A(_194_), .B(_191_), .C(_196_), .Y(_2__1_) );
INVX1 INVX1_72 ( .A(_2__1_), .Y(_201_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_202_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_203_) );
NAND3X1 NAND3X1_17 ( .A(_201_), .B(_203_), .C(_202_), .Y(_204_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_198_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_199_) );
OAI21X1 OAI21X1_45 ( .A(_198_), .B(_199_), .C(_2__1_), .Y(_200_) );
NAND2X1 NAND2X1_56 ( .A(_200_), .B(_204_), .Y(_0__5_) );
OAI21X1 OAI21X1_46 ( .A(_201_), .B(_198_), .C(_203_), .Y(_2__2_) );
INVX1 INVX1_73 ( .A(_2__2_), .Y(_208_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_209_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_210_) );
NAND3X1 NAND3X1_18 ( .A(_208_), .B(_210_), .C(_209_), .Y(_211_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_205_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_206_) );
OAI21X1 OAI21X1_47 ( .A(_205_), .B(_206_), .C(_2__2_), .Y(_207_) );
NAND2X1 NAND2X1_58 ( .A(_207_), .B(_211_), .Y(_0__6_) );
OAI21X1 OAI21X1_48 ( .A(_208_), .B(_205_), .C(_210_), .Y(_2__3_) );
INVX1 INVX1_74 ( .A(_2__3_), .Y(_215_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_216_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_217_) );
NAND3X1 NAND3X1_19 ( .A(_215_), .B(_217_), .C(_216_), .Y(_218_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_212_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_213_) );
OAI21X1 OAI21X1_49 ( .A(_212_), .B(_213_), .C(_2__3_), .Y(_214_) );
NAND2X1 NAND2X1_60 ( .A(_214_), .B(_218_), .Y(_0__7_) );
OAI21X1 OAI21X1_50 ( .A(_215_), .B(_212_), .C(_217_), .Y(_1_) );
INVX1 INVX1_75 ( .A(w_cout_1_), .Y(_222_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_223_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_224_) );
NAND3X1 NAND3X1_20 ( .A(_222_), .B(_224_), .C(_223_), .Y(_225_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_219_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_220_) );
OAI21X1 OAI21X1_51 ( .A(_219_), .B(_220_), .C(w_cout_1_), .Y(_221_) );
NAND2X1 NAND2X1_62 ( .A(_221_), .B(_225_), .Y(_0__8_) );
OAI21X1 OAI21X1_52 ( .A(_222_), .B(_219_), .C(_224_), .Y(_5__1_) );
INVX1 INVX1_76 ( .A(_5__1_), .Y(_229_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_230_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_231_) );
NAND3X1 NAND3X1_21 ( .A(_229_), .B(_231_), .C(_230_), .Y(_232_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_226_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_227_) );
OAI21X1 OAI21X1_53 ( .A(_226_), .B(_227_), .C(_5__1_), .Y(_228_) );
NAND2X1 NAND2X1_64 ( .A(_228_), .B(_232_), .Y(_0__9_) );
OAI21X1 OAI21X1_54 ( .A(_229_), .B(_226_), .C(_231_), .Y(_5__2_) );
INVX1 INVX1_77 ( .A(_5__2_), .Y(_236_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_237_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_238_) );
NAND3X1 NAND3X1_22 ( .A(_236_), .B(_238_), .C(_237_), .Y(_239_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_233_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_234_) );
OAI21X1 OAI21X1_55 ( .A(_233_), .B(_234_), .C(_5__2_), .Y(_235_) );
NAND2X1 NAND2X1_66 ( .A(_235_), .B(_239_), .Y(_0__10_) );
OAI21X1 OAI21X1_56 ( .A(_236_), .B(_233_), .C(_238_), .Y(_5__3_) );
INVX1 INVX1_78 ( .A(_5__3_), .Y(_243_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_244_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_245_) );
NAND3X1 NAND3X1_23 ( .A(_243_), .B(_245_), .C(_244_), .Y(_246_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_240_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_241_) );
OAI21X1 OAI21X1_57 ( .A(_240_), .B(_241_), .C(_5__3_), .Y(_242_) );
NAND2X1 NAND2X1_68 ( .A(_242_), .B(_246_), .Y(_0__11_) );
OAI21X1 OAI21X1_58 ( .A(_243_), .B(_240_), .C(_245_), .Y(_4_) );
INVX1 INVX1_79 ( .A(w_cout_2_), .Y(_250_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_251_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_252_) );
NAND3X1 NAND3X1_24 ( .A(_250_), .B(_252_), .C(_251_), .Y(_253_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_247_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_248_) );
OAI21X1 OAI21X1_59 ( .A(_247_), .B(_248_), .C(w_cout_2_), .Y(_249_) );
NAND2X1 NAND2X1_70 ( .A(_249_), .B(_253_), .Y(_0__12_) );
OAI21X1 OAI21X1_60 ( .A(_250_), .B(_247_), .C(_252_), .Y(_8__1_) );
INVX1 INVX1_80 ( .A(_8__1_), .Y(_257_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_258_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_259_) );
NAND3X1 NAND3X1_25 ( .A(_257_), .B(_259_), .C(_258_), .Y(_260_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_254_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_255_) );
OAI21X1 OAI21X1_61 ( .A(_254_), .B(_255_), .C(_8__1_), .Y(_256_) );
NAND2X1 NAND2X1_72 ( .A(_256_), .B(_260_), .Y(_0__13_) );
OAI21X1 OAI21X1_62 ( .A(_257_), .B(_254_), .C(_259_), .Y(_8__2_) );
INVX1 INVX1_81 ( .A(_8__2_), .Y(_264_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_265_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_266_) );
NAND3X1 NAND3X1_26 ( .A(_264_), .B(_266_), .C(_265_), .Y(_267_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_261_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_262_) );
OAI21X1 OAI21X1_63 ( .A(_261_), .B(_262_), .C(_8__2_), .Y(_263_) );
NAND2X1 NAND2X1_74 ( .A(_263_), .B(_267_), .Y(_0__14_) );
OAI21X1 OAI21X1_64 ( .A(_264_), .B(_261_), .C(_266_), .Y(_8__3_) );
INVX1 INVX1_82 ( .A(_8__3_), .Y(_271_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_272_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_273_) );
NAND3X1 NAND3X1_27 ( .A(_271_), .B(_273_), .C(_272_), .Y(_274_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_268_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_269_) );
OAI21X1 OAI21X1_65 ( .A(_268_), .B(_269_), .C(_8__3_), .Y(_270_) );
NAND2X1 NAND2X1_76 ( .A(_270_), .B(_274_), .Y(_0__15_) );
OAI21X1 OAI21X1_66 ( .A(_271_), .B(_268_), .C(_273_), .Y(_7_) );
INVX1 INVX1_83 ( .A(w_cout_3_), .Y(_278_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_279_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_280_) );
NAND3X1 NAND3X1_28 ( .A(_278_), .B(_280_), .C(_279_), .Y(_281_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_275_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_276_) );
OAI21X1 OAI21X1_67 ( .A(_275_), .B(_276_), .C(w_cout_3_), .Y(_277_) );
NAND2X1 NAND2X1_78 ( .A(_277_), .B(_281_), .Y(_0__16_) );
OAI21X1 OAI21X1_68 ( .A(_278_), .B(_275_), .C(_280_), .Y(_11__1_) );
INVX1 INVX1_84 ( .A(_11__1_), .Y(_285_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_286_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_287_) );
NAND3X1 NAND3X1_29 ( .A(_285_), .B(_287_), .C(_286_), .Y(_288_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_282_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_283_) );
OAI21X1 OAI21X1_69 ( .A(_282_), .B(_283_), .C(_11__1_), .Y(_284_) );
NAND2X1 NAND2X1_80 ( .A(_284_), .B(_288_), .Y(_0__17_) );
OAI21X1 OAI21X1_70 ( .A(_285_), .B(_282_), .C(_287_), .Y(_11__2_) );
INVX1 INVX1_85 ( .A(_11__2_), .Y(_292_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_293_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_294_) );
NAND3X1 NAND3X1_30 ( .A(_292_), .B(_294_), .C(_293_), .Y(_295_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_289_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_290_) );
OAI21X1 OAI21X1_71 ( .A(_289_), .B(_290_), .C(_11__2_), .Y(_291_) );
NAND2X1 NAND2X1_82 ( .A(_291_), .B(_295_), .Y(_0__18_) );
OAI21X1 OAI21X1_72 ( .A(_292_), .B(_289_), .C(_294_), .Y(_11__3_) );
INVX1 INVX1_86 ( .A(_11__3_), .Y(_299_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_300_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_301_) );
NAND3X1 NAND3X1_31 ( .A(_299_), .B(_301_), .C(_300_), .Y(_302_) );
NOR2X1 NOR2X1_108 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_296_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_297_) );
OAI21X1 OAI21X1_73 ( .A(_296_), .B(_297_), .C(_11__3_), .Y(_298_) );
NAND2X1 NAND2X1_84 ( .A(_298_), .B(_302_), .Y(_0__19_) );
OAI21X1 OAI21X1_74 ( .A(_299_), .B(_296_), .C(_301_), .Y(_10_) );
INVX1 INVX1_87 ( .A(w_cout_4_), .Y(_306_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_307_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_308_) );
NAND3X1 NAND3X1_32 ( .A(_306_), .B(_308_), .C(_307_), .Y(_309_) );
NOR2X1 NOR2X1_109 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_303_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_304_) );
OAI21X1 OAI21X1_75 ( .A(_303_), .B(_304_), .C(w_cout_4_), .Y(_305_) );
NAND2X1 NAND2X1_86 ( .A(_305_), .B(_309_), .Y(_0__20_) );
OAI21X1 OAI21X1_76 ( .A(_306_), .B(_303_), .C(_308_), .Y(_14__1_) );
INVX1 INVX1_88 ( .A(_14__1_), .Y(_313_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_314_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_315_) );
NAND3X1 NAND3X1_33 ( .A(_313_), .B(_315_), .C(_314_), .Y(_316_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_310_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_311_) );
OAI21X1 OAI21X1_77 ( .A(_310_), .B(_311_), .C(_14__1_), .Y(_312_) );
NAND2X1 NAND2X1_88 ( .A(_312_), .B(_316_), .Y(_0__21_) );
OAI21X1 OAI21X1_78 ( .A(_313_), .B(_310_), .C(_315_), .Y(_14__2_) );
INVX1 INVX1_89 ( .A(_14__2_), .Y(_320_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_321_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_322_) );
NAND3X1 NAND3X1_34 ( .A(_320_), .B(_322_), .C(_321_), .Y(_323_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_317_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_318_) );
OAI21X1 OAI21X1_79 ( .A(_317_), .B(_318_), .C(_14__2_), .Y(_319_) );
NAND2X1 NAND2X1_90 ( .A(_319_), .B(_323_), .Y(_0__22_) );
OAI21X1 OAI21X1_80 ( .A(_320_), .B(_317_), .C(_322_), .Y(_14__3_) );
INVX1 INVX1_90 ( .A(_14__3_), .Y(_327_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_328_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_329_) );
NAND3X1 NAND3X1_35 ( .A(_327_), .B(_329_), .C(_328_), .Y(_330_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_324_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_325_) );
OAI21X1 OAI21X1_81 ( .A(_324_), .B(_325_), .C(_14__3_), .Y(_326_) );
NAND2X1 NAND2X1_92 ( .A(_326_), .B(_330_), .Y(_0__23_) );
OAI21X1 OAI21X1_82 ( .A(_327_), .B(_324_), .C(_329_), .Y(_13_) );
INVX1 INVX1_91 ( .A(w_cout_5_), .Y(_334_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_335_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_336_) );
NAND3X1 NAND3X1_36 ( .A(_334_), .B(_336_), .C(_335_), .Y(_337_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_331_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_332_) );
OAI21X1 OAI21X1_83 ( .A(_331_), .B(_332_), .C(w_cout_5_), .Y(_333_) );
NAND2X1 NAND2X1_94 ( .A(_333_), .B(_337_), .Y(_0__24_) );
OAI21X1 OAI21X1_84 ( .A(_334_), .B(_331_), .C(_336_), .Y(_17__1_) );
INVX1 INVX1_92 ( .A(_17__1_), .Y(_341_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_342_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_343_) );
NAND3X1 NAND3X1_37 ( .A(_341_), .B(_343_), .C(_342_), .Y(_344_) );
NOR2X1 NOR2X1_114 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_338_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_339_) );
OAI21X1 OAI21X1_85 ( .A(_338_), .B(_339_), .C(_17__1_), .Y(_340_) );
NAND2X1 NAND2X1_96 ( .A(_340_), .B(_344_), .Y(_0__25_) );
OAI21X1 OAI21X1_86 ( .A(_341_), .B(_338_), .C(_343_), .Y(_17__2_) );
INVX1 INVX1_93 ( .A(_17__2_), .Y(_348_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_349_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_350_) );
NAND3X1 NAND3X1_38 ( .A(_348_), .B(_350_), .C(_349_), .Y(_351_) );
NOR2X1 NOR2X1_115 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_345_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_346_) );
OAI21X1 OAI21X1_87 ( .A(_345_), .B(_346_), .C(_17__2_), .Y(_347_) );
NAND2X1 NAND2X1_98 ( .A(_347_), .B(_351_), .Y(_0__26_) );
OAI21X1 OAI21X1_88 ( .A(_348_), .B(_345_), .C(_350_), .Y(_17__3_) );
INVX1 INVX1_94 ( .A(_17__3_), .Y(_355_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_356_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_357_) );
NAND3X1 NAND3X1_39 ( .A(_355_), .B(_357_), .C(_356_), .Y(_358_) );
NOR2X1 NOR2X1_116 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_352_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_353_) );
OAI21X1 OAI21X1_89 ( .A(_352_), .B(_353_), .C(_17__3_), .Y(_354_) );
NAND2X1 NAND2X1_100 ( .A(_354_), .B(_358_), .Y(_0__27_) );
OAI21X1 OAI21X1_90 ( .A(_355_), .B(_352_), .C(_357_), .Y(_16_) );
INVX1 INVX1_95 ( .A(w_cout_6_), .Y(_362_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_363_) );
NAND2X1 NAND2X1_101 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_364_) );
NAND3X1 NAND3X1_40 ( .A(_362_), .B(_364_), .C(_363_), .Y(_365_) );
NOR2X1 NOR2X1_117 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_359_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_360_) );
OAI21X1 OAI21X1_91 ( .A(_359_), .B(_360_), .C(w_cout_6_), .Y(_361_) );
NAND2X1 NAND2X1_102 ( .A(_361_), .B(_365_), .Y(_0__28_) );
OAI21X1 OAI21X1_92 ( .A(_362_), .B(_359_), .C(_364_), .Y(_20__1_) );
INVX1 INVX1_96 ( .A(_20__1_), .Y(_369_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_370_) );
NAND2X1 NAND2X1_103 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_371_) );
NAND3X1 NAND3X1_41 ( .A(_369_), .B(_371_), .C(_370_), .Y(_372_) );
NOR2X1 NOR2X1_118 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_366_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_367_) );
OAI21X1 OAI21X1_93 ( .A(_366_), .B(_367_), .C(_20__1_), .Y(_368_) );
NAND2X1 NAND2X1_104 ( .A(_368_), .B(_372_), .Y(_0__29_) );
OAI21X1 OAI21X1_94 ( .A(_369_), .B(_366_), .C(_371_), .Y(_20__2_) );
INVX1 INVX1_97 ( .A(_20__2_), .Y(_376_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_377_) );
NAND2X1 NAND2X1_105 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_378_) );
NAND3X1 NAND3X1_42 ( .A(_376_), .B(_378_), .C(_377_), .Y(_379_) );
NOR2X1 NOR2X1_119 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_373_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_374_) );
OAI21X1 OAI21X1_95 ( .A(_373_), .B(_374_), .C(_20__2_), .Y(_375_) );
NAND2X1 NAND2X1_106 ( .A(_375_), .B(_379_), .Y(_0__30_) );
OAI21X1 OAI21X1_96 ( .A(_376_), .B(_373_), .C(_378_), .Y(_20__3_) );
INVX1 INVX1_98 ( .A(_20__3_), .Y(_383_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_384_) );
NAND2X1 NAND2X1_107 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_385_) );
NAND3X1 NAND3X1_43 ( .A(_383_), .B(_385_), .C(_384_), .Y(_386_) );
NOR2X1 NOR2X1_120 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_380_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_381_) );
OAI21X1 OAI21X1_97 ( .A(_380_), .B(_381_), .C(_20__3_), .Y(_382_) );
NAND2X1 NAND2X1_108 ( .A(_382_), .B(_386_), .Y(_0__31_) );
OAI21X1 OAI21X1_98 ( .A(_383_), .B(_380_), .C(_385_), .Y(_19_) );
INVX1 INVX1_99 ( .A(w_cout_7_), .Y(_390_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_391_) );
NAND2X1 NAND2X1_109 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_392_) );
NAND3X1 NAND3X1_44 ( .A(_390_), .B(_392_), .C(_391_), .Y(_393_) );
NOR2X1 NOR2X1_121 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_387_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_388_) );
OAI21X1 OAI21X1_99 ( .A(_387_), .B(_388_), .C(w_cout_7_), .Y(_389_) );
NAND2X1 NAND2X1_110 ( .A(_389_), .B(_393_), .Y(_0__32_) );
BUFX2 BUFX2_46 ( .A(skip0_cin_next), .Y(_2__0_) );
BUFX2 BUFX2_47 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_48 ( .A(w_cout_1_), .Y(_5__0_) );
BUFX2 BUFX2_49 ( .A(_4_), .Y(_5__4_) );
BUFX2 BUFX2_50 ( .A(w_cout_2_), .Y(_8__0_) );
BUFX2 BUFX2_51 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_52 ( .A(w_cout_3_), .Y(_11__0_) );
BUFX2 BUFX2_53 ( .A(_10_), .Y(_11__4_) );
BUFX2 BUFX2_54 ( .A(w_cout_4_), .Y(_14__0_) );
BUFX2 BUFX2_55 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_56 ( .A(w_cout_5_), .Y(_17__0_) );
BUFX2 BUFX2_57 ( .A(_16_), .Y(_17__4_) );
BUFX2 BUFX2_58 ( .A(w_cout_6_), .Y(_20__0_) );
BUFX2 BUFX2_59 ( .A(_19_), .Y(_20__4_) );
BUFX2 BUFX2_60 ( .A(w_cout_7_), .Y(_23__0_) );
BUFX2 BUFX2_61 ( .A(_22_), .Y(_23__4_) );
BUFX2 BUFX2_62 ( .A(w_cout_8_), .Y(_26__0_) );
BUFX2 BUFX2_63 ( .A(_25_), .Y(_26__4_) );
BUFX2 BUFX2_64 ( .A(w_cout_9_), .Y(_29__0_) );
BUFX2 BUFX2_65 ( .A(_28_), .Y(_29__4_) );
BUFX2 BUFX2_66 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_67 ( .A(cout0), .Y(rca_inst_w_CARRY_4_) );
BUFX2 BUFX2_68 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
