module CSkipA_57bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term1[45], i_add_term1[46], i_add_term1[47], i_add_term1[48], i_add_term1[49], i_add_term1[50], i_add_term1[51], i_add_term1[52], i_add_term1[53], i_add_term1[54], i_add_term1[55], i_add_term1[56], i_add_term1[57], i_add_term1[58], i_add_term1[59], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], i_add_term2[45], i_add_term2[46], i_add_term2[47], i_add_term2[48], i_add_term2[49], i_add_term2[50], i_add_term2[51], i_add_term2[52], i_add_term2[53], i_add_term2[54], i_add_term2[55], i_add_term2[56], i_add_term2[57], i_add_term2[58], i_add_term2[59], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], sum[45], sum[46], sum[47], sum[48], sum[49], sum[50], sum[51], sum[52], sum[53], sum[54], sum[55], sum[56], sum[57], sum[58], sum[59], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term1[45];
input i_add_term1[46];
input i_add_term1[47];
input i_add_term1[48];
input i_add_term1[49];
input i_add_term1[50];
input i_add_term1[51];
input i_add_term1[52];
input i_add_term1[53];
input i_add_term1[54];
input i_add_term1[55];
input i_add_term1[56];
input i_add_term1[57];
input i_add_term1[58];
input i_add_term1[59];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
input i_add_term2[45];
input i_add_term2[46];
input i_add_term2[47];
input i_add_term2[48];
input i_add_term2[49];
input i_add_term2[50];
input i_add_term2[51];
input i_add_term2[52];
input i_add_term2[53];
input i_add_term2[54];
input i_add_term2[55];
input i_add_term2[56];
input i_add_term2[57];
input i_add_term2[58];
input i_add_term2[59];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output sum[45];
output sum[46];
output sum[47];
output sum[48];
output sum[49];
output sum[50];
output sum[51];
output sum[52];
output sum[53];
output sum[54];
output sum[55];
output sum[56];
output sum[57];
output sum[58];
output sum[59];
output cout;

AND2X2 AND2X2_1 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_345_) );
OAI21X1 OAI21X1_1 ( .A(_344_), .B(_345_), .C(_18__1_), .Y(_346_) );
NAND2X1 NAND2X1_1 ( .A(_346_), .B(_350_), .Y(_0__37_) );
OAI21X1 OAI21X1_2 ( .A(_347_), .B(_344_), .C(_349_), .Y(_18__2_) );
INVX1 INVX1_1 ( .A(_18__2_), .Y(_354_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_355_) );
NAND2X1 NAND2X1_2 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_356_) );
NAND3X1 NAND3X1_1 ( .A(_354_), .B(_356_), .C(_355_), .Y(_357_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_351_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_352_) );
OAI21X1 OAI21X1_3 ( .A(_351_), .B(_352_), .C(_18__2_), .Y(_353_) );
NAND2X1 NAND2X1_3 ( .A(_353_), .B(_357_), .Y(_0__38_) );
OAI21X1 OAI21X1_4 ( .A(_354_), .B(_351_), .C(_356_), .Y(_18__3_) );
INVX1 INVX1_2 ( .A(_18__3_), .Y(_361_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_362_) );
NAND2X1 NAND2X1_4 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_363_) );
NAND3X1 NAND3X1_2 ( .A(_361_), .B(_363_), .C(_362_), .Y(_364_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_358_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_359_) );
OAI21X1 OAI21X1_5 ( .A(_358_), .B(_359_), .C(_18__3_), .Y(_360_) );
NAND2X1 NAND2X1_5 ( .A(_360_), .B(_364_), .Y(_0__39_) );
OAI21X1 OAI21X1_6 ( .A(_361_), .B(_358_), .C(_363_), .Y(_17_) );
INVX1 INVX1_3 ( .A(w_cout_9_), .Y(_368_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_369_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_370_) );
NAND3X1 NAND3X1_3 ( .A(_368_), .B(_370_), .C(_369_), .Y(_371_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_365_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_366_) );
OAI21X1 OAI21X1_7 ( .A(_365_), .B(_366_), .C(w_cout_9_), .Y(_367_) );
NAND2X1 NAND2X1_7 ( .A(_367_), .B(_371_), .Y(_0__40_) );
OAI21X1 OAI21X1_8 ( .A(_368_), .B(_365_), .C(_370_), .Y(_20__1_) );
INVX1 INVX1_4 ( .A(_20__1_), .Y(_375_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_376_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_377_) );
NAND3X1 NAND3X1_4 ( .A(_375_), .B(_377_), .C(_376_), .Y(_378_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_372_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_373_) );
OAI21X1 OAI21X1_9 ( .A(_372_), .B(_373_), .C(_20__1_), .Y(_374_) );
NAND2X1 NAND2X1_9 ( .A(_374_), .B(_378_), .Y(_0__41_) );
OAI21X1 OAI21X1_10 ( .A(_375_), .B(_372_), .C(_377_), .Y(_20__2_) );
INVX1 INVX1_5 ( .A(_20__2_), .Y(_382_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_383_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_384_) );
NAND3X1 NAND3X1_5 ( .A(_382_), .B(_384_), .C(_383_), .Y(_385_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_379_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_380_) );
OAI21X1 OAI21X1_11 ( .A(_379_), .B(_380_), .C(_20__2_), .Y(_381_) );
NAND2X1 NAND2X1_11 ( .A(_381_), .B(_385_), .Y(_0__42_) );
OAI21X1 OAI21X1_12 ( .A(_382_), .B(_379_), .C(_384_), .Y(_20__3_) );
INVX1 INVX1_6 ( .A(_20__3_), .Y(_389_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_390_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_391_) );
NAND3X1 NAND3X1_6 ( .A(_389_), .B(_391_), .C(_390_), .Y(_392_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_386_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_387_) );
OAI21X1 OAI21X1_13 ( .A(_386_), .B(_387_), .C(_20__3_), .Y(_388_) );
NAND2X1 NAND2X1_13 ( .A(_388_), .B(_392_), .Y(_0__43_) );
OAI21X1 OAI21X1_14 ( .A(_389_), .B(_386_), .C(_391_), .Y(_19_) );
INVX1 INVX1_7 ( .A(w_cout_10_), .Y(_396_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_397_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_398_) );
NAND3X1 NAND3X1_7 ( .A(_396_), .B(_398_), .C(_397_), .Y(_399_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_393_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_394_) );
OAI21X1 OAI21X1_15 ( .A(_393_), .B(_394_), .C(w_cout_10_), .Y(_395_) );
NAND2X1 NAND2X1_15 ( .A(_395_), .B(_399_), .Y(_0__44_) );
OAI21X1 OAI21X1_16 ( .A(_396_), .B(_393_), .C(_398_), .Y(_22__1_) );
INVX1 INVX1_8 ( .A(_22__1_), .Y(_403_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_404_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_405_) );
NAND3X1 NAND3X1_8 ( .A(_403_), .B(_405_), .C(_404_), .Y(_406_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_400_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_401_) );
OAI21X1 OAI21X1_17 ( .A(_400_), .B(_401_), .C(_22__1_), .Y(_402_) );
NAND2X1 NAND2X1_17 ( .A(_402_), .B(_406_), .Y(_0__45_) );
OAI21X1 OAI21X1_18 ( .A(_403_), .B(_400_), .C(_405_), .Y(_22__2_) );
INVX1 INVX1_9 ( .A(_22__2_), .Y(_410_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_411_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_412_) );
NAND3X1 NAND3X1_9 ( .A(_410_), .B(_412_), .C(_411_), .Y(_413_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_407_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_408_) );
OAI21X1 OAI21X1_19 ( .A(_407_), .B(_408_), .C(_22__2_), .Y(_409_) );
NAND2X1 NAND2X1_19 ( .A(_409_), .B(_413_), .Y(_0__46_) );
OAI21X1 OAI21X1_20 ( .A(_410_), .B(_407_), .C(_412_), .Y(_22__3_) );
INVX1 INVX1_10 ( .A(_22__3_), .Y(_417_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_418_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_419_) );
NAND3X1 NAND3X1_10 ( .A(_417_), .B(_419_), .C(_418_), .Y(_420_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_414_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_415_) );
OAI21X1 OAI21X1_21 ( .A(_414_), .B(_415_), .C(_22__3_), .Y(_416_) );
NAND2X1 NAND2X1_21 ( .A(_416_), .B(_420_), .Y(_0__47_) );
OAI21X1 OAI21X1_22 ( .A(_417_), .B(_414_), .C(_419_), .Y(_21_) );
INVX1 INVX1_11 ( .A(w_cout_11_), .Y(_424_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_425_) );
NAND2X1 NAND2X1_22 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_426_) );
NAND3X1 NAND3X1_11 ( .A(_424_), .B(_426_), .C(_425_), .Y(_427_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_421_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_422_) );
OAI21X1 OAI21X1_23 ( .A(_421_), .B(_422_), .C(w_cout_11_), .Y(_423_) );
NAND2X1 NAND2X1_23 ( .A(_423_), .B(_427_), .Y(_0__48_) );
OAI21X1 OAI21X1_24 ( .A(_424_), .B(_421_), .C(_426_), .Y(_24__1_) );
INVX1 INVX1_12 ( .A(_24__1_), .Y(_431_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_432_) );
NAND2X1 NAND2X1_24 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_433_) );
NAND3X1 NAND3X1_12 ( .A(_431_), .B(_433_), .C(_432_), .Y(_434_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_428_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_429_) );
OAI21X1 OAI21X1_25 ( .A(_428_), .B(_429_), .C(_24__1_), .Y(_430_) );
NAND2X1 NAND2X1_25 ( .A(_430_), .B(_434_), .Y(_0__49_) );
OAI21X1 OAI21X1_26 ( .A(_431_), .B(_428_), .C(_433_), .Y(_24__2_) );
INVX1 INVX1_13 ( .A(_24__2_), .Y(_438_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_439_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_440_) );
NAND3X1 NAND3X1_13 ( .A(_438_), .B(_440_), .C(_439_), .Y(_441_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_435_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_436_) );
OAI21X1 OAI21X1_27 ( .A(_435_), .B(_436_), .C(_24__2_), .Y(_437_) );
NAND2X1 NAND2X1_27 ( .A(_437_), .B(_441_), .Y(_0__50_) );
OAI21X1 OAI21X1_28 ( .A(_438_), .B(_435_), .C(_440_), .Y(_24__3_) );
INVX1 INVX1_14 ( .A(_24__3_), .Y(_445_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_446_) );
NAND2X1 NAND2X1_28 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_447_) );
NAND3X1 NAND3X1_14 ( .A(_445_), .B(_447_), .C(_446_), .Y(_448_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_442_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_443_) );
OAI21X1 OAI21X1_29 ( .A(_442_), .B(_443_), .C(_24__3_), .Y(_444_) );
NAND2X1 NAND2X1_29 ( .A(_444_), .B(_448_), .Y(_0__51_) );
OAI21X1 OAI21X1_30 ( .A(_445_), .B(_442_), .C(_447_), .Y(_23_) );
INVX1 INVX1_15 ( .A(w_cout_12_), .Y(_452_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_453_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_454_) );
NAND3X1 NAND3X1_15 ( .A(_452_), .B(_454_), .C(_453_), .Y(_455_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_449_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_450_) );
OAI21X1 OAI21X1_31 ( .A(_449_), .B(_450_), .C(w_cout_12_), .Y(_451_) );
NAND2X1 NAND2X1_31 ( .A(_451_), .B(_455_), .Y(_0__52_) );
OAI21X1 OAI21X1_32 ( .A(_452_), .B(_449_), .C(_454_), .Y(_26__1_) );
INVX1 INVX1_16 ( .A(_26__1_), .Y(_459_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_460_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_461_) );
NAND3X1 NAND3X1_16 ( .A(_459_), .B(_461_), .C(_460_), .Y(_462_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_456_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_457_) );
OAI21X1 OAI21X1_33 ( .A(_456_), .B(_457_), .C(_26__1_), .Y(_458_) );
NAND2X1 NAND2X1_33 ( .A(_458_), .B(_462_), .Y(_0__53_) );
OAI21X1 OAI21X1_34 ( .A(_459_), .B(_456_), .C(_461_), .Y(_26__2_) );
INVX1 INVX1_17 ( .A(_26__2_), .Y(_466_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_467_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_468_) );
NAND3X1 NAND3X1_17 ( .A(_466_), .B(_468_), .C(_467_), .Y(_469_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_463_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_464_) );
OAI21X1 OAI21X1_35 ( .A(_463_), .B(_464_), .C(_26__2_), .Y(_465_) );
NAND2X1 NAND2X1_35 ( .A(_465_), .B(_469_), .Y(_0__54_) );
OAI21X1 OAI21X1_36 ( .A(_466_), .B(_463_), .C(_468_), .Y(_26__3_) );
INVX1 INVX1_18 ( .A(_26__3_), .Y(_473_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_474_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_475_) );
NAND3X1 NAND3X1_18 ( .A(_473_), .B(_475_), .C(_474_), .Y(_476_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_470_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_471_) );
OAI21X1 OAI21X1_37 ( .A(_470_), .B(_471_), .C(_26__3_), .Y(_472_) );
NAND2X1 NAND2X1_37 ( .A(_472_), .B(_476_), .Y(_0__55_) );
OAI21X1 OAI21X1_38 ( .A(_473_), .B(_470_), .C(_475_), .Y(_25_) );
INVX1 INVX1_19 ( .A(w_cout_13_), .Y(_480_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_481_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_482_) );
NAND3X1 NAND3X1_19 ( .A(_480_), .B(_482_), .C(_481_), .Y(_483_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_477_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_478_) );
OAI21X1 OAI21X1_39 ( .A(_477_), .B(_478_), .C(w_cout_13_), .Y(_479_) );
NAND2X1 NAND2X1_39 ( .A(_479_), .B(_483_), .Y(_0__56_) );
OAI21X1 OAI21X1_40 ( .A(_480_), .B(_477_), .C(_482_), .Y(_28__1_) );
INVX1 INVX1_20 ( .A(_28__1_), .Y(_487_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_488_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_489_) );
NAND3X1 NAND3X1_20 ( .A(_487_), .B(_489_), .C(_488_), .Y(_490_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_484_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_485_) );
OAI21X1 OAI21X1_41 ( .A(_484_), .B(_485_), .C(_28__1_), .Y(_486_) );
NAND2X1 NAND2X1_41 ( .A(_486_), .B(_490_), .Y(_0__57_) );
OAI21X1 OAI21X1_42 ( .A(_487_), .B(_484_), .C(_489_), .Y(_28__2_) );
INVX1 INVX1_21 ( .A(_28__2_), .Y(_494_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_495_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_496_) );
NAND3X1 NAND3X1_21 ( .A(_494_), .B(_496_), .C(_495_), .Y(_497_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_491_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_492_) );
OAI21X1 OAI21X1_43 ( .A(_491_), .B(_492_), .C(_28__2_), .Y(_493_) );
NAND2X1 NAND2X1_43 ( .A(_493_), .B(_497_), .Y(_0__58_) );
OAI21X1 OAI21X1_44 ( .A(_494_), .B(_491_), .C(_496_), .Y(_28__3_) );
INVX1 INVX1_22 ( .A(_28__3_), .Y(_501_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_502_) );
NAND2X1 NAND2X1_44 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_503_) );
NAND3X1 NAND3X1_22 ( .A(_501_), .B(_503_), .C(_502_), .Y(_504_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_498_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_499_) );
OAI21X1 OAI21X1_45 ( .A(_498_), .B(_499_), .C(_28__3_), .Y(_500_) );
NAND2X1 NAND2X1_45 ( .A(_500_), .B(_504_), .Y(_0__59_) );
OAI21X1 OAI21X1_46 ( .A(_501_), .B(_498_), .C(_503_), .Y(_27_) );
INVX1 INVX1_23 ( .A(1'b0), .Y(_508_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_509_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_510_) );
NAND3X1 NAND3X1_23 ( .A(_508_), .B(_510_), .C(_509_), .Y(_511_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_505_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_506_) );
OAI21X1 OAI21X1_47 ( .A(_505_), .B(_506_), .C(1'b0), .Y(_507_) );
NAND2X1 NAND2X1_47 ( .A(_507_), .B(_511_), .Y(_0__0_) );
OAI21X1 OAI21X1_48 ( .A(_508_), .B(_505_), .C(_510_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_24 ( .A(rca_inst_w_CARRY_1_), .Y(_515_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_516_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_517_) );
NAND3X1 NAND3X1_24 ( .A(_515_), .B(_517_), .C(_516_), .Y(_518_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_512_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_513_) );
OAI21X1 OAI21X1_49 ( .A(_512_), .B(_513_), .C(rca_inst_w_CARRY_1_), .Y(_514_) );
NAND2X1 NAND2X1_49 ( .A(_514_), .B(_518_), .Y(_0__1_) );
OAI21X1 OAI21X1_50 ( .A(_515_), .B(_512_), .C(_517_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_25 ( .A(rca_inst_w_CARRY_2_), .Y(_522_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_523_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_524_) );
NAND3X1 NAND3X1_25 ( .A(_522_), .B(_524_), .C(_523_), .Y(_525_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_519_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_520_) );
OAI21X1 OAI21X1_51 ( .A(_519_), .B(_520_), .C(rca_inst_w_CARRY_2_), .Y(_521_) );
NAND2X1 NAND2X1_51 ( .A(_521_), .B(_525_), .Y(_0__2_) );
OAI21X1 OAI21X1_52 ( .A(_522_), .B(_519_), .C(_524_), .Y(rca_inst_w_CARRY_3_) );
INVX1 INVX1_26 ( .A(rca_inst_w_CARRY_3_), .Y(_529_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_530_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_531_) );
NAND3X1 NAND3X1_26 ( .A(_529_), .B(_531_), .C(_530_), .Y(_532_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_526_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_527_) );
OAI21X1 OAI21X1_53 ( .A(_526_), .B(_527_), .C(rca_inst_w_CARRY_3_), .Y(_528_) );
NAND2X1 NAND2X1_53 ( .A(_528_), .B(_532_), .Y(_0__3_) );
OAI21X1 OAI21X1_54 ( .A(_529_), .B(_526_), .C(_531_), .Y(cout0) );
INVX1 INVX1_27 ( .A(cout0), .Y(_533_) );
OAI21X1 OAI21X1_55 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .C(1'b0), .Y(_534_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_535_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_536_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_537_) );
NAND3X1 NAND3X1_27 ( .A(_535_), .B(_536_), .C(_537_), .Y(_538_) );
OAI21X1 OAI21X1_56 ( .A(_534_), .B(_538_), .C(_533_), .Y(skip0_cin_next) );
BUFX2 BUFX2_1 ( .A(w_cout_14_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .A(_0__54_), .Y(sum[54]) );
BUFX2 BUFX2_57 ( .A(_0__55_), .Y(sum[55]) );
BUFX2 BUFX2_58 ( .A(_0__56_), .Y(sum[56]) );
BUFX2 BUFX2_59 ( .A(_0__57_), .Y(sum[57]) );
BUFX2 BUFX2_60 ( .A(_0__58_), .Y(sum[58]) );
BUFX2 BUFX2_61 ( .A(_0__59_), .Y(sum[59]) );
INVX1 INVX1_28 ( .A(_1_), .Y(_29_) );
OAI21X1 OAI21X1_57 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .C(1'b0), .Y(_30_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_31_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_32_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_33_) );
NAND3X1 NAND3X1_28 ( .A(_31_), .B(_32_), .C(_33_), .Y(_34_) );
OAI21X1 OAI21X1_58 ( .A(_30_), .B(_34_), .C(_29_), .Y(w_cout_1_) );
INVX1 INVX1_29 ( .A(_3_), .Y(_35_) );
OAI21X1 OAI21X1_59 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .C(1'b0), .Y(_36_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_37_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_38_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_39_) );
NAND3X1 NAND3X1_29 ( .A(_37_), .B(_38_), .C(_39_), .Y(_40_) );
OAI21X1 OAI21X1_60 ( .A(_36_), .B(_40_), .C(_35_), .Y(w_cout_2_) );
INVX1 INVX1_30 ( .A(_5_), .Y(_41_) );
OAI21X1 OAI21X1_61 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .C(1'b0), .Y(_42_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_43_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_44_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_45_) );
NAND3X1 NAND3X1_30 ( .A(_43_), .B(_44_), .C(_45_), .Y(_46_) );
OAI21X1 OAI21X1_62 ( .A(_42_), .B(_46_), .C(_41_), .Y(w_cout_3_) );
INVX1 INVX1_31 ( .A(_7_), .Y(_47_) );
OAI21X1 OAI21X1_63 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .C(1'b0), .Y(_48_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_49_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_50_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_51_) );
NAND3X1 NAND3X1_31 ( .A(_49_), .B(_50_), .C(_51_), .Y(_52_) );
OAI21X1 OAI21X1_64 ( .A(_48_), .B(_52_), .C(_47_), .Y(w_cout_4_) );
INVX1 INVX1_32 ( .A(_9_), .Y(_53_) );
OAI21X1 OAI21X1_65 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .C(1'b0), .Y(_54_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_55_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_56_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_57_) );
NAND3X1 NAND3X1_32 ( .A(_55_), .B(_56_), .C(_57_), .Y(_58_) );
OAI21X1 OAI21X1_66 ( .A(_54_), .B(_58_), .C(_53_), .Y(w_cout_5_) );
INVX1 INVX1_33 ( .A(_11_), .Y(_59_) );
OAI21X1 OAI21X1_67 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .C(1'b0), .Y(_60_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_61_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_62_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_63_) );
NAND3X1 NAND3X1_33 ( .A(_61_), .B(_62_), .C(_63_), .Y(_64_) );
OAI21X1 OAI21X1_68 ( .A(_60_), .B(_64_), .C(_59_), .Y(w_cout_6_) );
INVX1 INVX1_34 ( .A(_13_), .Y(_65_) );
OAI21X1 OAI21X1_69 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .C(1'b0), .Y(_66_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_67_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_68_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_69_) );
NAND3X1 NAND3X1_34 ( .A(_67_), .B(_68_), .C(_69_), .Y(_70_) );
OAI21X1 OAI21X1_70 ( .A(_66_), .B(_70_), .C(_65_), .Y(w_cout_7_) );
INVX1 INVX1_35 ( .A(_15_), .Y(_71_) );
OAI21X1 OAI21X1_71 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .C(1'b0), .Y(_72_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_73_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_74_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_75_) );
NAND3X1 NAND3X1_35 ( .A(_73_), .B(_74_), .C(_75_), .Y(_76_) );
OAI21X1 OAI21X1_72 ( .A(_72_), .B(_76_), .C(_71_), .Y(w_cout_8_) );
INVX1 INVX1_36 ( .A(_17_), .Y(_77_) );
OAI21X1 OAI21X1_73 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .C(1'b0), .Y(_78_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_79_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_80_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_81_) );
NAND3X1 NAND3X1_36 ( .A(_79_), .B(_80_), .C(_81_), .Y(_82_) );
OAI21X1 OAI21X1_74 ( .A(_78_), .B(_82_), .C(_77_), .Y(w_cout_9_) );
INVX1 INVX1_37 ( .A(_19_), .Y(_83_) );
OAI21X1 OAI21X1_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .C(1'b0), .Y(_84_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_85_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_86_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_87_) );
NAND3X1 NAND3X1_37 ( .A(_85_), .B(_86_), .C(_87_), .Y(_88_) );
OAI21X1 OAI21X1_76 ( .A(_84_), .B(_88_), .C(_83_), .Y(w_cout_10_) );
INVX1 INVX1_38 ( .A(_21_), .Y(_89_) );
OAI21X1 OAI21X1_77 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .C(1'b0), .Y(_90_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_91_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_92_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_93_) );
NAND3X1 NAND3X1_38 ( .A(_91_), .B(_92_), .C(_93_), .Y(_94_) );
OAI21X1 OAI21X1_78 ( .A(_90_), .B(_94_), .C(_89_), .Y(w_cout_11_) );
INVX1 INVX1_39 ( .A(_23_), .Y(_95_) );
OAI21X1 OAI21X1_79 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .C(1'b0), .Y(_96_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_97_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_98_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_99_) );
NAND3X1 NAND3X1_39 ( .A(_97_), .B(_98_), .C(_99_), .Y(_100_) );
OAI21X1 OAI21X1_80 ( .A(_96_), .B(_100_), .C(_95_), .Y(w_cout_12_) );
INVX1 INVX1_40 ( .A(_25_), .Y(_101_) );
OAI21X1 OAI21X1_81 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .C(1'b0), .Y(_102_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_103_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_104_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_105_) );
NAND3X1 NAND3X1_40 ( .A(_103_), .B(_104_), .C(_105_), .Y(_106_) );
OAI21X1 OAI21X1_82 ( .A(_102_), .B(_106_), .C(_101_), .Y(w_cout_13_) );
INVX1 INVX1_41 ( .A(_27_), .Y(_107_) );
OAI21X1 OAI21X1_83 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .C(1'b0), .Y(_108_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_109_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_110_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_111_) );
NAND3X1 NAND3X1_41 ( .A(_109_), .B(_110_), .C(_111_), .Y(_112_) );
OAI21X1 OAI21X1_84 ( .A(_108_), .B(_112_), .C(_107_), .Y(w_cout_14_) );
INVX1 INVX1_42 ( .A(skip0_cin_next), .Y(_116_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_117_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_118_) );
NAND3X1 NAND3X1_42 ( .A(_116_), .B(_118_), .C(_117_), .Y(_119_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_113_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_114_) );
OAI21X1 OAI21X1_85 ( .A(_113_), .B(_114_), .C(skip0_cin_next), .Y(_115_) );
NAND2X1 NAND2X1_55 ( .A(_115_), .B(_119_), .Y(_0__4_) );
OAI21X1 OAI21X1_86 ( .A(_116_), .B(_113_), .C(_118_), .Y(_2__1_) );
INVX1 INVX1_43 ( .A(_2__1_), .Y(_123_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_124_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_125_) );
NAND3X1 NAND3X1_43 ( .A(_123_), .B(_125_), .C(_124_), .Y(_126_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_120_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_121_) );
OAI21X1 OAI21X1_87 ( .A(_120_), .B(_121_), .C(_2__1_), .Y(_122_) );
NAND2X1 NAND2X1_57 ( .A(_122_), .B(_126_), .Y(_0__5_) );
OAI21X1 OAI21X1_88 ( .A(_123_), .B(_120_), .C(_125_), .Y(_2__2_) );
INVX1 INVX1_44 ( .A(_2__2_), .Y(_130_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_131_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_132_) );
NAND3X1 NAND3X1_44 ( .A(_130_), .B(_132_), .C(_131_), .Y(_133_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_127_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_128_) );
OAI21X1 OAI21X1_89 ( .A(_127_), .B(_128_), .C(_2__2_), .Y(_129_) );
NAND2X1 NAND2X1_59 ( .A(_129_), .B(_133_), .Y(_0__6_) );
OAI21X1 OAI21X1_90 ( .A(_130_), .B(_127_), .C(_132_), .Y(_2__3_) );
INVX1 INVX1_45 ( .A(_2__3_), .Y(_137_) );
OR2X2 OR2X2_75 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_138_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_139_) );
NAND3X1 NAND3X1_45 ( .A(_137_), .B(_139_), .C(_138_), .Y(_140_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_134_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_135_) );
OAI21X1 OAI21X1_91 ( .A(_134_), .B(_135_), .C(_2__3_), .Y(_136_) );
NAND2X1 NAND2X1_61 ( .A(_136_), .B(_140_), .Y(_0__7_) );
OAI21X1 OAI21X1_92 ( .A(_137_), .B(_134_), .C(_139_), .Y(_1_) );
INVX1 INVX1_46 ( .A(w_cout_1_), .Y(_144_) );
OR2X2 OR2X2_76 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_145_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_146_) );
NAND3X1 NAND3X1_46 ( .A(_144_), .B(_146_), .C(_145_), .Y(_147_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_141_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_142_) );
OAI21X1 OAI21X1_93 ( .A(_141_), .B(_142_), .C(w_cout_1_), .Y(_143_) );
NAND2X1 NAND2X1_63 ( .A(_143_), .B(_147_), .Y(_0__8_) );
OAI21X1 OAI21X1_94 ( .A(_144_), .B(_141_), .C(_146_), .Y(_4__1_) );
INVX1 INVX1_47 ( .A(_4__1_), .Y(_151_) );
OR2X2 OR2X2_77 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_152_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_153_) );
NAND3X1 NAND3X1_47 ( .A(_151_), .B(_153_), .C(_152_), .Y(_154_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_148_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_149_) );
OAI21X1 OAI21X1_95 ( .A(_148_), .B(_149_), .C(_4__1_), .Y(_150_) );
NAND2X1 NAND2X1_65 ( .A(_150_), .B(_154_), .Y(_0__9_) );
OAI21X1 OAI21X1_96 ( .A(_151_), .B(_148_), .C(_153_), .Y(_4__2_) );
INVX1 INVX1_48 ( .A(_4__2_), .Y(_158_) );
OR2X2 OR2X2_78 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_159_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_160_) );
NAND3X1 NAND3X1_48 ( .A(_158_), .B(_160_), .C(_159_), .Y(_161_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_155_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_156_) );
OAI21X1 OAI21X1_97 ( .A(_155_), .B(_156_), .C(_4__2_), .Y(_157_) );
NAND2X1 NAND2X1_67 ( .A(_157_), .B(_161_), .Y(_0__10_) );
OAI21X1 OAI21X1_98 ( .A(_158_), .B(_155_), .C(_160_), .Y(_4__3_) );
INVX1 INVX1_49 ( .A(_4__3_), .Y(_165_) );
OR2X2 OR2X2_79 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_166_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_167_) );
NAND3X1 NAND3X1_49 ( .A(_165_), .B(_167_), .C(_166_), .Y(_168_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_162_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_163_) );
OAI21X1 OAI21X1_99 ( .A(_162_), .B(_163_), .C(_4__3_), .Y(_164_) );
NAND2X1 NAND2X1_69 ( .A(_164_), .B(_168_), .Y(_0__11_) );
OAI21X1 OAI21X1_100 ( .A(_165_), .B(_162_), .C(_167_), .Y(_3_) );
INVX1 INVX1_50 ( .A(w_cout_2_), .Y(_172_) );
OR2X2 OR2X2_80 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_173_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_174_) );
NAND3X1 NAND3X1_50 ( .A(_172_), .B(_174_), .C(_173_), .Y(_175_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_169_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_170_) );
OAI21X1 OAI21X1_101 ( .A(_169_), .B(_170_), .C(w_cout_2_), .Y(_171_) );
NAND2X1 NAND2X1_71 ( .A(_171_), .B(_175_), .Y(_0__12_) );
OAI21X1 OAI21X1_102 ( .A(_172_), .B(_169_), .C(_174_), .Y(_6__1_) );
INVX1 INVX1_51 ( .A(_6__1_), .Y(_179_) );
OR2X2 OR2X2_81 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_180_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_181_) );
NAND3X1 NAND3X1_51 ( .A(_179_), .B(_181_), .C(_180_), .Y(_182_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_176_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_177_) );
OAI21X1 OAI21X1_103 ( .A(_176_), .B(_177_), .C(_6__1_), .Y(_178_) );
NAND2X1 NAND2X1_73 ( .A(_178_), .B(_182_), .Y(_0__13_) );
OAI21X1 OAI21X1_104 ( .A(_179_), .B(_176_), .C(_181_), .Y(_6__2_) );
INVX1 INVX1_52 ( .A(_6__2_), .Y(_186_) );
OR2X2 OR2X2_82 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_187_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_188_) );
NAND3X1 NAND3X1_52 ( .A(_186_), .B(_188_), .C(_187_), .Y(_189_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_183_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_184_) );
OAI21X1 OAI21X1_105 ( .A(_183_), .B(_184_), .C(_6__2_), .Y(_185_) );
NAND2X1 NAND2X1_75 ( .A(_185_), .B(_189_), .Y(_0__14_) );
OAI21X1 OAI21X1_106 ( .A(_186_), .B(_183_), .C(_188_), .Y(_6__3_) );
INVX1 INVX1_53 ( .A(_6__3_), .Y(_193_) );
OR2X2 OR2X2_83 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_194_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_195_) );
NAND3X1 NAND3X1_53 ( .A(_193_), .B(_195_), .C(_194_), .Y(_196_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_190_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_191_) );
OAI21X1 OAI21X1_107 ( .A(_190_), .B(_191_), .C(_6__3_), .Y(_192_) );
NAND2X1 NAND2X1_77 ( .A(_192_), .B(_196_), .Y(_0__15_) );
OAI21X1 OAI21X1_108 ( .A(_193_), .B(_190_), .C(_195_), .Y(_5_) );
INVX1 INVX1_54 ( .A(w_cout_3_), .Y(_200_) );
OR2X2 OR2X2_84 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_201_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_202_) );
NAND3X1 NAND3X1_54 ( .A(_200_), .B(_202_), .C(_201_), .Y(_203_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_197_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_198_) );
OAI21X1 OAI21X1_109 ( .A(_197_), .B(_198_), .C(w_cout_3_), .Y(_199_) );
NAND2X1 NAND2X1_79 ( .A(_199_), .B(_203_), .Y(_0__16_) );
OAI21X1 OAI21X1_110 ( .A(_200_), .B(_197_), .C(_202_), .Y(_8__1_) );
INVX1 INVX1_55 ( .A(_8__1_), .Y(_207_) );
OR2X2 OR2X2_85 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_208_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_209_) );
NAND3X1 NAND3X1_55 ( .A(_207_), .B(_209_), .C(_208_), .Y(_210_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_204_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_205_) );
OAI21X1 OAI21X1_111 ( .A(_204_), .B(_205_), .C(_8__1_), .Y(_206_) );
NAND2X1 NAND2X1_81 ( .A(_206_), .B(_210_), .Y(_0__17_) );
OAI21X1 OAI21X1_112 ( .A(_207_), .B(_204_), .C(_209_), .Y(_8__2_) );
INVX1 INVX1_56 ( .A(_8__2_), .Y(_214_) );
OR2X2 OR2X2_86 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_215_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_216_) );
NAND3X1 NAND3X1_56 ( .A(_214_), .B(_216_), .C(_215_), .Y(_217_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_211_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_212_) );
OAI21X1 OAI21X1_113 ( .A(_211_), .B(_212_), .C(_8__2_), .Y(_213_) );
NAND2X1 NAND2X1_83 ( .A(_213_), .B(_217_), .Y(_0__18_) );
OAI21X1 OAI21X1_114 ( .A(_214_), .B(_211_), .C(_216_), .Y(_8__3_) );
INVX1 INVX1_57 ( .A(_8__3_), .Y(_221_) );
OR2X2 OR2X2_87 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_222_) );
NAND2X1 NAND2X1_84 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_223_) );
NAND3X1 NAND3X1_57 ( .A(_221_), .B(_223_), .C(_222_), .Y(_224_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_218_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_219_) );
OAI21X1 OAI21X1_115 ( .A(_218_), .B(_219_), .C(_8__3_), .Y(_220_) );
NAND2X1 NAND2X1_85 ( .A(_220_), .B(_224_), .Y(_0__19_) );
OAI21X1 OAI21X1_116 ( .A(_221_), .B(_218_), .C(_223_), .Y(_7_) );
INVX1 INVX1_58 ( .A(w_cout_4_), .Y(_228_) );
OR2X2 OR2X2_88 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_229_) );
NAND2X1 NAND2X1_86 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_230_) );
NAND3X1 NAND3X1_58 ( .A(_228_), .B(_230_), .C(_229_), .Y(_231_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_225_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_226_) );
OAI21X1 OAI21X1_117 ( .A(_225_), .B(_226_), .C(w_cout_4_), .Y(_227_) );
NAND2X1 NAND2X1_87 ( .A(_227_), .B(_231_), .Y(_0__20_) );
OAI21X1 OAI21X1_118 ( .A(_228_), .B(_225_), .C(_230_), .Y(_10__1_) );
INVX1 INVX1_59 ( .A(_10__1_), .Y(_235_) );
OR2X2 OR2X2_89 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_236_) );
NAND2X1 NAND2X1_88 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_237_) );
NAND3X1 NAND3X1_59 ( .A(_235_), .B(_237_), .C(_236_), .Y(_238_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_232_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_233_) );
OAI21X1 OAI21X1_119 ( .A(_232_), .B(_233_), .C(_10__1_), .Y(_234_) );
NAND2X1 NAND2X1_89 ( .A(_234_), .B(_238_), .Y(_0__21_) );
OAI21X1 OAI21X1_120 ( .A(_235_), .B(_232_), .C(_237_), .Y(_10__2_) );
INVX1 INVX1_60 ( .A(_10__2_), .Y(_242_) );
OR2X2 OR2X2_90 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_243_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_244_) );
NAND3X1 NAND3X1_60 ( .A(_242_), .B(_244_), .C(_243_), .Y(_245_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_239_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_240_) );
OAI21X1 OAI21X1_121 ( .A(_239_), .B(_240_), .C(_10__2_), .Y(_241_) );
NAND2X1 NAND2X1_91 ( .A(_241_), .B(_245_), .Y(_0__22_) );
OAI21X1 OAI21X1_122 ( .A(_242_), .B(_239_), .C(_244_), .Y(_10__3_) );
INVX1 INVX1_61 ( .A(_10__3_), .Y(_249_) );
OR2X2 OR2X2_91 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_250_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_251_) );
NAND3X1 NAND3X1_61 ( .A(_249_), .B(_251_), .C(_250_), .Y(_252_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_246_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_247_) );
OAI21X1 OAI21X1_123 ( .A(_246_), .B(_247_), .C(_10__3_), .Y(_248_) );
NAND2X1 NAND2X1_93 ( .A(_248_), .B(_252_), .Y(_0__23_) );
OAI21X1 OAI21X1_124 ( .A(_249_), .B(_246_), .C(_251_), .Y(_9_) );
INVX1 INVX1_62 ( .A(w_cout_5_), .Y(_256_) );
OR2X2 OR2X2_92 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_257_) );
NAND2X1 NAND2X1_94 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_258_) );
NAND3X1 NAND3X1_62 ( .A(_256_), .B(_258_), .C(_257_), .Y(_259_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_253_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_254_) );
OAI21X1 OAI21X1_125 ( .A(_253_), .B(_254_), .C(w_cout_5_), .Y(_255_) );
NAND2X1 NAND2X1_95 ( .A(_255_), .B(_259_), .Y(_0__24_) );
OAI21X1 OAI21X1_126 ( .A(_256_), .B(_253_), .C(_258_), .Y(_12__1_) );
INVX1 INVX1_63 ( .A(_12__1_), .Y(_263_) );
OR2X2 OR2X2_93 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_264_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_265_) );
NAND3X1 NAND3X1_63 ( .A(_263_), .B(_265_), .C(_264_), .Y(_266_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_260_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_261_) );
OAI21X1 OAI21X1_127 ( .A(_260_), .B(_261_), .C(_12__1_), .Y(_262_) );
NAND2X1 NAND2X1_97 ( .A(_262_), .B(_266_), .Y(_0__25_) );
OAI21X1 OAI21X1_128 ( .A(_263_), .B(_260_), .C(_265_), .Y(_12__2_) );
INVX1 INVX1_64 ( .A(_12__2_), .Y(_270_) );
OR2X2 OR2X2_94 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_271_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_272_) );
NAND3X1 NAND3X1_64 ( .A(_270_), .B(_272_), .C(_271_), .Y(_273_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_267_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_268_) );
OAI21X1 OAI21X1_129 ( .A(_267_), .B(_268_), .C(_12__2_), .Y(_269_) );
NAND2X1 NAND2X1_99 ( .A(_269_), .B(_273_), .Y(_0__26_) );
OAI21X1 OAI21X1_130 ( .A(_270_), .B(_267_), .C(_272_), .Y(_12__3_) );
INVX1 INVX1_65 ( .A(_12__3_), .Y(_277_) );
OR2X2 OR2X2_95 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_278_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_279_) );
NAND3X1 NAND3X1_65 ( .A(_277_), .B(_279_), .C(_278_), .Y(_280_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_274_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_275_) );
OAI21X1 OAI21X1_131 ( .A(_274_), .B(_275_), .C(_12__3_), .Y(_276_) );
NAND2X1 NAND2X1_101 ( .A(_276_), .B(_280_), .Y(_0__27_) );
OAI21X1 OAI21X1_132 ( .A(_277_), .B(_274_), .C(_279_), .Y(_11_) );
INVX1 INVX1_66 ( .A(w_cout_6_), .Y(_284_) );
OR2X2 OR2X2_96 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_285_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_286_) );
NAND3X1 NAND3X1_66 ( .A(_284_), .B(_286_), .C(_285_), .Y(_287_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_281_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_282_) );
OAI21X1 OAI21X1_133 ( .A(_281_), .B(_282_), .C(w_cout_6_), .Y(_283_) );
NAND2X1 NAND2X1_103 ( .A(_283_), .B(_287_), .Y(_0__28_) );
OAI21X1 OAI21X1_134 ( .A(_284_), .B(_281_), .C(_286_), .Y(_14__1_) );
INVX1 INVX1_67 ( .A(_14__1_), .Y(_291_) );
OR2X2 OR2X2_97 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_292_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_293_) );
NAND3X1 NAND3X1_67 ( .A(_291_), .B(_293_), .C(_292_), .Y(_294_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_288_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_289_) );
OAI21X1 OAI21X1_135 ( .A(_288_), .B(_289_), .C(_14__1_), .Y(_290_) );
NAND2X1 NAND2X1_105 ( .A(_290_), .B(_294_), .Y(_0__29_) );
OAI21X1 OAI21X1_136 ( .A(_291_), .B(_288_), .C(_293_), .Y(_14__2_) );
INVX1 INVX1_68 ( .A(_14__2_), .Y(_298_) );
OR2X2 OR2X2_98 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_299_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_300_) );
NAND3X1 NAND3X1_68 ( .A(_298_), .B(_300_), .C(_299_), .Y(_301_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_295_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_296_) );
OAI21X1 OAI21X1_137 ( .A(_295_), .B(_296_), .C(_14__2_), .Y(_297_) );
NAND2X1 NAND2X1_107 ( .A(_297_), .B(_301_), .Y(_0__30_) );
OAI21X1 OAI21X1_138 ( .A(_298_), .B(_295_), .C(_300_), .Y(_14__3_) );
INVX1 INVX1_69 ( .A(_14__3_), .Y(_305_) );
OR2X2 OR2X2_99 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_306_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_307_) );
NAND3X1 NAND3X1_69 ( .A(_305_), .B(_307_), .C(_306_), .Y(_308_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_302_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_303_) );
OAI21X1 OAI21X1_139 ( .A(_302_), .B(_303_), .C(_14__3_), .Y(_304_) );
NAND2X1 NAND2X1_109 ( .A(_304_), .B(_308_), .Y(_0__31_) );
OAI21X1 OAI21X1_140 ( .A(_305_), .B(_302_), .C(_307_), .Y(_13_) );
INVX1 INVX1_70 ( .A(w_cout_7_), .Y(_312_) );
OR2X2 OR2X2_100 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_313_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_314_) );
NAND3X1 NAND3X1_70 ( .A(_312_), .B(_314_), .C(_313_), .Y(_315_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_309_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_310_) );
OAI21X1 OAI21X1_141 ( .A(_309_), .B(_310_), .C(w_cout_7_), .Y(_311_) );
NAND2X1 NAND2X1_111 ( .A(_311_), .B(_315_), .Y(_0__32_) );
OAI21X1 OAI21X1_142 ( .A(_312_), .B(_309_), .C(_314_), .Y(_16__1_) );
INVX1 INVX1_71 ( .A(_16__1_), .Y(_319_) );
OR2X2 OR2X2_101 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_320_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_321_) );
NAND3X1 NAND3X1_71 ( .A(_319_), .B(_321_), .C(_320_), .Y(_322_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_316_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_317_) );
OAI21X1 OAI21X1_143 ( .A(_316_), .B(_317_), .C(_16__1_), .Y(_318_) );
NAND2X1 NAND2X1_113 ( .A(_318_), .B(_322_), .Y(_0__33_) );
OAI21X1 OAI21X1_144 ( .A(_319_), .B(_316_), .C(_321_), .Y(_16__2_) );
INVX1 INVX1_72 ( .A(_16__2_), .Y(_326_) );
OR2X2 OR2X2_102 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_327_) );
NAND2X1 NAND2X1_114 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_328_) );
NAND3X1 NAND3X1_72 ( .A(_326_), .B(_328_), .C(_327_), .Y(_329_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_323_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_324_) );
OAI21X1 OAI21X1_145 ( .A(_323_), .B(_324_), .C(_16__2_), .Y(_325_) );
NAND2X1 NAND2X1_115 ( .A(_325_), .B(_329_), .Y(_0__34_) );
OAI21X1 OAI21X1_146 ( .A(_326_), .B(_323_), .C(_328_), .Y(_16__3_) );
INVX1 INVX1_73 ( .A(_16__3_), .Y(_333_) );
OR2X2 OR2X2_103 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_334_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_335_) );
NAND3X1 NAND3X1_73 ( .A(_333_), .B(_335_), .C(_334_), .Y(_336_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_330_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_331_) );
OAI21X1 OAI21X1_147 ( .A(_330_), .B(_331_), .C(_16__3_), .Y(_332_) );
NAND2X1 NAND2X1_117 ( .A(_332_), .B(_336_), .Y(_0__35_) );
OAI21X1 OAI21X1_148 ( .A(_333_), .B(_330_), .C(_335_), .Y(_15_) );
INVX1 INVX1_74 ( .A(w_cout_8_), .Y(_340_) );
OR2X2 OR2X2_104 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_341_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_342_) );
NAND3X1 NAND3X1_74 ( .A(_340_), .B(_342_), .C(_341_), .Y(_343_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_337_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_338_) );
OAI21X1 OAI21X1_149 ( .A(_337_), .B(_338_), .C(w_cout_8_), .Y(_339_) );
NAND2X1 NAND2X1_119 ( .A(_339_), .B(_343_), .Y(_0__36_) );
OAI21X1 OAI21X1_150 ( .A(_340_), .B(_337_), .C(_342_), .Y(_18__1_) );
INVX1 INVX1_75 ( .A(_18__1_), .Y(_347_) );
OR2X2 OR2X2_105 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_348_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_349_) );
NAND3X1 NAND3X1_75 ( .A(_347_), .B(_349_), .C(_348_), .Y(_350_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_344_) );
BUFX2 BUFX2_62 ( .A(skip0_cin_next), .Y(_2__0_) );
BUFX2 BUFX2_63 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_64 ( .A(w_cout_1_), .Y(_4__0_) );
BUFX2 BUFX2_65 ( .A(_3_), .Y(_4__4_) );
BUFX2 BUFX2_66 ( .A(w_cout_2_), .Y(_6__0_) );
BUFX2 BUFX2_67 ( .A(_5_), .Y(_6__4_) );
BUFX2 BUFX2_68 ( .A(w_cout_3_), .Y(_8__0_) );
BUFX2 BUFX2_69 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_70 ( .A(w_cout_4_), .Y(_10__0_) );
BUFX2 BUFX2_71 ( .A(_9_), .Y(_10__4_) );
BUFX2 BUFX2_72 ( .A(w_cout_5_), .Y(_12__0_) );
BUFX2 BUFX2_73 ( .A(_11_), .Y(_12__4_) );
BUFX2 BUFX2_74 ( .A(w_cout_6_), .Y(_14__0_) );
BUFX2 BUFX2_75 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_76 ( .A(w_cout_7_), .Y(_16__0_) );
BUFX2 BUFX2_77 ( .A(_15_), .Y(_16__4_) );
BUFX2 BUFX2_78 ( .A(w_cout_8_), .Y(_18__0_) );
BUFX2 BUFX2_79 ( .A(_17_), .Y(_18__4_) );
BUFX2 BUFX2_80 ( .A(w_cout_9_), .Y(_20__0_) );
BUFX2 BUFX2_81 ( .A(_19_), .Y(_20__4_) );
BUFX2 BUFX2_82 ( .A(w_cout_10_), .Y(_22__0_) );
BUFX2 BUFX2_83 ( .A(_21_), .Y(_22__4_) );
BUFX2 BUFX2_84 ( .A(w_cout_11_), .Y(_24__0_) );
BUFX2 BUFX2_85 ( .A(_23_), .Y(_24__4_) );
BUFX2 BUFX2_86 ( .A(w_cout_12_), .Y(_26__0_) );
BUFX2 BUFX2_87 ( .A(_25_), .Y(_26__4_) );
BUFX2 BUFX2_88 ( .A(w_cout_13_), .Y(_28__0_) );
BUFX2 BUFX2_89 ( .A(_27_), .Y(_28__4_) );
BUFX2 BUFX2_90 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_91 ( .A(cout0), .Y(rca_inst_w_CARRY_4_) );
BUFX2 BUFX2_92 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
