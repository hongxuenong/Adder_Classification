module CSkipA_24bit ( gnd, vdd, i_add_term1, i_add_term2, sum, cout);

input gnd, vdd;
output cout;
input [23:0] i_add_term1;
input [23:0] i_add_term2;
output [23:0] sum;

BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .Y(cout) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_0__23_), .Y(sum[23]) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(skip0_cin_next), .Y(_19_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_20_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_21_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_21_), .C(_20_), .Y(_22_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_16_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_17_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_17_), .C(skip0_cin_next), .Y(_18_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_22_), .Y(_0__4_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_16_), .C(_21_), .Y(_2__1_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_2__3_), .Y(_26_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_27_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_28_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_28_), .C(_27_), .Y(_29_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_23_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_24_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_24_), .C(_2__3_), .Y(_25_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_29_), .Y(_0__7_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_23_), .C(_28_), .Y(_1_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_2__1_), .Y(_33_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_34_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_35_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_35_), .C(_34_), .Y(_36_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_30_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_31_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_31_), .C(_2__1_), .Y(_32_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_36_), .Y(_0__5_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_30_), .C(_35_), .Y(_2__2_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_2__2_), .Y(_40_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_41_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_42_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_42_), .C(_41_), .Y(_43_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_37_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_38_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_38_), .C(_2__2_), .Y(_39_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_43_), .Y(_0__6_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_37_), .C(_42_), .Y(_2__3_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .Y(_44_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[4]), .B(_44_), .Y(_45_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[4]), .Y(_46_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(_46_), .Y(_47_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[5]), .Y(_48_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(_48_), .Y(_49_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .Y(_50_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[5]), .B(_50_), .Y(_51_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_47_), .C(_49_), .D(_51_), .Y(_52_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_53_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_54_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_54_), .Y(_55_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_56_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_56_), .Y(_57_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_57_), .Y(_3_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_58_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_3_), .Y(_59_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_58_), .C(_59_), .Y(w_cout_1_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .Y(_63_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_64_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_65_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_65_), .C(_64_), .Y(_66_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_60_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_61_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_61_), .C(w_cout_1_), .Y(_62_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_66_), .Y(_0__8_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_60_), .C(_65_), .Y(_5__1_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_5__3_), .Y(_70_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_71_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_72_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_72_), .C(_71_), .Y(_73_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_67_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_68_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_68_), .C(_5__3_), .Y(_69_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_73_), .Y(_0__11_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_67_), .C(_72_), .Y(_4_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_5__1_), .Y(_77_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_78_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_79_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_79_), .C(_78_), .Y(_80_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_74_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_75_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_75_), .C(_5__1_), .Y(_76_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_80_), .Y(_0__9_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_74_), .C(_79_), .Y(_5__2_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_5__2_), .Y(_84_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_85_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_86_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_86_), .C(_85_), .Y(_87_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_81_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_82_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_82_), .C(_5__2_), .Y(_83_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_87_), .Y(_0__10_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_81_), .C(_86_), .Y(_5__3_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .Y(_88_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[8]), .B(_88_), .Y(_89_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[8]), .Y(_90_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(_90_), .Y(_91_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[9]), .Y(_92_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(_92_), .Y(_93_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .Y(_94_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[9]), .B(_94_), .Y(_95_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_91_), .C(_93_), .D(_95_), .Y(_96_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_97_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_98_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_98_), .Y(_99_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_100_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_100_), .Y(_101_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_101_), .Y(_6_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(_102_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_6_), .Y(_103_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_102_), .C(_103_), .Y(w_cout_2_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .Y(_107_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_108_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_109_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_109_), .C(_108_), .Y(_110_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_104_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_105_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_105_), .C(w_cout_2_), .Y(_106_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_106_), .B(_110_), .Y(_0__12_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_104_), .C(_109_), .Y(_8__1_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_8__3_), .Y(_114_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_115_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_116_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_116_), .C(_115_), .Y(_117_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_111_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_112_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_112_), .C(_8__3_), .Y(_113_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_117_), .Y(_0__15_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_111_), .C(_116_), .Y(_7_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_8__1_), .Y(_121_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_122_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_123_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_123_), .C(_122_), .Y(_124_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_118_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_119_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_119_), .C(_8__1_), .Y(_120_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_124_), .Y(_0__13_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_118_), .C(_123_), .Y(_8__2_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_8__2_), .Y(_128_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_129_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_130_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_130_), .C(_129_), .Y(_131_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_125_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_126_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_126_), .C(_8__2_), .Y(_127_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_131_), .Y(_0__14_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_125_), .C(_130_), .Y(_8__3_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .Y(_132_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[12]), .B(_132_), .Y(_133_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[12]), .Y(_134_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(_134_), .Y(_135_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[13]), .Y(_136_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(_136_), .Y(_137_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .Y(_138_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[13]), .B(_138_), .Y(_139_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_135_), .C(_137_), .D(_139_), .Y(_140_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_141_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_142_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_142_), .Y(_143_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_144_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_144_), .Y(_145_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_145_), .Y(_9_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_146_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_9_), .Y(_147_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_146_), .C(_147_), .Y(w_cout_3_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .Y(_151_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_152_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_153_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_153_), .C(_152_), .Y(_154_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_148_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_149_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_149_), .C(w_cout_3_), .Y(_150_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_154_), .Y(_0__16_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_148_), .C(_153_), .Y(_11__1_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_11__3_), .Y(_158_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_159_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_160_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_160_), .C(_159_), .Y(_161_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_155_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_156_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_156_), .C(_11__3_), .Y(_157_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_161_), .Y(_0__19_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_155_), .C(_160_), .Y(_10_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_11__1_), .Y(_165_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_166_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_167_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_167_), .C(_166_), .Y(_168_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_162_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_163_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_163_), .C(_11__1_), .Y(_164_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_168_), .Y(_0__17_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_162_), .C(_167_), .Y(_11__2_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_11__2_), .Y(_172_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_173_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_174_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_174_), .C(_173_), .Y(_175_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_169_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_170_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_170_), .C(_11__2_), .Y(_171_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_175_), .Y(_0__18_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_169_), .C(_174_), .Y(_11__3_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .Y(_176_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[16]), .B(_176_), .Y(_177_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[16]), .Y(_178_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(_178_), .Y(_179_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[17]), .Y(_180_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(_180_), .Y(_181_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .Y(_182_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[17]), .B(_182_), .Y(_183_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_179_), .C(_181_), .D(_183_), .Y(_184_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_185_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_186_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_186_), .Y(_187_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_188_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(_188_), .Y(_189_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_189_), .Y(_12_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(_190_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_12_), .Y(_191_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_190_), .C(_191_), .Y(w_cout_4_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .Y(_195_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_196_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_197_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_197_), .C(_196_), .Y(_198_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_192_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_193_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(_193_), .C(w_cout_4_), .Y(_194_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_198_), .Y(_0__20_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_192_), .C(_197_), .Y(_14__1_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_14__3_), .Y(_202_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_203_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_204_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_204_), .C(_203_), .Y(_205_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_199_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_200_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_200_), .C(_14__3_), .Y(_201_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_205_), .Y(_0__23_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_199_), .C(_204_), .Y(_13_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_14__1_), .Y(_209_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_210_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_211_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_211_), .C(_210_), .Y(_212_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_206_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_207_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_207_), .C(_14__1_), .Y(_208_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_212_), .Y(_0__21_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_206_), .C(_211_), .Y(_14__2_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_14__2_), .Y(_216_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_217_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_218_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_218_), .C(_217_), .Y(_219_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_213_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_214_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_214_), .C(_14__2_), .Y(_215_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_219_), .Y(_0__22_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_213_), .C(_218_), .Y(_14__3_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .Y(_220_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[20]), .B(_220_), .Y(_221_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[20]), .Y(_222_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(_222_), .Y(_223_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[21]), .Y(_224_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(_224_), .Y(_225_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .Y(_226_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[21]), .B(_226_), .Y(_227_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_223_), .C(_225_), .D(_227_), .Y(_228_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_229_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_230_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_230_), .Y(_231_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_232_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_232_), .Y(_233_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_233_), .Y(_15_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_234_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_15_), .Y(_235_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_234_), .C(_235_), .Y(w_cout_5_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_239_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_240_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_241_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_241_), .C(_240_), .Y(_242_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_236_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_237_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_237_), .C(gnd), .Y(_238_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_238_), .B(_242_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_236_), .C(_241_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_i_carry), .Y(_246_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_247_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_248_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_248_), .C(_247_), .Y(_249_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_243_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_244_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_244_), .C(rca_inst_fa3_i_carry), .Y(_245_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_249_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_243_), .C(_248_), .Y(cout0) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_carry), .Y(_253_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_254_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_255_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_253_), .B(_255_), .C(_254_), .Y(_256_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_250_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_251_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_251_), .C(rca_inst_fa0_o_carry), .Y(_252_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_256_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_253_), .B(_250_), .C(_255_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_carry), .Y(_260_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_261_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_262_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_262_), .C(_261_), .Y(_263_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_257_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_258_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_258_), .C(rca_inst_fa_1__o_carry), .Y(_259_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_263_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_257_), .C(_262_), .Y(rca_inst_fa3_i_carry) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .Y(_264_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .B(_264_), .Y(_265_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .Y(_266_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(_266_), .Y(_267_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .Y(_268_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(_268_), .Y(_269_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .Y(_270_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .B(_270_), .Y(_271_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_267_), .C(_269_), .D(_271_), .Y(_272_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_273_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_274_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_274_), .Y(_275_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_276_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_276_), .Y(_277_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_277_), .Y(skip0_P) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(cout0), .Y(_278_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(skip0_P), .Y(_279_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(skip0_P), .B(_278_), .C(_279_), .Y(skip0_cin_next) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
