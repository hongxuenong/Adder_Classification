module csa_40bit ( gnd, vdd, i_add_term1, i_add_term2, sum, cout);

input gnd, vdd;
output cout;
input [39:0] i_add_term1;
input [39:0] i_add_term2;
output [39:0] sum;

OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_264_), .C(gnd), .Y(_265_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_269_), .Y(_21__0_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_263_), .C(_268_), .Y(_23__1_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_23__3_), .Y(_273_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_274_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_275_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_275_), .C(_274_), .Y(_276_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_270_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_271_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_271_), .C(_23__3_), .Y(_272_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_276_), .Y(_21__3_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_270_), .C(_275_), .Y(_19_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_23__1_), .Y(_280_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_281_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_282_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_282_), .C(_281_), .Y(_283_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_277_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_278_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_278_), .C(_23__1_), .Y(_279_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_279_), .B(_283_), .Y(_21__1_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_277_), .C(_282_), .Y(_23__2_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_23__2_), .Y(_287_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_288_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_289_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_287_), .B(_289_), .C(_288_), .Y(_290_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_284_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_285_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_285_), .C(_23__2_), .Y(_286_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_290_), .Y(_21__2_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_287_), .B(_284_), .C(_289_), .Y(_23__3_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_294_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_295_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_296_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_296_), .C(_295_), .Y(_297_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_291_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_292_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_292_), .C(vdd), .Y(_293_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_297_), .Y(_22__0_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_291_), .C(_296_), .Y(_24__1_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_24__3_), .Y(_301_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_302_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_303_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_303_), .C(_302_), .Y(_304_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_298_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_299_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_299_), .C(_24__3_), .Y(_300_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_304_), .Y(_22__3_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_298_), .C(_303_), .Y(_20_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_24__1_), .Y(_308_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_309_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_310_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_310_), .C(_309_), .Y(_311_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_305_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_306_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_306_), .C(_24__1_), .Y(_307_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_311_), .Y(_22__1_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_305_), .C(_310_), .Y(_24__2_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_24__2_), .Y(_315_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_316_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_317_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_317_), .C(_316_), .Y(_318_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_312_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_313_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_313_), .C(_24__2_), .Y(_314_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_318_), .Y(_22__2_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_312_), .C(_317_), .Y(_24__3_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(_319_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(w_cout_4_), .Y(_320_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_319_), .C(_320_), .Y(w_cout_5_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_27__0_), .Y(_321_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_28__0_), .B(w_cout_4_), .Y(_322_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_321_), .C(_322_), .Y(_0__20_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_27__1_), .Y(_323_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_28__1_), .Y(_324_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_323_), .C(_324_), .Y(_0__21_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_27__2_), .Y(_325_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_28__2_), .Y(_326_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_325_), .C(_326_), .Y(_0__22_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_27__3_), .Y(_327_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_28__3_), .Y(_328_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_327_), .C(_328_), .Y(_0__23_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_332_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_333_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_334_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_334_), .C(_333_), .Y(_335_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_329_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_330_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_330_), .C(gnd), .Y(_331_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_335_), .Y(_27__0_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_329_), .C(_334_), .Y(_29__1_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_29__3_), .Y(_339_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_340_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_341_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_341_), .C(_340_), .Y(_342_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_336_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_337_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_337_), .C(_29__3_), .Y(_338_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_342_), .Y(_27__3_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_336_), .C(_341_), .Y(_25_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_29__1_), .Y(_346_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_347_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_348_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_348_), .C(_347_), .Y(_349_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_343_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_344_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_344_), .C(_29__1_), .Y(_345_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_349_), .Y(_27__1_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_343_), .C(_348_), .Y(_29__2_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_29__2_), .Y(_353_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_354_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_355_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_355_), .C(_354_), .Y(_356_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_350_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_351_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_351_), .C(_29__2_), .Y(_352_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_356_), .Y(_27__2_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_350_), .C(_355_), .Y(_29__3_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_360_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_361_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_362_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_362_), .C(_361_), .Y(_363_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_357_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_358_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_358_), .C(vdd), .Y(_359_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_363_), .Y(_28__0_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_357_), .C(_362_), .Y(_30__1_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_30__3_), .Y(_367_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_368_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_369_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_369_), .C(_368_), .Y(_370_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_364_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_365_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_365_), .C(_30__3_), .Y(_366_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_370_), .Y(_28__3_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_364_), .C(_369_), .Y(_26_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_30__1_), .Y(_374_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_375_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_376_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_376_), .C(_375_), .Y(_377_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_371_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_372_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_372_), .C(_30__1_), .Y(_373_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_373_), .B(_377_), .Y(_28__1_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_371_), .C(_376_), .Y(_30__2_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_30__2_), .Y(_381_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_382_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_383_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_383_), .C(_382_), .Y(_384_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_378_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_379_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_379_), .C(_30__2_), .Y(_380_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_384_), .Y(_28__2_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_378_), .C(_383_), .Y(_30__3_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_31_), .Y(_385_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(w_cout_5_), .Y(_386_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_385_), .C(_386_), .Y(w_cout_6_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_33__0_), .Y(_387_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_34__0_), .B(w_cout_5_), .Y(_388_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_387_), .C(_388_), .Y(_0__24_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_33__1_), .Y(_389_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_34__1_), .Y(_390_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_389_), .C(_390_), .Y(_0__25_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_33__2_), .Y(_391_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_34__2_), .Y(_392_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_391_), .C(_392_), .Y(_0__26_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_33__3_), .Y(_393_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_34__3_), .Y(_394_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_393_), .C(_394_), .Y(_0__27_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_398_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_399_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_400_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_400_), .C(_399_), .Y(_401_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_395_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_396_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_396_), .C(gnd), .Y(_397_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_401_), .Y(_33__0_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_395_), .C(_400_), .Y(_35__1_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_35__3_), .Y(_405_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_406_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_407_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_407_), .C(_406_), .Y(_408_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_402_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_403_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_403_), .C(_35__3_), .Y(_404_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_408_), .Y(_33__3_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_402_), .C(_407_), .Y(_31_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_35__1_), .Y(_412_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_413_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_414_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_414_), .C(_413_), .Y(_415_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_409_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_410_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_410_), .C(_35__1_), .Y(_411_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_415_), .Y(_33__1_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_409_), .C(_414_), .Y(_35__2_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_35__2_), .Y(_419_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_420_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_421_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_421_), .C(_420_), .Y(_422_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_416_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_417_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_417_), .C(_35__2_), .Y(_418_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_422_), .Y(_33__2_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_416_), .C(_421_), .Y(_35__3_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_426_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_427_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_428_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_428_), .C(_427_), .Y(_429_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_423_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_424_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_424_), .C(vdd), .Y(_425_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(_429_), .Y(_34__0_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_423_), .C(_428_), .Y(_36__1_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_36__3_), .Y(_433_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_434_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_435_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_435_), .C(_434_), .Y(_436_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_430_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_431_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_431_), .C(_36__3_), .Y(_432_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_432_), .B(_436_), .Y(_34__3_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_430_), .C(_435_), .Y(_32_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_36__1_), .Y(_440_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_441_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_442_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_442_), .C(_441_), .Y(_443_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_437_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_438_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_438_), .C(_36__1_), .Y(_439_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_443_), .Y(_34__1_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_437_), .C(_442_), .Y(_36__2_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_36__2_), .Y(_447_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_448_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_449_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_449_), .C(_448_), .Y(_450_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_444_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_445_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_445_), .C(_36__2_), .Y(_446_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(_450_), .Y(_34__2_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_444_), .C(_449_), .Y(_36__3_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_37_), .Y(_451_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(w_cout_6_), .Y(_452_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_451_), .C(_452_), .Y(w_cout_7_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_39__0_), .Y(_453_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_40__0_), .B(w_cout_6_), .Y(_454_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_453_), .C(_454_), .Y(_0__28_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_39__1_), .Y(_455_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_40__1_), .Y(_456_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_455_), .C(_456_), .Y(_0__29_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_39__2_), .Y(_457_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_40__2_), .Y(_458_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_457_), .C(_458_), .Y(_0__30_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_39__3_), .Y(_459_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_40__3_), .Y(_460_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_459_), .C(_460_), .Y(_0__31_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_464_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_465_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_466_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_466_), .C(_465_), .Y(_467_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_461_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_462_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_462_), .C(gnd), .Y(_463_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_467_), .Y(_39__0_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_461_), .C(_466_), .Y(_41__1_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_41__3_), .Y(_471_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_472_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_473_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_473_), .C(_472_), .Y(_474_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_468_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_469_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_468_), .B(_469_), .C(_41__3_), .Y(_470_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_470_), .B(_474_), .Y(_39__3_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_468_), .C(_473_), .Y(_37_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_41__1_), .Y(_478_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_479_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_480_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_480_), .C(_479_), .Y(_481_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_475_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_476_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_476_), .C(_41__1_), .Y(_477_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_477_), .B(_481_), .Y(_39__1_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_475_), .C(_480_), .Y(_41__2_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_41__2_), .Y(_485_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_486_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_487_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_487_), .C(_486_), .Y(_488_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_482_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_483_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_482_), .B(_483_), .C(_41__2_), .Y(_484_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_484_), .B(_488_), .Y(_39__2_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_482_), .C(_487_), .Y(_41__3_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_492_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_493_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_494_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_492_), .B(_494_), .C(_493_), .Y(_495_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_489_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_490_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_490_), .C(vdd), .Y(_491_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_495_), .Y(_40__0_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_492_), .B(_489_), .C(_494_), .Y(_42__1_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_42__3_), .Y(_499_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_500_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_501_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_501_), .C(_500_), .Y(_502_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_496_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_497_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_497_), .C(_42__3_), .Y(_498_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_502_), .Y(_40__3_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_496_), .C(_501_), .Y(_38_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_42__1_), .Y(_506_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_507_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_508_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_508_), .C(_507_), .Y(_509_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_503_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_504_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_504_), .C(_42__1_), .Y(_505_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(_509_), .Y(_40__1_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_503_), .C(_508_), .Y(_42__2_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_42__2_), .Y(_513_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_514_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_515_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_515_), .C(_514_), .Y(_516_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_510_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_511_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_511_), .C(_42__2_), .Y(_512_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_516_), .Y(_40__2_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_510_), .C(_515_), .Y(_42__3_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(_517_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(w_cout_7_), .Y(_518_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_517_), .C(_518_), .Y(w_cout_8_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_45__0_), .Y(_519_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_46__0_), .B(w_cout_7_), .Y(_520_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_519_), .C(_520_), .Y(_0__32_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_45__1_), .Y(_521_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_46__1_), .Y(_522_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_521_), .C(_522_), .Y(_0__33_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_45__2_), .Y(_523_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_46__2_), .Y(_524_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_523_), .C(_524_), .Y(_0__34_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_45__3_), .Y(_525_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_46__3_), .Y(_526_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_525_), .C(_526_), .Y(_0__35_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_530_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_531_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_532_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_532_), .C(_531_), .Y(_533_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_527_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_528_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_528_), .C(gnd), .Y(_529_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_533_), .Y(_45__0_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_527_), .C(_532_), .Y(_47__1_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_47__3_), .Y(_537_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_538_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_539_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_539_), .C(_538_), .Y(_540_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_534_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_535_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_535_), .C(_47__3_), .Y(_536_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_536_), .B(_540_), .Y(_45__3_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_534_), .C(_539_), .Y(_43_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_47__1_), .Y(_544_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_545_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_546_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_546_), .C(_545_), .Y(_547_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_541_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_542_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_541_), .B(_542_), .C(_47__1_), .Y(_543_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_547_), .Y(_45__1_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_541_), .C(_546_), .Y(_47__2_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_47__2_), .Y(_551_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_552_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_553_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_551_), .B(_553_), .C(_552_), .Y(_554_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_548_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_549_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_549_), .C(_47__2_), .Y(_550_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_550_), .B(_554_), .Y(_45__2_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_551_), .B(_548_), .C(_553_), .Y(_47__3_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_558_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_559_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_560_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_560_), .C(_559_), .Y(_561_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_555_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_556_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_555_), .B(_556_), .C(vdd), .Y(_557_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_557_), .B(_561_), .Y(_46__0_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_555_), .C(_560_), .Y(_48__1_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_48__3_), .Y(_565_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_566_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_567_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_567_), .C(_566_), .Y(_568_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_562_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_563_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_562_), .B(_563_), .C(_48__3_), .Y(_564_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_564_), .B(_568_), .Y(_46__3_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_562_), .C(_567_), .Y(_44_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_48__1_), .Y(_572_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_573_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_574_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_574_), .C(_573_), .Y(_575_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_569_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_570_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_569_), .B(_570_), .C(_48__1_), .Y(_571_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_575_), .Y(_46__1_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_569_), .C(_574_), .Y(_48__2_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_48__2_), .Y(_579_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_580_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_581_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_581_), .C(_580_), .Y(_582_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_576_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_577_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_576_), .B(_577_), .C(_48__2_), .Y(_578_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_578_), .B(_582_), .Y(_46__2_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_576_), .C(_581_), .Y(_48__3_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_49_), .Y(_583_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(w_cout_8_), .Y(_584_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_583_), .C(_584_), .Y(w_cout_9_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_51__0_), .Y(_585_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_52__0_), .B(w_cout_8_), .Y(_586_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_585_), .C(_586_), .Y(_0__36_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_51__1_), .Y(_587_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_52__1_), .Y(_588_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_587_), .C(_588_), .Y(_0__37_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_51__2_), .Y(_589_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_52__2_), .Y(_590_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_589_), .C(_590_), .Y(_0__38_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_51__3_), .Y(_591_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_52__3_), .Y(_592_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_591_), .C(_592_), .Y(_0__39_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_596_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_597_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_598_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_598_), .C(_597_), .Y(_599_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_593_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_594_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_594_), .C(gnd), .Y(_595_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_595_), .B(_599_), .Y(_51__0_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_593_), .C(_598_), .Y(_53__1_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_53__3_), .Y(_603_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_604_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_605_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_603_), .B(_605_), .C(_604_), .Y(_606_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_600_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_601_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_601_), .C(_53__3_), .Y(_602_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_602_), .B(_606_), .Y(_51__3_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_603_), .B(_600_), .C(_605_), .Y(_49_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_53__1_), .Y(_610_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_611_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_612_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_612_), .C(_611_), .Y(_613_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_607_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_608_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_608_), .C(_53__1_), .Y(_609_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_609_), .B(_613_), .Y(_51__1_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_607_), .C(_612_), .Y(_53__2_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_53__2_), .Y(_617_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_618_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_619_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_617_), .B(_619_), .C(_618_), .Y(_620_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_614_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_615_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_615_), .C(_53__2_), .Y(_616_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_616_), .B(_620_), .Y(_51__2_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_617_), .B(_614_), .C(_619_), .Y(_53__3_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_624_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_625_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_626_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_624_), .B(_626_), .C(_625_), .Y(_627_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_621_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_622_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_622_), .C(vdd), .Y(_623_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_623_), .B(_627_), .Y(_52__0_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_624_), .B(_621_), .C(_626_), .Y(_54__1_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_54__3_), .Y(_631_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_632_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_633_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_631_), .B(_633_), .C(_632_), .Y(_634_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_628_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_629_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_629_), .C(_54__3_), .Y(_630_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_630_), .B(_634_), .Y(_52__3_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_631_), .B(_628_), .C(_633_), .Y(_50_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(_54__1_), .Y(_638_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_639_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_640_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_640_), .C(_639_), .Y(_641_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_635_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_636_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_636_), .C(_54__1_), .Y(_637_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_637_), .B(_641_), .Y(_52__1_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_635_), .C(_640_), .Y(_54__2_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_54__2_), .Y(_645_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_646_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_647_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_645_), .B(_647_), .C(_646_), .Y(_648_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_642_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_643_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_642_), .B(_643_), .C(_54__2_), .Y(_644_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_644_), .B(_648_), .Y(_52__2_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_645_), .B(_642_), .C(_647_), .Y(_54__3_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_652_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_653_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_654_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_654_), .C(_653_), .Y(_655_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_649_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_650_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_650_), .C(gnd), .Y(_651_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_651_), .B(_655_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_649_), .C(_654_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_i_carry), .Y(_659_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_660_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_661_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(_661_), .C(_660_), .Y(_662_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_656_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_657_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_656_), .B(_657_), .C(rca_inst_fa3_i_carry), .Y(_658_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_658_), .B(_662_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(_656_), .C(_661_), .Y(rca_inst_cout) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_carry), .Y(_666_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_667_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_668_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_666_), .B(_668_), .C(_667_), .Y(_669_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_663_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_664_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(_664_), .C(rca_inst_fa0_o_carry), .Y(_665_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_665_), .B(_669_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_666_), .B(_663_), .C(_668_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_carry), .Y(_673_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_674_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_675_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(_675_), .C(_674_), .Y(_676_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_670_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_671_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(_671_), .C(rca_inst_fa_1__o_carry), .Y(_672_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_672_), .B(_676_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(_670_), .C(_675_), .Y(rca_inst_fa3_i_carry) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .Y(cout) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_0__39_), .Y(sum[39]) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_55_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(rca_inst_cout), .Y(_56_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_55_), .C(_56_), .Y(w_cout_1_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_3__0_), .Y(_57_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_4__0_), .B(rca_inst_cout), .Y(_58_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_57_), .C(_58_), .Y(_0__4_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(_3__1_), .Y(_59_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_4__1_), .Y(_60_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_59_), .C(_60_), .Y(_0__5_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_3__2_), .Y(_61_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_4__2_), .Y(_62_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_61_), .C(_62_), .Y(_0__6_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_3__3_), .Y(_63_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_4__3_), .Y(_64_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_63_), .C(_64_), .Y(_0__7_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_68_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_69_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_70_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_70_), .C(_69_), .Y(_71_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_65_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_66_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_66_), .C(gnd), .Y(_67_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_71_), .Y(_3__0_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_65_), .C(_70_), .Y(_5__1_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_5__3_), .Y(_75_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_76_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_77_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_77_), .C(_76_), .Y(_78_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_72_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_73_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_73_), .C(_5__3_), .Y(_74_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_78_), .Y(_3__3_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_72_), .C(_77_), .Y(_1_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(_5__1_), .Y(_82_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_83_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_84_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_84_), .C(_83_), .Y(_85_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_79_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_80_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_80_), .C(_5__1_), .Y(_81_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_85_), .Y(_3__1_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_79_), .C(_84_), .Y(_5__2_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_5__2_), .Y(_89_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_90_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_91_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_91_), .C(_90_), .Y(_92_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_86_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_87_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_87_), .C(_5__2_), .Y(_88_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_92_), .Y(_3__2_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_86_), .C(_91_), .Y(_5__3_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_96_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_97_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_98_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_98_), .C(_97_), .Y(_99_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_93_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_94_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_94_), .C(vdd), .Y(_95_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_99_), .Y(_4__0_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_93_), .C(_98_), .Y(_6__1_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(_6__3_), .Y(_103_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_104_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_105_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_105_), .C(_104_), .Y(_106_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_100_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_101_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_101_), .C(_6__3_), .Y(_102_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_106_), .Y(_4__3_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_100_), .C(_105_), .Y(_2_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(_6__1_), .Y(_110_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_111_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_112_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_112_), .C(_111_), .Y(_113_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_107_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_108_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_108_), .C(_6__1_), .Y(_109_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_113_), .Y(_4__1_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_107_), .C(_112_), .Y(_6__2_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(_6__2_), .Y(_117_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_118_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_119_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_119_), .C(_118_), .Y(_120_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_114_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_115_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_115_), .C(_6__2_), .Y(_116_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_120_), .Y(_4__2_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_114_), .C(_119_), .Y(_6__3_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_121_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(w_cout_1_), .Y(_122_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_121_), .C(_122_), .Y(w_cout_2_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(_9__0_), .Y(_123_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_10__0_), .B(w_cout_1_), .Y(_124_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_123_), .C(_124_), .Y(_0__8_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(_9__1_), .Y(_125_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_10__1_), .Y(_126_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_125_), .C(_126_), .Y(_0__9_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(_9__2_), .Y(_127_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_10__2_), .Y(_128_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_127_), .C(_128_), .Y(_0__10_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_9__3_), .Y(_129_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_10__3_), .Y(_130_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_129_), .C(_130_), .Y(_0__11_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_134_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_135_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_136_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_136_), .C(_135_), .Y(_137_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_131_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_132_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_132_), .C(gnd), .Y(_133_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_137_), .Y(_9__0_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_131_), .C(_136_), .Y(_11__1_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(_11__3_), .Y(_141_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_142_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_143_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_143_), .C(_142_), .Y(_144_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_138_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_139_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_139_), .C(_11__3_), .Y(_140_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_144_), .Y(_9__3_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_138_), .C(_143_), .Y(_7_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(_11__1_), .Y(_148_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_149_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_150_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_150_), .C(_149_), .Y(_151_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_145_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_146_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_146_), .C(_11__1_), .Y(_147_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_151_), .Y(_9__1_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_145_), .C(_150_), .Y(_11__2_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(_11__2_), .Y(_155_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_156_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_157_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_157_), .C(_156_), .Y(_158_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_152_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_153_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_153_), .C(_11__2_), .Y(_154_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_158_), .Y(_9__2_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_152_), .C(_157_), .Y(_11__3_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_162_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_163_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_164_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_164_), .C(_163_), .Y(_165_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_159_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_160_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_159_), .B(_160_), .C(vdd), .Y(_161_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_165_), .Y(_10__0_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_159_), .C(_164_), .Y(_12__1_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(_12__3_), .Y(_169_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_170_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_171_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_171_), .C(_170_), .Y(_172_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_166_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_167_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_167_), .C(_12__3_), .Y(_168_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_172_), .Y(_10__3_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_166_), .C(_171_), .Y(_8_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(_12__1_), .Y(_176_) );
OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_177_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_178_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_178_), .C(_177_), .Y(_179_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_173_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_174_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(_174_), .C(_12__1_), .Y(_175_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_175_), .B(_179_), .Y(_10__1_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_173_), .C(_178_), .Y(_12__2_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(_12__2_), .Y(_183_) );
OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_184_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_185_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_185_), .C(_184_), .Y(_186_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_180_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_181_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_181_), .C(_12__2_), .Y(_182_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_186_), .Y(_10__2_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_180_), .C(_185_), .Y(_12__3_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_187_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(w_cout_2_), .Y(_188_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_187_), .C(_188_), .Y(w_cout_3_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(_15__0_), .Y(_189_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_16__0_), .B(w_cout_2_), .Y(_190_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_189_), .C(_190_), .Y(_0__12_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_15__1_), .Y(_191_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_16__1_), .Y(_192_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_191_), .C(_192_), .Y(_0__13_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_15__2_), .Y(_193_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_16__2_), .Y(_194_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_193_), .C(_194_), .Y(_0__14_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_15__3_), .Y(_195_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_16__3_), .Y(_196_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_195_), .C(_196_), .Y(_0__15_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_200_) );
OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_201_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_202_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_202_), .C(_201_), .Y(_203_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_197_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_198_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_198_), .C(gnd), .Y(_199_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_203_), .Y(_15__0_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_197_), .C(_202_), .Y(_17__1_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_17__3_), .Y(_207_) );
OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_208_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_209_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_209_), .C(_208_), .Y(_210_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_204_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_205_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_205_), .C(_17__3_), .Y(_206_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_210_), .Y(_15__3_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_204_), .C(_209_), .Y(_13_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(_17__1_), .Y(_214_) );
OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_215_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_216_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_216_), .C(_215_), .Y(_217_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_211_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_212_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_212_), .C(_17__1_), .Y(_213_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_217_), .Y(_15__1_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_211_), .C(_216_), .Y(_17__2_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_17__2_), .Y(_221_) );
OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_222_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_223_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_223_), .C(_222_), .Y(_224_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_218_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_219_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(_219_), .C(_17__2_), .Y(_220_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_224_), .Y(_15__2_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_218_), .C(_223_), .Y(_17__3_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_228_) );
OR2X2 OR2X2_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_229_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_230_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_230_), .C(_229_), .Y(_231_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_225_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_226_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_226_), .C(vdd), .Y(_227_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_231_), .Y(_16__0_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_225_), .C(_230_), .Y(_18__1_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(_18__3_), .Y(_235_) );
OR2X2 OR2X2_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_236_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_237_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_237_), .C(_236_), .Y(_238_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_232_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_233_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_233_), .C(_18__3_), .Y(_234_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_238_), .Y(_16__3_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_232_), .C(_237_), .Y(_14_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(_18__1_), .Y(_242_) );
OR2X2 OR2X2_74 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_243_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_244_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_244_), .C(_243_), .Y(_245_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_239_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_240_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_240_), .C(_18__1_), .Y(_241_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_245_), .Y(_16__1_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_239_), .C(_244_), .Y(_18__2_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(_18__2_), .Y(_249_) );
OR2X2 OR2X2_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_250_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_251_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_251_), .C(_250_), .Y(_252_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_246_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_247_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_247_), .C(_18__2_), .Y(_248_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_252_), .Y(_16__2_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_246_), .C(_251_), .Y(_18__3_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_253_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(w_cout_3_), .Y(_254_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_253_), .C(_254_), .Y(w_cout_4_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(_21__0_), .Y(_255_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_22__0_), .B(w_cout_3_), .Y(_256_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_255_), .C(_256_), .Y(_0__16_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(_21__1_), .Y(_257_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_22__1_), .Y(_258_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_257_), .C(_258_), .Y(_0__17_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(_21__2_), .Y(_259_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_22__2_), .Y(_260_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_259_), .C(_260_), .Y(_0__18_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(_21__3_), .Y(_261_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_22__3_), .Y(_262_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_261_), .C(_262_), .Y(_0__19_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_266_) );
OR2X2 OR2X2_76 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_267_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_268_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_268_), .C(_267_), .Y(_269_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_263_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_264_) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .Y(w_cout_0_) );
endmodule
