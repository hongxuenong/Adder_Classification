module cla_25bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add1[19], i_add1[20], i_add1[21], i_add1[22], i_add1[23], i_add1[24], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], i_add2[19], i_add2[20], i_add2[21], i_add2[22], i_add2[23], i_add2[24], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21], o_result[22], o_result[23], o_result[24], o_result[25]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add1[19];
input i_add1[20];
input i_add1[21];
input i_add1[22];
input i_add1[23];
input i_add1[24];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
input i_add2[19];
input i_add2[20];
input i_add2[21];
input i_add2[22];
input i_add2[23];
input i_add2[24];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];
output o_result[22];
output o_result[23];
output o_result[24];
output o_result[25];

NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_106_) );
INVX1 INVX1_1 ( .A(_106_), .Y(w_C_1_) );
NAND2X1 NAND2X1_2 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_107_) );
NAND2X1 NAND2X1_3 ( .A(_106_), .B(_107_), .Y(_108_) );
OAI21X1 OAI21X1_1 ( .A(i_add2[1]), .B(i_add1[1]), .C(_108_), .Y(_109_) );
INVX1 INVX1_2 ( .A(_109_), .Y(w_C_2_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_110_) );
OR2X2 OR2X2_1 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_111_) );
OR2X2 OR2X2_2 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_112_) );
NAND3X1 NAND3X1_1 ( .A(_111_), .B(_112_), .C(_108_), .Y(_113_) );
NAND2X1 NAND2X1_5 ( .A(_110_), .B(_113_), .Y(w_C_3_) );
OR2X2 OR2X2_3 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_114_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_115_) );
NAND3X1 NAND3X1_2 ( .A(_110_), .B(_115_), .C(_113_), .Y(_116_) );
AND2X2 AND2X2_1 ( .A(_116_), .B(_114_), .Y(w_C_4_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_117_) );
OR2X2 OR2X2_4 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_118_) );
NAND3X1 NAND3X1_3 ( .A(_114_), .B(_118_), .C(_116_), .Y(_119_) );
NAND2X1 NAND2X1_8 ( .A(_117_), .B(_119_), .Y(w_C_5_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_120_) );
INVX1 INVX1_3 ( .A(_120_), .Y(_121_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_122_) );
NAND3X1 NAND3X1_4 ( .A(_117_), .B(_122_), .C(_119_), .Y(_123_) );
AND2X2 AND2X2_2 ( .A(_123_), .B(_121_), .Y(w_C_6_) );
AND2X2 AND2X2_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_0_) );
INVX1 INVX1_4 ( .A(_0_), .Y(_1_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_2_) );
INVX1 INVX1_5 ( .A(_2_), .Y(_3_) );
NAND3X1 NAND3X1_5 ( .A(_121_), .B(_3_), .C(_123_), .Y(_4_) );
AND2X2 AND2X2_4 ( .A(_4_), .B(_1_), .Y(_5_) );
INVX1 INVX1_6 ( .A(_5_), .Y(w_C_7_) );
AND2X2 AND2X2_5 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_6_) );
INVX1 INVX1_7 ( .A(_6_), .Y(_7_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_8_) );
OAI21X1 OAI21X1_2 ( .A(_8_), .B(_5_), .C(_7_), .Y(w_C_8_) );
AND2X2 AND2X2_6 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_9_) );
INVX1 INVX1_8 ( .A(_9_), .Y(_10_) );
INVX1 INVX1_9 ( .A(_8_), .Y(_11_) );
NAND3X1 NAND3X1_6 ( .A(_1_), .B(_7_), .C(_4_), .Y(_12_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_13_) );
INVX1 INVX1_10 ( .A(_13_), .Y(_14_) );
NAND3X1 NAND3X1_7 ( .A(_11_), .B(_14_), .C(_12_), .Y(_15_) );
AND2X2 AND2X2_7 ( .A(_15_), .B(_10_), .Y(_16_) );
INVX1 INVX1_11 ( .A(_16_), .Y(w_C_9_) );
AND2X2 AND2X2_8 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_17_) );
INVX1 INVX1_12 ( .A(_17_), .Y(_18_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_19_) );
OAI21X1 OAI21X1_3 ( .A(_19_), .B(_16_), .C(_18_), .Y(w_C_10_) );
INVX1 INVX1_13 ( .A(i_add2[10]), .Y(_20_) );
INVX1 INVX1_14 ( .A(i_add1[10]), .Y(_21_) );
INVX1 INVX1_15 ( .A(_19_), .Y(_22_) );
NAND3X1 NAND3X1_8 ( .A(_10_), .B(_18_), .C(_15_), .Y(_23_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_24_) );
INVX1 INVX1_16 ( .A(_24_), .Y(_25_) );
NAND3X1 NAND3X1_9 ( .A(_22_), .B(_25_), .C(_23_), .Y(_26_) );
OAI21X1 OAI21X1_4 ( .A(_20_), .B(_21_), .C(_26_), .Y(w_C_11_) );
NOR2X1 NOR2X1_7 ( .A(_20_), .B(_21_), .Y(_27_) );
INVX1 INVX1_17 ( .A(_27_), .Y(_28_) );
AND2X2 AND2X2_9 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_29_) );
INVX1 INVX1_18 ( .A(_29_), .Y(_30_) );
NAND3X1 NAND3X1_10 ( .A(_28_), .B(_30_), .C(_26_), .Y(_31_) );
OAI21X1 OAI21X1_5 ( .A(i_add2[11]), .B(i_add1[11]), .C(_31_), .Y(_32_) );
INVX1 INVX1_19 ( .A(_32_), .Y(w_C_12_) );
INVX1 INVX1_20 ( .A(i_add2[12]), .Y(_33_) );
INVX1 INVX1_21 ( .A(i_add1[12]), .Y(_34_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_35_) );
INVX1 INVX1_22 ( .A(_35_), .Y(_36_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_37_) );
INVX1 INVX1_23 ( .A(_37_), .Y(_38_) );
NAND3X1 NAND3X1_11 ( .A(_36_), .B(_38_), .C(_31_), .Y(_39_) );
OAI21X1 OAI21X1_6 ( .A(_33_), .B(_34_), .C(_39_), .Y(w_C_13_) );
NOR2X1 NOR2X1_10 ( .A(_33_), .B(_34_), .Y(_40_) );
INVX1 INVX1_24 ( .A(_40_), .Y(_41_) );
AND2X2 AND2X2_10 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_42_) );
INVX1 INVX1_25 ( .A(_42_), .Y(_43_) );
NAND3X1 NAND3X1_12 ( .A(_41_), .B(_43_), .C(_39_), .Y(_44_) );
OAI21X1 OAI21X1_7 ( .A(i_add2[13]), .B(i_add1[13]), .C(_44_), .Y(_45_) );
INVX1 INVX1_26 ( .A(_45_), .Y(w_C_14_) );
INVX1 INVX1_27 ( .A(i_add2[14]), .Y(_46_) );
INVX1 INVX1_28 ( .A(i_add1[14]), .Y(_47_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_48_) );
INVX1 INVX1_29 ( .A(_48_), .Y(_49_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_50_) );
INVX1 INVX1_30 ( .A(_50_), .Y(_51_) );
NAND3X1 NAND3X1_13 ( .A(_49_), .B(_51_), .C(_44_), .Y(_52_) );
OAI21X1 OAI21X1_8 ( .A(_46_), .B(_47_), .C(_52_), .Y(w_C_15_) );
NOR2X1 NOR2X1_13 ( .A(_46_), .B(_47_), .Y(_53_) );
INVX1 INVX1_31 ( .A(_53_), .Y(_54_) );
AND2X2 AND2X2_11 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_55_) );
INVX1 INVX1_32 ( .A(_55_), .Y(_56_) );
NAND3X1 NAND3X1_14 ( .A(_54_), .B(_56_), .C(_52_), .Y(_57_) );
OAI21X1 OAI21X1_9 ( .A(i_add2[15]), .B(i_add1[15]), .C(_57_), .Y(_58_) );
INVX1 INVX1_33 ( .A(_58_), .Y(w_C_16_) );
INVX1 INVX1_34 ( .A(i_add2[16]), .Y(_59_) );
INVX1 INVX1_35 ( .A(i_add1[16]), .Y(_60_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_61_) );
INVX1 INVX1_36 ( .A(_61_), .Y(_62_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_63_) );
INVX1 INVX1_37 ( .A(_63_), .Y(_64_) );
NAND3X1 NAND3X1_15 ( .A(_62_), .B(_64_), .C(_57_), .Y(_65_) );
OAI21X1 OAI21X1_10 ( .A(_59_), .B(_60_), .C(_65_), .Y(w_C_17_) );
NOR2X1 NOR2X1_16 ( .A(_59_), .B(_60_), .Y(_66_) );
INVX1 INVX1_38 ( .A(_66_), .Y(_67_) );
AND2X2 AND2X2_12 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_68_) );
INVX1 INVX1_39 ( .A(_68_), .Y(_69_) );
NAND3X1 NAND3X1_16 ( .A(_67_), .B(_69_), .C(_65_), .Y(_70_) );
OAI21X1 OAI21X1_11 ( .A(i_add2[17]), .B(i_add1[17]), .C(_70_), .Y(_71_) );
INVX1 INVX1_40 ( .A(_71_), .Y(w_C_18_) );
INVX1 INVX1_41 ( .A(i_add2[18]), .Y(_72_) );
INVX1 INVX1_42 ( .A(i_add1[18]), .Y(_73_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_74_) );
INVX1 INVX1_43 ( .A(_74_), .Y(_75_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_76_) );
INVX1 INVX1_44 ( .A(_76_), .Y(_77_) );
NAND3X1 NAND3X1_17 ( .A(_75_), .B(_77_), .C(_70_), .Y(_78_) );
OAI21X1 OAI21X1_12 ( .A(_72_), .B(_73_), .C(_78_), .Y(w_C_19_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_79_) );
INVX1 INVX1_45 ( .A(_79_), .Y(_80_) );
NOR2X1 NOR2X1_20 ( .A(_72_), .B(_73_), .Y(_81_) );
INVX1 INVX1_46 ( .A(_81_), .Y(_82_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_83_) );
NAND3X1 NAND3X1_18 ( .A(_82_), .B(_83_), .C(_78_), .Y(_84_) );
AND2X2 AND2X2_13 ( .A(_84_), .B(_80_), .Y(w_C_20_) );
INVX1 INVX1_47 ( .A(i_add2[20]), .Y(_85_) );
INVX1 INVX1_48 ( .A(i_add1[20]), .Y(_86_) );
NAND2X1 NAND2X1_11 ( .A(_85_), .B(_86_), .Y(_87_) );
NAND3X1 NAND3X1_19 ( .A(_80_), .B(_87_), .C(_84_), .Y(_88_) );
OAI21X1 OAI21X1_13 ( .A(_85_), .B(_86_), .C(_88_), .Y(w_C_21_) );
INVX1 INVX1_49 ( .A(i_add2[21]), .Y(_89_) );
INVX1 INVX1_50 ( .A(i_add1[21]), .Y(_90_) );
NAND2X1 NAND2X1_12 ( .A(_89_), .B(_90_), .Y(_91_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_92_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_93_) );
NAND3X1 NAND3X1_20 ( .A(_92_), .B(_93_), .C(_88_), .Y(_94_) );
AND2X2 AND2X2_14 ( .A(_94_), .B(_91_), .Y(w_C_22_) );
INVX1 INVX1_51 ( .A(i_add2[22]), .Y(_95_) );
INVX1 INVX1_52 ( .A(i_add1[22]), .Y(_96_) );
NAND2X1 NAND2X1_15 ( .A(_95_), .B(_96_), .Y(_97_) );
NAND3X1 NAND3X1_21 ( .A(_91_), .B(_97_), .C(_94_), .Y(_98_) );
OAI21X1 OAI21X1_14 ( .A(_95_), .B(_96_), .C(_98_), .Y(w_C_23_) );
OR2X2 OR2X2_5 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_99_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_100_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_101_) );
NAND3X1 NAND3X1_22 ( .A(_100_), .B(_101_), .C(_98_), .Y(_102_) );
AND2X2 AND2X2_15 ( .A(_102_), .B(_99_), .Y(w_C_24_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_103_) );
OR2X2 OR2X2_6 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_104_) );
NAND3X1 NAND3X1_23 ( .A(_99_), .B(_104_), .C(_102_), .Y(_105_) );
NAND2X1 NAND2X1_19 ( .A(_103_), .B(_105_), .Y(w_C_25_) );
BUFX2 BUFX2_1 ( .A(_124__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_124__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_124__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_124__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_124__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_124__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_124__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_124__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_124__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_124__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_124__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_124__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_124__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_124__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_124__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_124__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_124__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_124__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_124__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_124__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_124__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_124__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_124__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_124__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_124__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(w_C_25_), .Y(o_result[25]) );
INVX1 INVX1_53 ( .A(w_C_4_), .Y(_128_) );
OR2X2 OR2X2_7 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_129_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_130_) );
NAND3X1 NAND3X1_24 ( .A(_128_), .B(_130_), .C(_129_), .Y(_131_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_125_) );
AND2X2 AND2X2_16 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_126_) );
OAI21X1 OAI21X1_15 ( .A(_125_), .B(_126_), .C(w_C_4_), .Y(_127_) );
NAND2X1 NAND2X1_21 ( .A(_127_), .B(_131_), .Y(_124__4_) );
INVX1 INVX1_54 ( .A(w_C_5_), .Y(_135_) );
OR2X2 OR2X2_8 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_136_) );
NAND2X1 NAND2X1_22 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_137_) );
NAND3X1 NAND3X1_25 ( .A(_135_), .B(_137_), .C(_136_), .Y(_138_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_132_) );
AND2X2 AND2X2_17 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_133_) );
OAI21X1 OAI21X1_16 ( .A(_132_), .B(_133_), .C(w_C_5_), .Y(_134_) );
NAND2X1 NAND2X1_23 ( .A(_134_), .B(_138_), .Y(_124__5_) );
INVX1 INVX1_55 ( .A(w_C_6_), .Y(_142_) );
OR2X2 OR2X2_9 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_143_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_144_) );
NAND3X1 NAND3X1_26 ( .A(_142_), .B(_144_), .C(_143_), .Y(_145_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_139_) );
AND2X2 AND2X2_18 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_140_) );
OAI21X1 OAI21X1_17 ( .A(_139_), .B(_140_), .C(w_C_6_), .Y(_141_) );
NAND2X1 NAND2X1_25 ( .A(_141_), .B(_145_), .Y(_124__6_) );
INVX1 INVX1_56 ( .A(w_C_7_), .Y(_149_) );
OR2X2 OR2X2_10 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_150_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_151_) );
NAND3X1 NAND3X1_27 ( .A(_149_), .B(_151_), .C(_150_), .Y(_152_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_146_) );
AND2X2 AND2X2_19 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_147_) );
OAI21X1 OAI21X1_18 ( .A(_146_), .B(_147_), .C(w_C_7_), .Y(_148_) );
NAND2X1 NAND2X1_27 ( .A(_148_), .B(_152_), .Y(_124__7_) );
INVX1 INVX1_57 ( .A(w_C_8_), .Y(_156_) );
OR2X2 OR2X2_11 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_157_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_158_) );
NAND3X1 NAND3X1_28 ( .A(_156_), .B(_158_), .C(_157_), .Y(_159_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_153_) );
AND2X2 AND2X2_20 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_154_) );
OAI21X1 OAI21X1_19 ( .A(_153_), .B(_154_), .C(w_C_8_), .Y(_155_) );
NAND2X1 NAND2X1_29 ( .A(_155_), .B(_159_), .Y(_124__8_) );
INVX1 INVX1_58 ( .A(w_C_9_), .Y(_163_) );
OR2X2 OR2X2_12 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_164_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_165_) );
NAND3X1 NAND3X1_29 ( .A(_163_), .B(_165_), .C(_164_), .Y(_166_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_160_) );
AND2X2 AND2X2_21 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_161_) );
OAI21X1 OAI21X1_20 ( .A(_160_), .B(_161_), .C(w_C_9_), .Y(_162_) );
NAND2X1 NAND2X1_31 ( .A(_162_), .B(_166_), .Y(_124__9_) );
INVX1 INVX1_59 ( .A(w_C_10_), .Y(_170_) );
OR2X2 OR2X2_13 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_171_) );
NAND2X1 NAND2X1_32 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_172_) );
NAND3X1 NAND3X1_30 ( .A(_170_), .B(_172_), .C(_171_), .Y(_173_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_167_) );
AND2X2 AND2X2_22 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_168_) );
OAI21X1 OAI21X1_21 ( .A(_167_), .B(_168_), .C(w_C_10_), .Y(_169_) );
NAND2X1 NAND2X1_33 ( .A(_169_), .B(_173_), .Y(_124__10_) );
INVX1 INVX1_60 ( .A(w_C_11_), .Y(_177_) );
OR2X2 OR2X2_14 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_178_) );
NAND2X1 NAND2X1_34 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_179_) );
NAND3X1 NAND3X1_31 ( .A(_177_), .B(_179_), .C(_178_), .Y(_180_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_174_) );
AND2X2 AND2X2_23 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_175_) );
OAI21X1 OAI21X1_22 ( .A(_174_), .B(_175_), .C(w_C_11_), .Y(_176_) );
NAND2X1 NAND2X1_35 ( .A(_176_), .B(_180_), .Y(_124__11_) );
INVX1 INVX1_61 ( .A(w_C_12_), .Y(_184_) );
OR2X2 OR2X2_15 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_185_) );
NAND2X1 NAND2X1_36 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_186_) );
NAND3X1 NAND3X1_32 ( .A(_184_), .B(_186_), .C(_185_), .Y(_187_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_181_) );
AND2X2 AND2X2_24 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_182_) );
OAI21X1 OAI21X1_23 ( .A(_181_), .B(_182_), .C(w_C_12_), .Y(_183_) );
NAND2X1 NAND2X1_37 ( .A(_183_), .B(_187_), .Y(_124__12_) );
INVX1 INVX1_62 ( .A(w_C_13_), .Y(_191_) );
OR2X2 OR2X2_16 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_192_) );
NAND2X1 NAND2X1_38 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_193_) );
NAND3X1 NAND3X1_33 ( .A(_191_), .B(_193_), .C(_192_), .Y(_194_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_188_) );
AND2X2 AND2X2_25 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_189_) );
OAI21X1 OAI21X1_24 ( .A(_188_), .B(_189_), .C(w_C_13_), .Y(_190_) );
NAND2X1 NAND2X1_39 ( .A(_190_), .B(_194_), .Y(_124__13_) );
INVX1 INVX1_63 ( .A(w_C_14_), .Y(_198_) );
OR2X2 OR2X2_17 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_199_) );
NAND2X1 NAND2X1_40 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_200_) );
NAND3X1 NAND3X1_34 ( .A(_198_), .B(_200_), .C(_199_), .Y(_201_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_195_) );
AND2X2 AND2X2_26 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_196_) );
OAI21X1 OAI21X1_25 ( .A(_195_), .B(_196_), .C(w_C_14_), .Y(_197_) );
NAND2X1 NAND2X1_41 ( .A(_197_), .B(_201_), .Y(_124__14_) );
INVX1 INVX1_64 ( .A(w_C_15_), .Y(_205_) );
OR2X2 OR2X2_18 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_206_) );
NAND2X1 NAND2X1_42 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_207_) );
NAND3X1 NAND3X1_35 ( .A(_205_), .B(_207_), .C(_206_), .Y(_208_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_202_) );
AND2X2 AND2X2_27 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_203_) );
OAI21X1 OAI21X1_26 ( .A(_202_), .B(_203_), .C(w_C_15_), .Y(_204_) );
NAND2X1 NAND2X1_43 ( .A(_204_), .B(_208_), .Y(_124__15_) );
INVX1 INVX1_65 ( .A(w_C_16_), .Y(_212_) );
OR2X2 OR2X2_19 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_213_) );
NAND2X1 NAND2X1_44 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_214_) );
NAND3X1 NAND3X1_36 ( .A(_212_), .B(_214_), .C(_213_), .Y(_215_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_209_) );
AND2X2 AND2X2_28 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_210_) );
OAI21X1 OAI21X1_27 ( .A(_209_), .B(_210_), .C(w_C_16_), .Y(_211_) );
NAND2X1 NAND2X1_45 ( .A(_211_), .B(_215_), .Y(_124__16_) );
INVX1 INVX1_66 ( .A(w_C_17_), .Y(_219_) );
OR2X2 OR2X2_20 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_220_) );
NAND2X1 NAND2X1_46 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_221_) );
NAND3X1 NAND3X1_37 ( .A(_219_), .B(_221_), .C(_220_), .Y(_222_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_216_) );
AND2X2 AND2X2_29 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_217_) );
OAI21X1 OAI21X1_28 ( .A(_216_), .B(_217_), .C(w_C_17_), .Y(_218_) );
NAND2X1 NAND2X1_47 ( .A(_218_), .B(_222_), .Y(_124__17_) );
INVX1 INVX1_67 ( .A(w_C_18_), .Y(_226_) );
OR2X2 OR2X2_21 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_227_) );
NAND2X1 NAND2X1_48 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_228_) );
NAND3X1 NAND3X1_38 ( .A(_226_), .B(_228_), .C(_227_), .Y(_229_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_223_) );
AND2X2 AND2X2_30 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_224_) );
OAI21X1 OAI21X1_29 ( .A(_223_), .B(_224_), .C(w_C_18_), .Y(_225_) );
NAND2X1 NAND2X1_49 ( .A(_225_), .B(_229_), .Y(_124__18_) );
INVX1 INVX1_68 ( .A(w_C_19_), .Y(_233_) );
OR2X2 OR2X2_22 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_234_) );
NAND2X1 NAND2X1_50 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_235_) );
NAND3X1 NAND3X1_39 ( .A(_233_), .B(_235_), .C(_234_), .Y(_236_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_230_) );
AND2X2 AND2X2_31 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_231_) );
OAI21X1 OAI21X1_30 ( .A(_230_), .B(_231_), .C(w_C_19_), .Y(_232_) );
NAND2X1 NAND2X1_51 ( .A(_232_), .B(_236_), .Y(_124__19_) );
INVX1 INVX1_69 ( .A(w_C_20_), .Y(_240_) );
OR2X2 OR2X2_23 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_241_) );
NAND2X1 NAND2X1_52 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_242_) );
NAND3X1 NAND3X1_40 ( .A(_240_), .B(_242_), .C(_241_), .Y(_243_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_237_) );
AND2X2 AND2X2_32 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_238_) );
OAI21X1 OAI21X1_31 ( .A(_237_), .B(_238_), .C(w_C_20_), .Y(_239_) );
NAND2X1 NAND2X1_53 ( .A(_239_), .B(_243_), .Y(_124__20_) );
INVX1 INVX1_70 ( .A(w_C_21_), .Y(_247_) );
OR2X2 OR2X2_24 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_248_) );
NAND2X1 NAND2X1_54 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_249_) );
NAND3X1 NAND3X1_41 ( .A(_247_), .B(_249_), .C(_248_), .Y(_250_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_244_) );
AND2X2 AND2X2_33 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_245_) );
OAI21X1 OAI21X1_32 ( .A(_244_), .B(_245_), .C(w_C_21_), .Y(_246_) );
NAND2X1 NAND2X1_55 ( .A(_246_), .B(_250_), .Y(_124__21_) );
INVX1 INVX1_71 ( .A(w_C_22_), .Y(_254_) );
OR2X2 OR2X2_25 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_255_) );
NAND2X1 NAND2X1_56 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_256_) );
NAND3X1 NAND3X1_42 ( .A(_254_), .B(_256_), .C(_255_), .Y(_257_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_251_) );
AND2X2 AND2X2_34 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_252_) );
OAI21X1 OAI21X1_33 ( .A(_251_), .B(_252_), .C(w_C_22_), .Y(_253_) );
NAND2X1 NAND2X1_57 ( .A(_253_), .B(_257_), .Y(_124__22_) );
INVX1 INVX1_72 ( .A(w_C_23_), .Y(_261_) );
OR2X2 OR2X2_26 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_262_) );
NAND2X1 NAND2X1_58 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_263_) );
NAND3X1 NAND3X1_43 ( .A(_261_), .B(_263_), .C(_262_), .Y(_264_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_258_) );
AND2X2 AND2X2_35 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_259_) );
OAI21X1 OAI21X1_34 ( .A(_258_), .B(_259_), .C(w_C_23_), .Y(_260_) );
NAND2X1 NAND2X1_59 ( .A(_260_), .B(_264_), .Y(_124__23_) );
INVX1 INVX1_73 ( .A(w_C_24_), .Y(_268_) );
OR2X2 OR2X2_27 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_269_) );
NAND2X1 NAND2X1_60 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_270_) );
NAND3X1 NAND3X1_44 ( .A(_268_), .B(_270_), .C(_269_), .Y(_271_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_265_) );
AND2X2 AND2X2_36 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_266_) );
OAI21X1 OAI21X1_35 ( .A(_265_), .B(_266_), .C(w_C_24_), .Y(_267_) );
NAND2X1 NAND2X1_61 ( .A(_267_), .B(_271_), .Y(_124__24_) );
INVX1 INVX1_74 ( .A(1'b0), .Y(_275_) );
OR2X2 OR2X2_28 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_276_) );
NAND2X1 NAND2X1_62 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_277_) );
NAND3X1 NAND3X1_45 ( .A(_275_), .B(_277_), .C(_276_), .Y(_278_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_272_) );
AND2X2 AND2X2_37 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_273_) );
OAI21X1 OAI21X1_36 ( .A(_272_), .B(_273_), .C(1'b0), .Y(_274_) );
NAND2X1 NAND2X1_63 ( .A(_274_), .B(_278_), .Y(_124__0_) );
INVX1 INVX1_75 ( .A(w_C_1_), .Y(_282_) );
OR2X2 OR2X2_29 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_283_) );
NAND2X1 NAND2X1_64 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_284_) );
NAND3X1 NAND3X1_46 ( .A(_282_), .B(_284_), .C(_283_), .Y(_285_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_279_) );
AND2X2 AND2X2_38 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_280_) );
OAI21X1 OAI21X1_37 ( .A(_279_), .B(_280_), .C(w_C_1_), .Y(_281_) );
NAND2X1 NAND2X1_65 ( .A(_281_), .B(_285_), .Y(_124__1_) );
INVX1 INVX1_76 ( .A(w_C_2_), .Y(_289_) );
OR2X2 OR2X2_30 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_290_) );
NAND2X1 NAND2X1_66 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_291_) );
NAND3X1 NAND3X1_47 ( .A(_289_), .B(_291_), .C(_290_), .Y(_292_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_286_) );
AND2X2 AND2X2_39 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_287_) );
OAI21X1 OAI21X1_38 ( .A(_286_), .B(_287_), .C(w_C_2_), .Y(_288_) );
NAND2X1 NAND2X1_67 ( .A(_288_), .B(_292_), .Y(_124__2_) );
INVX1 INVX1_77 ( .A(w_C_3_), .Y(_296_) );
OR2X2 OR2X2_31 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_297_) );
NAND2X1 NAND2X1_68 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_298_) );
NAND3X1 NAND3X1_48 ( .A(_296_), .B(_298_), .C(_297_), .Y(_299_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_293_) );
AND2X2 AND2X2_40 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_294_) );
OAI21X1 OAI21X1_39 ( .A(_293_), .B(_294_), .C(w_C_3_), .Y(_295_) );
NAND2X1 NAND2X1_69 ( .A(_295_), .B(_299_), .Y(_124__3_) );
BUFX2 BUFX2_27 ( .A(w_C_25_), .Y(_124__25_) );
BUFX2 BUFX2_28 ( .A(1'b0), .Y(w_C_0_) );
endmodule
