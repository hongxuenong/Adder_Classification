module cla_24bit (i_add1, i_add2, o_result);

input [23:0] i_add1;
input [23:0] i_add2;
output [24:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_100_) );
INVX1 INVX1_1 ( .A(_100_), .Y(w_C_1_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_101_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_102_) );
NOR2X1 NOR2X1_2 ( .A(_101_), .B(_102_), .Y(w_C_2_) );
INVX1 INVX1_2 ( .A(i_add2[2]), .Y(_103_) );
INVX1 INVX1_3 ( .A(i_add1[2]), .Y(_104_) );
NAND2X1 NAND2X1_2 ( .A(_103_), .B(_104_), .Y(_105_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_106_) );
OAI21X1 OAI21X1_1 ( .A(_101_), .B(_102_), .C(_106_), .Y(_107_) );
AND2X2 AND2X2_1 ( .A(_107_), .B(_105_), .Y(w_C_3_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_108_) );
OR2X2 OR2X2_1 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_109_) );
NAND3X1 NAND3X1_1 ( .A(_105_), .B(_109_), .C(_107_), .Y(_110_) );
NAND2X1 NAND2X1_5 ( .A(_108_), .B(_110_), .Y(w_C_4_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_111_) );
INVX1 INVX1_4 ( .A(_111_), .Y(_112_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_113_) );
NAND3X1 NAND3X1_2 ( .A(_108_), .B(_113_), .C(_110_), .Y(_114_) );
AND2X2 AND2X2_2 ( .A(_114_), .B(_112_), .Y(w_C_5_) );
AND2X2 AND2X2_3 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_115_) );
INVX1 INVX1_5 ( .A(_115_), .Y(_116_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_117_) );
INVX1 INVX1_6 ( .A(_117_), .Y(_118_) );
NAND3X1 NAND3X1_3 ( .A(_112_), .B(_118_), .C(_114_), .Y(_119_) );
AND2X2 AND2X2_4 ( .A(_119_), .B(_116_), .Y(_120_) );
INVX1 INVX1_7 ( .A(_120_), .Y(w_C_6_) );
AND2X2 AND2X2_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_0_) );
INVX1 INVX1_8 ( .A(_0_), .Y(_1_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_2_) );
OAI21X1 OAI21X1_2 ( .A(_2_), .B(_120_), .C(_1_), .Y(w_C_7_) );
AND2X2 AND2X2_6 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_3_) );
INVX1 INVX1_9 ( .A(_3_), .Y(_4_) );
INVX1 INVX1_10 ( .A(_2_), .Y(_5_) );
NAND3X1 NAND3X1_4 ( .A(_116_), .B(_1_), .C(_119_), .Y(_6_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_7_) );
INVX1 INVX1_11 ( .A(_7_), .Y(_8_) );
NAND3X1 NAND3X1_5 ( .A(_5_), .B(_8_), .C(_6_), .Y(_9_) );
AND2X2 AND2X2_7 ( .A(_9_), .B(_4_), .Y(_10_) );
INVX1 INVX1_12 ( .A(_10_), .Y(w_C_8_) );
AND2X2 AND2X2_8 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_11_) );
INVX1 INVX1_13 ( .A(_11_), .Y(_12_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_13_) );
OAI21X1 OAI21X1_3 ( .A(_13_), .B(_10_), .C(_12_), .Y(w_C_9_) );
INVX1 INVX1_14 ( .A(i_add2[9]), .Y(_14_) );
INVX1 INVX1_15 ( .A(i_add1[9]), .Y(_15_) );
INVX1 INVX1_16 ( .A(_13_), .Y(_16_) );
NAND3X1 NAND3X1_6 ( .A(_4_), .B(_12_), .C(_9_), .Y(_17_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_18_) );
INVX1 INVX1_17 ( .A(_18_), .Y(_19_) );
NAND3X1 NAND3X1_7 ( .A(_16_), .B(_19_), .C(_17_), .Y(_20_) );
OAI21X1 OAI21X1_4 ( .A(_14_), .B(_15_), .C(_20_), .Y(w_C_10_) );
NOR2X1 NOR2X1_9 ( .A(_14_), .B(_15_), .Y(_21_) );
INVX1 INVX1_18 ( .A(_21_), .Y(_22_) );
AND2X2 AND2X2_9 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_23_) );
INVX1 INVX1_19 ( .A(_23_), .Y(_24_) );
NAND3X1 NAND3X1_8 ( .A(_22_), .B(_24_), .C(_20_), .Y(_25_) );
OAI21X1 OAI21X1_5 ( .A(i_add2[10]), .B(i_add1[10]), .C(_25_), .Y(_26_) );
INVX1 INVX1_20 ( .A(_26_), .Y(w_C_11_) );
INVX1 INVX1_21 ( .A(i_add2[11]), .Y(_27_) );
INVX1 INVX1_22 ( .A(i_add1[11]), .Y(_28_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_29_) );
INVX1 INVX1_23 ( .A(_29_), .Y(_30_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_31_) );
INVX1 INVX1_24 ( .A(_31_), .Y(_32_) );
NAND3X1 NAND3X1_9 ( .A(_30_), .B(_32_), .C(_25_), .Y(_33_) );
OAI21X1 OAI21X1_6 ( .A(_27_), .B(_28_), .C(_33_), .Y(w_C_12_) );
NOR2X1 NOR2X1_12 ( .A(_27_), .B(_28_), .Y(_34_) );
INVX1 INVX1_25 ( .A(_34_), .Y(_35_) );
AND2X2 AND2X2_10 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_36_) );
INVX1 INVX1_26 ( .A(_36_), .Y(_37_) );
NAND3X1 NAND3X1_10 ( .A(_35_), .B(_37_), .C(_33_), .Y(_38_) );
OAI21X1 OAI21X1_7 ( .A(i_add2[12]), .B(i_add1[12]), .C(_38_), .Y(_39_) );
INVX1 INVX1_27 ( .A(_39_), .Y(w_C_13_) );
INVX1 INVX1_28 ( .A(i_add2[13]), .Y(_40_) );
INVX1 INVX1_29 ( .A(i_add1[13]), .Y(_41_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_42_) );
INVX1 INVX1_30 ( .A(_42_), .Y(_43_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_44_) );
INVX1 INVX1_31 ( .A(_44_), .Y(_45_) );
NAND3X1 NAND3X1_11 ( .A(_43_), .B(_45_), .C(_38_), .Y(_46_) );
OAI21X1 OAI21X1_8 ( .A(_40_), .B(_41_), .C(_46_), .Y(w_C_14_) );
NOR2X1 NOR2X1_15 ( .A(_40_), .B(_41_), .Y(_47_) );
INVX1 INVX1_32 ( .A(_47_), .Y(_48_) );
AND2X2 AND2X2_11 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_49_) );
INVX1 INVX1_33 ( .A(_49_), .Y(_50_) );
NAND3X1 NAND3X1_12 ( .A(_48_), .B(_50_), .C(_46_), .Y(_51_) );
OAI21X1 OAI21X1_9 ( .A(i_add2[14]), .B(i_add1[14]), .C(_51_), .Y(_52_) );
INVX1 INVX1_34 ( .A(_52_), .Y(w_C_15_) );
INVX1 INVX1_35 ( .A(i_add2[15]), .Y(_53_) );
INVX1 INVX1_36 ( .A(i_add1[15]), .Y(_54_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_55_) );
INVX1 INVX1_37 ( .A(_55_), .Y(_56_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_57_) );
INVX1 INVX1_38 ( .A(_57_), .Y(_58_) );
NAND3X1 NAND3X1_13 ( .A(_56_), .B(_58_), .C(_51_), .Y(_59_) );
OAI21X1 OAI21X1_10 ( .A(_53_), .B(_54_), .C(_59_), .Y(w_C_16_) );
NOR2X1 NOR2X1_18 ( .A(_53_), .B(_54_), .Y(_60_) );
INVX1 INVX1_39 ( .A(_60_), .Y(_61_) );
AND2X2 AND2X2_12 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_62_) );
INVX1 INVX1_40 ( .A(_62_), .Y(_63_) );
NAND3X1 NAND3X1_14 ( .A(_61_), .B(_63_), .C(_59_), .Y(_64_) );
OAI21X1 OAI21X1_11 ( .A(i_add2[16]), .B(i_add1[16]), .C(_64_), .Y(_65_) );
INVX1 INVX1_41 ( .A(_65_), .Y(w_C_17_) );
INVX1 INVX1_42 ( .A(i_add2[17]), .Y(_66_) );
INVX1 INVX1_43 ( .A(i_add1[17]), .Y(_67_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_68_) );
INVX1 INVX1_44 ( .A(_68_), .Y(_69_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_70_) );
INVX1 INVX1_45 ( .A(_70_), .Y(_71_) );
NAND3X1 NAND3X1_15 ( .A(_69_), .B(_71_), .C(_64_), .Y(_72_) );
OAI21X1 OAI21X1_12 ( .A(_66_), .B(_67_), .C(_72_), .Y(w_C_18_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_73_) );
INVX1 INVX1_46 ( .A(_73_), .Y(_74_) );
NOR2X1 NOR2X1_22 ( .A(_66_), .B(_67_), .Y(_75_) );
INVX1 INVX1_47 ( .A(_75_), .Y(_76_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_77_) );
NAND3X1 NAND3X1_16 ( .A(_76_), .B(_77_), .C(_72_), .Y(_78_) );
AND2X2 AND2X2_13 ( .A(_78_), .B(_74_), .Y(w_C_19_) );
INVX1 INVX1_48 ( .A(i_add2[19]), .Y(_79_) );
INVX1 INVX1_49 ( .A(i_add1[19]), .Y(_80_) );
NAND2X1 NAND2X1_8 ( .A(_79_), .B(_80_), .Y(_81_) );
NAND3X1 NAND3X1_17 ( .A(_74_), .B(_81_), .C(_78_), .Y(_82_) );
OAI21X1 OAI21X1_13 ( .A(_79_), .B(_80_), .C(_82_), .Y(w_C_20_) );
INVX1 INVX1_50 ( .A(i_add2[20]), .Y(_83_) );
INVX1 INVX1_51 ( .A(i_add1[20]), .Y(_84_) );
NAND2X1 NAND2X1_9 ( .A(_83_), .B(_84_), .Y(_85_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_86_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_87_) );
NAND3X1 NAND3X1_18 ( .A(_86_), .B(_87_), .C(_82_), .Y(_88_) );
AND2X2 AND2X2_14 ( .A(_88_), .B(_85_), .Y(w_C_21_) );
INVX1 INVX1_52 ( .A(i_add2[21]), .Y(_89_) );
INVX1 INVX1_53 ( .A(i_add1[21]), .Y(_90_) );
NAND2X1 NAND2X1_12 ( .A(_89_), .B(_90_), .Y(_91_) );
NAND3X1 NAND3X1_19 ( .A(_85_), .B(_91_), .C(_88_), .Y(_92_) );
OAI21X1 OAI21X1_14 ( .A(_89_), .B(_90_), .C(_92_), .Y(w_C_22_) );
OR2X2 OR2X2_2 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_93_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_94_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_95_) );
NAND3X1 NAND3X1_20 ( .A(_94_), .B(_95_), .C(_92_), .Y(_96_) );
AND2X2 AND2X2_15 ( .A(_96_), .B(_93_), .Y(w_C_23_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_97_) );
OR2X2 OR2X2_3 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_98_) );
NAND3X1 NAND3X1_21 ( .A(_93_), .B(_98_), .C(_96_), .Y(_99_) );
NAND2X1 NAND2X1_16 ( .A(_97_), .B(_99_), .Y(w_C_24_) );
BUFX2 BUFX2_1 ( .A(_121__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_121__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_121__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_121__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_121__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_121__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_121__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_121__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_121__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_121__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_121__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_121__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_121__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_121__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_121__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_121__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_121__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_121__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_121__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_121__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_121__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_121__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_121__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_121__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(w_C_24_), .Y(o_result[24]) );
INVX1 INVX1_54 ( .A(w_C_4_), .Y(_125_) );
OR2X2 OR2X2_4 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_126_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_127_) );
NAND3X1 NAND3X1_22 ( .A(_125_), .B(_127_), .C(_126_), .Y(_128_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_122_) );
AND2X2 AND2X2_16 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_123_) );
OAI21X1 OAI21X1_15 ( .A(_122_), .B(_123_), .C(w_C_4_), .Y(_124_) );
NAND2X1 NAND2X1_18 ( .A(_124_), .B(_128_), .Y(_121__4_) );
INVX1 INVX1_55 ( .A(w_C_5_), .Y(_132_) );
OR2X2 OR2X2_5 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_133_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_134_) );
NAND3X1 NAND3X1_23 ( .A(_132_), .B(_134_), .C(_133_), .Y(_135_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_129_) );
AND2X2 AND2X2_17 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_130_) );
OAI21X1 OAI21X1_16 ( .A(_129_), .B(_130_), .C(w_C_5_), .Y(_131_) );
NAND2X1 NAND2X1_20 ( .A(_131_), .B(_135_), .Y(_121__5_) );
INVX1 INVX1_56 ( .A(w_C_6_), .Y(_139_) );
OR2X2 OR2X2_6 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_140_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_141_) );
NAND3X1 NAND3X1_24 ( .A(_139_), .B(_141_), .C(_140_), .Y(_142_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_136_) );
AND2X2 AND2X2_18 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_137_) );
OAI21X1 OAI21X1_17 ( .A(_136_), .B(_137_), .C(w_C_6_), .Y(_138_) );
NAND2X1 NAND2X1_22 ( .A(_138_), .B(_142_), .Y(_121__6_) );
INVX1 INVX1_57 ( .A(w_C_7_), .Y(_146_) );
OR2X2 OR2X2_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_147_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_148_) );
NAND3X1 NAND3X1_25 ( .A(_146_), .B(_148_), .C(_147_), .Y(_149_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_143_) );
AND2X2 AND2X2_19 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_144_) );
OAI21X1 OAI21X1_18 ( .A(_143_), .B(_144_), .C(w_C_7_), .Y(_145_) );
NAND2X1 NAND2X1_24 ( .A(_145_), .B(_149_), .Y(_121__7_) );
INVX1 INVX1_58 ( .A(w_C_8_), .Y(_153_) );
OR2X2 OR2X2_8 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_154_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_155_) );
NAND3X1 NAND3X1_26 ( .A(_153_), .B(_155_), .C(_154_), .Y(_156_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_150_) );
AND2X2 AND2X2_20 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_151_) );
OAI21X1 OAI21X1_19 ( .A(_150_), .B(_151_), .C(w_C_8_), .Y(_152_) );
NAND2X1 NAND2X1_26 ( .A(_152_), .B(_156_), .Y(_121__8_) );
INVX1 INVX1_59 ( .A(w_C_9_), .Y(_160_) );
OR2X2 OR2X2_9 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_161_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_162_) );
NAND3X1 NAND3X1_27 ( .A(_160_), .B(_162_), .C(_161_), .Y(_163_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_157_) );
AND2X2 AND2X2_21 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_158_) );
OAI21X1 OAI21X1_20 ( .A(_157_), .B(_158_), .C(w_C_9_), .Y(_159_) );
NAND2X1 NAND2X1_28 ( .A(_159_), .B(_163_), .Y(_121__9_) );
INVX1 INVX1_60 ( .A(w_C_10_), .Y(_167_) );
OR2X2 OR2X2_10 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_168_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_169_) );
NAND3X1 NAND3X1_28 ( .A(_167_), .B(_169_), .C(_168_), .Y(_170_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_164_) );
AND2X2 AND2X2_22 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_165_) );
OAI21X1 OAI21X1_21 ( .A(_164_), .B(_165_), .C(w_C_10_), .Y(_166_) );
NAND2X1 NAND2X1_30 ( .A(_166_), .B(_170_), .Y(_121__10_) );
INVX1 INVX1_61 ( .A(w_C_11_), .Y(_174_) );
OR2X2 OR2X2_11 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_175_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_176_) );
NAND3X1 NAND3X1_29 ( .A(_174_), .B(_176_), .C(_175_), .Y(_177_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_171_) );
AND2X2 AND2X2_23 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_172_) );
OAI21X1 OAI21X1_22 ( .A(_171_), .B(_172_), .C(w_C_11_), .Y(_173_) );
NAND2X1 NAND2X1_32 ( .A(_173_), .B(_177_), .Y(_121__11_) );
INVX1 INVX1_62 ( .A(w_C_12_), .Y(_181_) );
OR2X2 OR2X2_12 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_182_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_183_) );
NAND3X1 NAND3X1_30 ( .A(_181_), .B(_183_), .C(_182_), .Y(_184_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_178_) );
AND2X2 AND2X2_24 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_179_) );
OAI21X1 OAI21X1_23 ( .A(_178_), .B(_179_), .C(w_C_12_), .Y(_180_) );
NAND2X1 NAND2X1_34 ( .A(_180_), .B(_184_), .Y(_121__12_) );
INVX1 INVX1_63 ( .A(w_C_13_), .Y(_188_) );
OR2X2 OR2X2_13 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_189_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_190_) );
NAND3X1 NAND3X1_31 ( .A(_188_), .B(_190_), .C(_189_), .Y(_191_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_185_) );
AND2X2 AND2X2_25 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_186_) );
OAI21X1 OAI21X1_24 ( .A(_185_), .B(_186_), .C(w_C_13_), .Y(_187_) );
NAND2X1 NAND2X1_36 ( .A(_187_), .B(_191_), .Y(_121__13_) );
INVX1 INVX1_64 ( .A(w_C_14_), .Y(_195_) );
OR2X2 OR2X2_14 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_196_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_197_) );
NAND3X1 NAND3X1_32 ( .A(_195_), .B(_197_), .C(_196_), .Y(_198_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_192_) );
AND2X2 AND2X2_26 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_193_) );
OAI21X1 OAI21X1_25 ( .A(_192_), .B(_193_), .C(w_C_14_), .Y(_194_) );
NAND2X1 NAND2X1_38 ( .A(_194_), .B(_198_), .Y(_121__14_) );
INVX1 INVX1_65 ( .A(w_C_15_), .Y(_202_) );
OR2X2 OR2X2_15 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_203_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_204_) );
NAND3X1 NAND3X1_33 ( .A(_202_), .B(_204_), .C(_203_), .Y(_205_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_199_) );
AND2X2 AND2X2_27 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_200_) );
OAI21X1 OAI21X1_26 ( .A(_199_), .B(_200_), .C(w_C_15_), .Y(_201_) );
NAND2X1 NAND2X1_40 ( .A(_201_), .B(_205_), .Y(_121__15_) );
INVX1 INVX1_66 ( .A(w_C_16_), .Y(_209_) );
OR2X2 OR2X2_16 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_210_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_211_) );
NAND3X1 NAND3X1_34 ( .A(_209_), .B(_211_), .C(_210_), .Y(_212_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_206_) );
AND2X2 AND2X2_28 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_207_) );
OAI21X1 OAI21X1_27 ( .A(_206_), .B(_207_), .C(w_C_16_), .Y(_208_) );
NAND2X1 NAND2X1_42 ( .A(_208_), .B(_212_), .Y(_121__16_) );
INVX1 INVX1_67 ( .A(w_C_17_), .Y(_216_) );
OR2X2 OR2X2_17 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_217_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_218_) );
NAND3X1 NAND3X1_35 ( .A(_216_), .B(_218_), .C(_217_), .Y(_219_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_213_) );
AND2X2 AND2X2_29 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_214_) );
OAI21X1 OAI21X1_28 ( .A(_213_), .B(_214_), .C(w_C_17_), .Y(_215_) );
NAND2X1 NAND2X1_44 ( .A(_215_), .B(_219_), .Y(_121__17_) );
INVX1 INVX1_68 ( .A(w_C_18_), .Y(_223_) );
OR2X2 OR2X2_18 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_224_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_225_) );
NAND3X1 NAND3X1_36 ( .A(_223_), .B(_225_), .C(_224_), .Y(_226_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_220_) );
AND2X2 AND2X2_30 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_221_) );
OAI21X1 OAI21X1_29 ( .A(_220_), .B(_221_), .C(w_C_18_), .Y(_222_) );
NAND2X1 NAND2X1_46 ( .A(_222_), .B(_226_), .Y(_121__18_) );
INVX1 INVX1_69 ( .A(w_C_19_), .Y(_230_) );
OR2X2 OR2X2_19 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_231_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_232_) );
NAND3X1 NAND3X1_37 ( .A(_230_), .B(_232_), .C(_231_), .Y(_233_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_227_) );
AND2X2 AND2X2_31 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_228_) );
OAI21X1 OAI21X1_30 ( .A(_227_), .B(_228_), .C(w_C_19_), .Y(_229_) );
NAND2X1 NAND2X1_48 ( .A(_229_), .B(_233_), .Y(_121__19_) );
INVX1 INVX1_70 ( .A(w_C_20_), .Y(_237_) );
OR2X2 OR2X2_20 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_238_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_239_) );
NAND3X1 NAND3X1_38 ( .A(_237_), .B(_239_), .C(_238_), .Y(_240_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_234_) );
AND2X2 AND2X2_32 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_235_) );
OAI21X1 OAI21X1_31 ( .A(_234_), .B(_235_), .C(w_C_20_), .Y(_236_) );
NAND2X1 NAND2X1_50 ( .A(_236_), .B(_240_), .Y(_121__20_) );
INVX1 INVX1_71 ( .A(w_C_21_), .Y(_244_) );
OR2X2 OR2X2_21 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_245_) );
NAND2X1 NAND2X1_51 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_246_) );
NAND3X1 NAND3X1_39 ( .A(_244_), .B(_246_), .C(_245_), .Y(_247_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_241_) );
AND2X2 AND2X2_33 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_242_) );
OAI21X1 OAI21X1_32 ( .A(_241_), .B(_242_), .C(w_C_21_), .Y(_243_) );
NAND2X1 NAND2X1_52 ( .A(_243_), .B(_247_), .Y(_121__21_) );
INVX1 INVX1_72 ( .A(w_C_22_), .Y(_251_) );
OR2X2 OR2X2_22 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_252_) );
NAND2X1 NAND2X1_53 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_253_) );
NAND3X1 NAND3X1_40 ( .A(_251_), .B(_253_), .C(_252_), .Y(_254_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_248_) );
AND2X2 AND2X2_34 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_249_) );
OAI21X1 OAI21X1_33 ( .A(_248_), .B(_249_), .C(w_C_22_), .Y(_250_) );
NAND2X1 NAND2X1_54 ( .A(_250_), .B(_254_), .Y(_121__22_) );
INVX1 INVX1_73 ( .A(w_C_23_), .Y(_258_) );
OR2X2 OR2X2_23 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_259_) );
NAND2X1 NAND2X1_55 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_260_) );
NAND3X1 NAND3X1_41 ( .A(_258_), .B(_260_), .C(_259_), .Y(_261_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_255_) );
AND2X2 AND2X2_35 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_256_) );
OAI21X1 OAI21X1_34 ( .A(_255_), .B(_256_), .C(w_C_23_), .Y(_257_) );
NAND2X1 NAND2X1_56 ( .A(_257_), .B(_261_), .Y(_121__23_) );
INVX1 INVX1_74 ( .A(gnd), .Y(_265_) );
OR2X2 OR2X2_24 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_266_) );
NAND2X1 NAND2X1_57 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_267_) );
NAND3X1 NAND3X1_42 ( .A(_265_), .B(_267_), .C(_266_), .Y(_268_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_262_) );
AND2X2 AND2X2_36 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_263_) );
OAI21X1 OAI21X1_35 ( .A(_262_), .B(_263_), .C(gnd), .Y(_264_) );
NAND2X1 NAND2X1_58 ( .A(_264_), .B(_268_), .Y(_121__0_) );
INVX1 INVX1_75 ( .A(w_C_1_), .Y(_272_) );
OR2X2 OR2X2_25 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_273_) );
NAND2X1 NAND2X1_59 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_274_) );
NAND3X1 NAND3X1_43 ( .A(_272_), .B(_274_), .C(_273_), .Y(_275_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_269_) );
AND2X2 AND2X2_37 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_270_) );
OAI21X1 OAI21X1_36 ( .A(_269_), .B(_270_), .C(w_C_1_), .Y(_271_) );
NAND2X1 NAND2X1_60 ( .A(_271_), .B(_275_), .Y(_121__1_) );
INVX1 INVX1_76 ( .A(w_C_2_), .Y(_279_) );
OR2X2 OR2X2_26 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_280_) );
NAND2X1 NAND2X1_61 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_281_) );
NAND3X1 NAND3X1_44 ( .A(_279_), .B(_281_), .C(_280_), .Y(_282_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_276_) );
AND2X2 AND2X2_38 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_277_) );
OAI21X1 OAI21X1_37 ( .A(_276_), .B(_277_), .C(w_C_2_), .Y(_278_) );
NAND2X1 NAND2X1_62 ( .A(_278_), .B(_282_), .Y(_121__2_) );
INVX1 INVX1_77 ( .A(w_C_3_), .Y(_286_) );
OR2X2 OR2X2_27 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_287_) );
NAND2X1 NAND2X1_63 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_288_) );
NAND3X1 NAND3X1_45 ( .A(_286_), .B(_288_), .C(_287_), .Y(_289_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_283_) );
AND2X2 AND2X2_39 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_284_) );
OAI21X1 OAI21X1_38 ( .A(_283_), .B(_284_), .C(w_C_3_), .Y(_285_) );
NAND2X1 NAND2X1_64 ( .A(_285_), .B(_289_), .Y(_121__3_) );
BUFX2 BUFX2_26 ( .A(w_C_24_), .Y(_121__24_) );
BUFX2 BUFX2_27 ( .A(gnd), .Y(w_C_0_) );
endmodule
