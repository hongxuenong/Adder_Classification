module CSkipA_45bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output cout;

NOR2X1 NOR2X1_1 ( .A(_379_), .B(_380_), .Y(_381_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_382_) );
NAND2X1 NAND2X1_1 ( .A(_381_), .B(_382_), .Y(_383_) );
NOR2X1 NOR2X1_2 ( .A(_378_), .B(_383_), .Y(_24_) );
INVX1 INVX1_1 ( .A(_22_), .Y(_384_) );
NAND2X1 NAND2X1_2 ( .A(1'b0), .B(_24_), .Y(_385_) );
OAI21X1 OAI21X1_1 ( .A(_24_), .B(_384_), .C(_385_), .Y(w_cout_8_) );
INVX1 INVX1_2 ( .A(w_cout_8_), .Y(_389_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_390_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_391_) );
NAND3X1 NAND3X1_1 ( .A(_389_), .B(_391_), .C(_390_), .Y(_392_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_386_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_387_) );
OAI21X1 OAI21X1_2 ( .A(_386_), .B(_387_), .C(w_cout_8_), .Y(_388_) );
NAND2X1 NAND2X1_4 ( .A(_388_), .B(_392_), .Y(_0__32_) );
OAI21X1 OAI21X1_3 ( .A(_389_), .B(_386_), .C(_391_), .Y(_26__1_) );
INVX1 INVX1_3 ( .A(_26__3_), .Y(_396_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_397_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_398_) );
NAND3X1 NAND3X1_2 ( .A(_396_), .B(_398_), .C(_397_), .Y(_399_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_393_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_394_) );
OAI21X1 OAI21X1_4 ( .A(_393_), .B(_394_), .C(_26__3_), .Y(_395_) );
NAND2X1 NAND2X1_6 ( .A(_395_), .B(_399_), .Y(_0__35_) );
OAI21X1 OAI21X1_5 ( .A(_396_), .B(_393_), .C(_398_), .Y(_25_) );
INVX1 INVX1_4 ( .A(_26__1_), .Y(_403_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_404_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_405_) );
NAND3X1 NAND3X1_3 ( .A(_403_), .B(_405_), .C(_404_), .Y(_406_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_400_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_401_) );
OAI21X1 OAI21X1_6 ( .A(_400_), .B(_401_), .C(_26__1_), .Y(_402_) );
NAND2X1 NAND2X1_8 ( .A(_402_), .B(_406_), .Y(_0__33_) );
OAI21X1 OAI21X1_7 ( .A(_403_), .B(_400_), .C(_405_), .Y(_26__2_) );
INVX1 INVX1_5 ( .A(_26__2_), .Y(_410_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_411_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_412_) );
NAND3X1 NAND3X1_4 ( .A(_410_), .B(_412_), .C(_411_), .Y(_413_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_407_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_408_) );
OAI21X1 OAI21X1_8 ( .A(_407_), .B(_408_), .C(_26__2_), .Y(_409_) );
NAND2X1 NAND2X1_10 ( .A(_409_), .B(_413_), .Y(_0__34_) );
OAI21X1 OAI21X1_9 ( .A(_410_), .B(_407_), .C(_412_), .Y(_26__3_) );
INVX1 INVX1_6 ( .A(i_add_term1[32]), .Y(_414_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[32]), .B(_414_), .Y(_415_) );
INVX1 INVX1_7 ( .A(i_add_term2[32]), .Y(_416_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term1[32]), .B(_416_), .Y(_417_) );
INVX1 INVX1_8 ( .A(i_add_term1[33]), .Y(_418_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[33]), .B(_418_), .Y(_419_) );
INVX1 INVX1_9 ( .A(i_add_term2[33]), .Y(_420_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term1[33]), .B(_420_), .Y(_421_) );
OAI22X1 OAI22X1_1 ( .A(_415_), .B(_417_), .C(_419_), .D(_421_), .Y(_422_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_423_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_424_) );
NOR2X1 NOR2X1_12 ( .A(_423_), .B(_424_), .Y(_425_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_426_) );
NAND2X1 NAND2X1_11 ( .A(_425_), .B(_426_), .Y(_427_) );
NOR2X1 NOR2X1_13 ( .A(_422_), .B(_427_), .Y(_27_) );
INVX1 INVX1_10 ( .A(_25_), .Y(_428_) );
NAND2X1 NAND2X1_12 ( .A(1'b0), .B(_27_), .Y(_429_) );
OAI21X1 OAI21X1_10 ( .A(_27_), .B(_428_), .C(_429_), .Y(w_cout_9_) );
INVX1 INVX1_11 ( .A(w_cout_9_), .Y(_433_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_434_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_435_) );
NAND3X1 NAND3X1_5 ( .A(_433_), .B(_435_), .C(_434_), .Y(_436_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_430_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_431_) );
OAI21X1 OAI21X1_11 ( .A(_430_), .B(_431_), .C(w_cout_9_), .Y(_432_) );
NAND2X1 NAND2X1_14 ( .A(_432_), .B(_436_), .Y(_0__36_) );
OAI21X1 OAI21X1_12 ( .A(_433_), .B(_430_), .C(_435_), .Y(_29__1_) );
INVX1 INVX1_12 ( .A(_29__3_), .Y(_440_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_441_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_442_) );
NAND3X1 NAND3X1_6 ( .A(_440_), .B(_442_), .C(_441_), .Y(_443_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_437_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_438_) );
OAI21X1 OAI21X1_13 ( .A(_437_), .B(_438_), .C(_29__3_), .Y(_439_) );
NAND2X1 NAND2X1_16 ( .A(_439_), .B(_443_), .Y(_0__39_) );
OAI21X1 OAI21X1_14 ( .A(_440_), .B(_437_), .C(_442_), .Y(_28_) );
INVX1 INVX1_13 ( .A(_29__1_), .Y(_447_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_448_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_449_) );
NAND3X1 NAND3X1_7 ( .A(_447_), .B(_449_), .C(_448_), .Y(_450_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_444_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_445_) );
OAI21X1 OAI21X1_15 ( .A(_444_), .B(_445_), .C(_29__1_), .Y(_446_) );
NAND2X1 NAND2X1_18 ( .A(_446_), .B(_450_), .Y(_0__37_) );
OAI21X1 OAI21X1_16 ( .A(_447_), .B(_444_), .C(_449_), .Y(_29__2_) );
INVX1 INVX1_14 ( .A(_29__2_), .Y(_454_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_455_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_456_) );
NAND3X1 NAND3X1_8 ( .A(_454_), .B(_456_), .C(_455_), .Y(_457_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_451_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_452_) );
OAI21X1 OAI21X1_17 ( .A(_451_), .B(_452_), .C(_29__2_), .Y(_453_) );
NAND2X1 NAND2X1_20 ( .A(_453_), .B(_457_), .Y(_0__38_) );
OAI21X1 OAI21X1_18 ( .A(_454_), .B(_451_), .C(_456_), .Y(_29__3_) );
INVX1 INVX1_15 ( .A(i_add_term1[36]), .Y(_458_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[36]), .B(_458_), .Y(_459_) );
INVX1 INVX1_16 ( .A(i_add_term2[36]), .Y(_460_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term1[36]), .B(_460_), .Y(_461_) );
INVX1 INVX1_17 ( .A(i_add_term1[37]), .Y(_462_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[37]), .B(_462_), .Y(_463_) );
INVX1 INVX1_18 ( .A(i_add_term2[37]), .Y(_464_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term1[37]), .B(_464_), .Y(_465_) );
OAI22X1 OAI22X1_2 ( .A(_459_), .B(_461_), .C(_463_), .D(_465_), .Y(_466_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_467_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_468_) );
NOR2X1 NOR2X1_23 ( .A(_467_), .B(_468_), .Y(_469_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_470_) );
NAND2X1 NAND2X1_21 ( .A(_469_), .B(_470_), .Y(_471_) );
NOR2X1 NOR2X1_24 ( .A(_466_), .B(_471_), .Y(_30_) );
INVX1 INVX1_19 ( .A(_28_), .Y(_472_) );
NAND2X1 NAND2X1_22 ( .A(1'b0), .B(_30_), .Y(_473_) );
OAI21X1 OAI21X1_19 ( .A(_30_), .B(_472_), .C(_473_), .Y(w_cout_10_) );
INVX1 INVX1_20 ( .A(w_cout_10_), .Y(_477_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_478_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_479_) );
NAND3X1 NAND3X1_9 ( .A(_477_), .B(_479_), .C(_478_), .Y(_480_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_474_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_475_) );
OAI21X1 OAI21X1_20 ( .A(_474_), .B(_475_), .C(w_cout_10_), .Y(_476_) );
NAND2X1 NAND2X1_24 ( .A(_476_), .B(_480_), .Y(_0__40_) );
OAI21X1 OAI21X1_21 ( .A(_477_), .B(_474_), .C(_479_), .Y(_32__1_) );
INVX1 INVX1_21 ( .A(_32__3_), .Y(_484_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_485_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_486_) );
NAND3X1 NAND3X1_10 ( .A(_484_), .B(_486_), .C(_485_), .Y(_487_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_481_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_482_) );
OAI21X1 OAI21X1_22 ( .A(_481_), .B(_482_), .C(_32__3_), .Y(_483_) );
NAND2X1 NAND2X1_26 ( .A(_483_), .B(_487_), .Y(_0__43_) );
OAI21X1 OAI21X1_23 ( .A(_484_), .B(_481_), .C(_486_), .Y(_31_) );
INVX1 INVX1_22 ( .A(_32__1_), .Y(_491_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_492_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_493_) );
NAND3X1 NAND3X1_11 ( .A(_491_), .B(_493_), .C(_492_), .Y(_494_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_488_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_489_) );
OAI21X1 OAI21X1_24 ( .A(_488_), .B(_489_), .C(_32__1_), .Y(_490_) );
NAND2X1 NAND2X1_28 ( .A(_490_), .B(_494_), .Y(_0__41_) );
OAI21X1 OAI21X1_25 ( .A(_491_), .B(_488_), .C(_493_), .Y(_32__2_) );
INVX1 INVX1_23 ( .A(_32__2_), .Y(_498_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_499_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_500_) );
NAND3X1 NAND3X1_12 ( .A(_498_), .B(_500_), .C(_499_), .Y(_501_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_495_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_496_) );
OAI21X1 OAI21X1_26 ( .A(_495_), .B(_496_), .C(_32__2_), .Y(_497_) );
NAND2X1 NAND2X1_30 ( .A(_497_), .B(_501_), .Y(_0__42_) );
OAI21X1 OAI21X1_27 ( .A(_498_), .B(_495_), .C(_500_), .Y(_32__3_) );
INVX1 INVX1_24 ( .A(i_add_term1[40]), .Y(_502_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[40]), .B(_502_), .Y(_503_) );
INVX1 INVX1_25 ( .A(i_add_term2[40]), .Y(_504_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term1[40]), .B(_504_), .Y(_505_) );
INVX1 INVX1_26 ( .A(i_add_term1[41]), .Y(_506_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[41]), .B(_506_), .Y(_507_) );
INVX1 INVX1_27 ( .A(i_add_term2[41]), .Y(_508_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term1[41]), .B(_508_), .Y(_509_) );
OAI22X1 OAI22X1_3 ( .A(_503_), .B(_505_), .C(_507_), .D(_509_), .Y(_510_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_511_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_512_) );
NOR2X1 NOR2X1_34 ( .A(_511_), .B(_512_), .Y(_513_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_514_) );
NAND2X1 NAND2X1_31 ( .A(_513_), .B(_514_), .Y(_515_) );
NOR2X1 NOR2X1_35 ( .A(_510_), .B(_515_), .Y(_33_) );
INVX1 INVX1_28 ( .A(_31_), .Y(_516_) );
NAND2X1 NAND2X1_32 ( .A(1'b0), .B(_33_), .Y(_517_) );
OAI21X1 OAI21X1_28 ( .A(_33_), .B(_516_), .C(_517_), .Y(cskip1_inst_cin) );
INVX1 INVX1_29 ( .A(cskip1_inst_cin), .Y(_521_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_522_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_523_) );
NAND3X1 NAND3X1_13 ( .A(_521_), .B(_523_), .C(_522_), .Y(_524_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_518_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_519_) );
OAI21X1 OAI21X1_29 ( .A(_518_), .B(_519_), .C(cskip1_inst_cin), .Y(_520_) );
NAND2X1 NAND2X1_34 ( .A(_520_), .B(_524_), .Y(cskip1_inst_rca0_fa0_o_sum) );
OAI21X1 OAI21X1_30 ( .A(_521_), .B(_518_), .C(_523_), .Y(cskip1_inst_cout0) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_525_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_526_) );
NOR2X1 NOR2X1_38 ( .A(_525_), .B(_526_), .Y(cskip1_inst_skip0_P) );
INVX1 INVX1_30 ( .A(cskip1_inst_cout0), .Y(_527_) );
NAND2X1 NAND2X1_35 ( .A(1'b0), .B(cskip1_inst_skip0_P), .Y(_528_) );
OAI21X1 OAI21X1_31 ( .A(cskip1_inst_skip0_P), .B(_527_), .C(_528_), .Y(w_cout_12_) );
BUFX2 BUFX2_1 ( .A(w_cout_12_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(cskip1_inst_rca0_fa0_o_sum), .Y(sum[44]) );
INVX1 INVX1_31 ( .A(1'b0), .Y(_37_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_38_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_39_) );
NAND3X1 NAND3X1_14 ( .A(_37_), .B(_39_), .C(_38_), .Y(_40_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_34_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_35_) );
OAI21X1 OAI21X1_32 ( .A(_34_), .B(_35_), .C(1'b0), .Y(_36_) );
NAND2X1 NAND2X1_37 ( .A(_36_), .B(_40_), .Y(_0__0_) );
OAI21X1 OAI21X1_33 ( .A(_37_), .B(_34_), .C(_39_), .Y(_2__1_) );
INVX1 INVX1_32 ( .A(_2__3_), .Y(_44_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_45_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_46_) );
NAND3X1 NAND3X1_15 ( .A(_44_), .B(_46_), .C(_45_), .Y(_47_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_41_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_42_) );
OAI21X1 OAI21X1_34 ( .A(_41_), .B(_42_), .C(_2__3_), .Y(_43_) );
NAND2X1 NAND2X1_39 ( .A(_43_), .B(_47_), .Y(_0__3_) );
OAI21X1 OAI21X1_35 ( .A(_44_), .B(_41_), .C(_46_), .Y(_1_) );
INVX1 INVX1_33 ( .A(_2__1_), .Y(_51_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_52_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_53_) );
NAND3X1 NAND3X1_16 ( .A(_51_), .B(_53_), .C(_52_), .Y(_54_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_48_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_49_) );
OAI21X1 OAI21X1_36 ( .A(_48_), .B(_49_), .C(_2__1_), .Y(_50_) );
NAND2X1 NAND2X1_41 ( .A(_50_), .B(_54_), .Y(_0__1_) );
OAI21X1 OAI21X1_37 ( .A(_51_), .B(_48_), .C(_53_), .Y(_2__2_) );
INVX1 INVX1_34 ( .A(_2__2_), .Y(_58_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_59_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_60_) );
NAND3X1 NAND3X1_17 ( .A(_58_), .B(_60_), .C(_59_), .Y(_61_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_55_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_56_) );
OAI21X1 OAI21X1_38 ( .A(_55_), .B(_56_), .C(_2__2_), .Y(_57_) );
NAND2X1 NAND2X1_43 ( .A(_57_), .B(_61_), .Y(_0__2_) );
OAI21X1 OAI21X1_39 ( .A(_58_), .B(_55_), .C(_60_), .Y(_2__3_) );
INVX1 INVX1_35 ( .A(i_add_term1[0]), .Y(_62_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[0]), .B(_62_), .Y(_63_) );
INVX1 INVX1_36 ( .A(i_add_term2[0]), .Y(_64_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term1[0]), .B(_64_), .Y(_65_) );
INVX1 INVX1_37 ( .A(i_add_term1[1]), .Y(_66_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[1]), .B(_66_), .Y(_67_) );
INVX1 INVX1_38 ( .A(i_add_term2[1]), .Y(_68_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term1[1]), .B(_68_), .Y(_69_) );
OAI22X1 OAI22X1_4 ( .A(_63_), .B(_65_), .C(_67_), .D(_69_), .Y(_70_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_71_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_72_) );
NOR2X1 NOR2X1_48 ( .A(_71_), .B(_72_), .Y(_73_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_74_) );
NAND2X1 NAND2X1_44 ( .A(_73_), .B(_74_), .Y(_75_) );
NOR2X1 NOR2X1_49 ( .A(_70_), .B(_75_), .Y(_3_) );
INVX1 INVX1_39 ( .A(_1_), .Y(_76_) );
NAND2X1 NAND2X1_45 ( .A(1'b0), .B(_3_), .Y(_77_) );
OAI21X1 OAI21X1_40 ( .A(_3_), .B(_76_), .C(_77_), .Y(w_cout_1_) );
INVX1 INVX1_40 ( .A(w_cout_1_), .Y(_81_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_82_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_83_) );
NAND3X1 NAND3X1_18 ( .A(_81_), .B(_83_), .C(_82_), .Y(_84_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_78_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_79_) );
OAI21X1 OAI21X1_41 ( .A(_78_), .B(_79_), .C(w_cout_1_), .Y(_80_) );
NAND2X1 NAND2X1_47 ( .A(_80_), .B(_84_), .Y(_0__4_) );
OAI21X1 OAI21X1_42 ( .A(_81_), .B(_78_), .C(_83_), .Y(_5__1_) );
INVX1 INVX1_41 ( .A(_5__3_), .Y(_88_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_89_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_90_) );
NAND3X1 NAND3X1_19 ( .A(_88_), .B(_90_), .C(_89_), .Y(_91_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_85_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_86_) );
OAI21X1 OAI21X1_43 ( .A(_85_), .B(_86_), .C(_5__3_), .Y(_87_) );
NAND2X1 NAND2X1_49 ( .A(_87_), .B(_91_), .Y(_0__7_) );
OAI21X1 OAI21X1_44 ( .A(_88_), .B(_85_), .C(_90_), .Y(_4_) );
INVX1 INVX1_42 ( .A(_5__1_), .Y(_95_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_96_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_97_) );
NAND3X1 NAND3X1_20 ( .A(_95_), .B(_97_), .C(_96_), .Y(_98_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_92_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_93_) );
OAI21X1 OAI21X1_45 ( .A(_92_), .B(_93_), .C(_5__1_), .Y(_94_) );
NAND2X1 NAND2X1_51 ( .A(_94_), .B(_98_), .Y(_0__5_) );
OAI21X1 OAI21X1_46 ( .A(_95_), .B(_92_), .C(_97_), .Y(_5__2_) );
INVX1 INVX1_43 ( .A(_5__2_), .Y(_102_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_103_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_104_) );
NAND3X1 NAND3X1_21 ( .A(_102_), .B(_104_), .C(_103_), .Y(_105_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_99_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_100_) );
OAI21X1 OAI21X1_47 ( .A(_99_), .B(_100_), .C(_5__2_), .Y(_101_) );
NAND2X1 NAND2X1_53 ( .A(_101_), .B(_105_), .Y(_0__6_) );
OAI21X1 OAI21X1_48 ( .A(_102_), .B(_99_), .C(_104_), .Y(_5__3_) );
INVX1 INVX1_44 ( .A(i_add_term1[4]), .Y(_106_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[4]), .B(_106_), .Y(_107_) );
INVX1 INVX1_45 ( .A(i_add_term2[4]), .Y(_108_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term1[4]), .B(_108_), .Y(_109_) );
INVX1 INVX1_46 ( .A(i_add_term1[5]), .Y(_110_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[5]), .B(_110_), .Y(_111_) );
INVX1 INVX1_47 ( .A(i_add_term2[5]), .Y(_112_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term1[5]), .B(_112_), .Y(_113_) );
OAI22X1 OAI22X1_5 ( .A(_107_), .B(_109_), .C(_111_), .D(_113_), .Y(_114_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_115_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_116_) );
NOR2X1 NOR2X1_59 ( .A(_115_), .B(_116_), .Y(_117_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_118_) );
NAND2X1 NAND2X1_54 ( .A(_117_), .B(_118_), .Y(_119_) );
NOR2X1 NOR2X1_60 ( .A(_114_), .B(_119_), .Y(_6_) );
INVX1 INVX1_48 ( .A(_4_), .Y(_120_) );
NAND2X1 NAND2X1_55 ( .A(1'b0), .B(_6_), .Y(_121_) );
OAI21X1 OAI21X1_49 ( .A(_6_), .B(_120_), .C(_121_), .Y(w_cout_2_) );
INVX1 INVX1_49 ( .A(w_cout_2_), .Y(_125_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_126_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_127_) );
NAND3X1 NAND3X1_22 ( .A(_125_), .B(_127_), .C(_126_), .Y(_128_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_122_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_123_) );
OAI21X1 OAI21X1_50 ( .A(_122_), .B(_123_), .C(w_cout_2_), .Y(_124_) );
NAND2X1 NAND2X1_57 ( .A(_124_), .B(_128_), .Y(_0__8_) );
OAI21X1 OAI21X1_51 ( .A(_125_), .B(_122_), .C(_127_), .Y(_8__1_) );
INVX1 INVX1_50 ( .A(_8__3_), .Y(_132_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_133_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_134_) );
NAND3X1 NAND3X1_23 ( .A(_132_), .B(_134_), .C(_133_), .Y(_135_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_129_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_130_) );
OAI21X1 OAI21X1_52 ( .A(_129_), .B(_130_), .C(_8__3_), .Y(_131_) );
NAND2X1 NAND2X1_59 ( .A(_131_), .B(_135_), .Y(_0__11_) );
OAI21X1 OAI21X1_53 ( .A(_132_), .B(_129_), .C(_134_), .Y(_7_) );
INVX1 INVX1_51 ( .A(_8__1_), .Y(_139_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_140_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_141_) );
NAND3X1 NAND3X1_24 ( .A(_139_), .B(_141_), .C(_140_), .Y(_142_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_136_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_137_) );
OAI21X1 OAI21X1_54 ( .A(_136_), .B(_137_), .C(_8__1_), .Y(_138_) );
NAND2X1 NAND2X1_61 ( .A(_138_), .B(_142_), .Y(_0__9_) );
OAI21X1 OAI21X1_55 ( .A(_139_), .B(_136_), .C(_141_), .Y(_8__2_) );
INVX1 INVX1_52 ( .A(_8__2_), .Y(_146_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_147_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_148_) );
NAND3X1 NAND3X1_25 ( .A(_146_), .B(_148_), .C(_147_), .Y(_149_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_143_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_144_) );
OAI21X1 OAI21X1_56 ( .A(_143_), .B(_144_), .C(_8__2_), .Y(_145_) );
NAND2X1 NAND2X1_63 ( .A(_145_), .B(_149_), .Y(_0__10_) );
OAI21X1 OAI21X1_57 ( .A(_146_), .B(_143_), .C(_148_), .Y(_8__3_) );
INVX1 INVX1_53 ( .A(i_add_term1[8]), .Y(_150_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[8]), .B(_150_), .Y(_151_) );
INVX1 INVX1_54 ( .A(i_add_term2[8]), .Y(_152_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term1[8]), .B(_152_), .Y(_153_) );
INVX1 INVX1_55 ( .A(i_add_term1[9]), .Y(_154_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[9]), .B(_154_), .Y(_155_) );
INVX1 INVX1_56 ( .A(i_add_term2[9]), .Y(_156_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term1[9]), .B(_156_), .Y(_157_) );
OAI22X1 OAI22X1_6 ( .A(_151_), .B(_153_), .C(_155_), .D(_157_), .Y(_158_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_159_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_160_) );
NOR2X1 NOR2X1_70 ( .A(_159_), .B(_160_), .Y(_161_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_162_) );
NAND2X1 NAND2X1_64 ( .A(_161_), .B(_162_), .Y(_163_) );
NOR2X1 NOR2X1_71 ( .A(_158_), .B(_163_), .Y(_9_) );
INVX1 INVX1_57 ( .A(_7_), .Y(_164_) );
NAND2X1 NAND2X1_65 ( .A(1'b0), .B(_9_), .Y(_165_) );
OAI21X1 OAI21X1_58 ( .A(_9_), .B(_164_), .C(_165_), .Y(w_cout_3_) );
INVX1 INVX1_58 ( .A(w_cout_3_), .Y(_169_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_170_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_171_) );
NAND3X1 NAND3X1_26 ( .A(_169_), .B(_171_), .C(_170_), .Y(_172_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_166_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_167_) );
OAI21X1 OAI21X1_59 ( .A(_166_), .B(_167_), .C(w_cout_3_), .Y(_168_) );
NAND2X1 NAND2X1_67 ( .A(_168_), .B(_172_), .Y(_0__12_) );
OAI21X1 OAI21X1_60 ( .A(_169_), .B(_166_), .C(_171_), .Y(_11__1_) );
INVX1 INVX1_59 ( .A(_11__3_), .Y(_176_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_177_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_178_) );
NAND3X1 NAND3X1_27 ( .A(_176_), .B(_178_), .C(_177_), .Y(_179_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_173_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_174_) );
OAI21X1 OAI21X1_61 ( .A(_173_), .B(_174_), .C(_11__3_), .Y(_175_) );
NAND2X1 NAND2X1_69 ( .A(_175_), .B(_179_), .Y(_0__15_) );
OAI21X1 OAI21X1_62 ( .A(_176_), .B(_173_), .C(_178_), .Y(_10_) );
INVX1 INVX1_60 ( .A(_11__1_), .Y(_183_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_184_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_185_) );
NAND3X1 NAND3X1_28 ( .A(_183_), .B(_185_), .C(_184_), .Y(_186_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_180_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_181_) );
OAI21X1 OAI21X1_63 ( .A(_180_), .B(_181_), .C(_11__1_), .Y(_182_) );
NAND2X1 NAND2X1_71 ( .A(_182_), .B(_186_), .Y(_0__13_) );
OAI21X1 OAI21X1_64 ( .A(_183_), .B(_180_), .C(_185_), .Y(_11__2_) );
INVX1 INVX1_61 ( .A(_11__2_), .Y(_190_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_191_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_192_) );
NAND3X1 NAND3X1_29 ( .A(_190_), .B(_192_), .C(_191_), .Y(_193_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_187_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_188_) );
OAI21X1 OAI21X1_65 ( .A(_187_), .B(_188_), .C(_11__2_), .Y(_189_) );
NAND2X1 NAND2X1_73 ( .A(_189_), .B(_193_), .Y(_0__14_) );
OAI21X1 OAI21X1_66 ( .A(_190_), .B(_187_), .C(_192_), .Y(_11__3_) );
INVX1 INVX1_62 ( .A(i_add_term1[12]), .Y(_194_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[12]), .B(_194_), .Y(_195_) );
INVX1 INVX1_63 ( .A(i_add_term2[12]), .Y(_196_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term1[12]), .B(_196_), .Y(_197_) );
INVX1 INVX1_64 ( .A(i_add_term1[13]), .Y(_198_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[13]), .B(_198_), .Y(_199_) );
INVX1 INVX1_65 ( .A(i_add_term2[13]), .Y(_200_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term1[13]), .B(_200_), .Y(_201_) );
OAI22X1 OAI22X1_7 ( .A(_195_), .B(_197_), .C(_199_), .D(_201_), .Y(_202_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_203_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_204_) );
NOR2X1 NOR2X1_81 ( .A(_203_), .B(_204_), .Y(_205_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_206_) );
NAND2X1 NAND2X1_74 ( .A(_205_), .B(_206_), .Y(_207_) );
NOR2X1 NOR2X1_82 ( .A(_202_), .B(_207_), .Y(_12_) );
INVX1 INVX1_66 ( .A(_10_), .Y(_208_) );
NAND2X1 NAND2X1_75 ( .A(1'b0), .B(_12_), .Y(_209_) );
OAI21X1 OAI21X1_67 ( .A(_12_), .B(_208_), .C(_209_), .Y(w_cout_4_) );
INVX1 INVX1_67 ( .A(w_cout_4_), .Y(_213_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_214_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_215_) );
NAND3X1 NAND3X1_30 ( .A(_213_), .B(_215_), .C(_214_), .Y(_216_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_210_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_211_) );
OAI21X1 OAI21X1_68 ( .A(_210_), .B(_211_), .C(w_cout_4_), .Y(_212_) );
NAND2X1 NAND2X1_77 ( .A(_212_), .B(_216_), .Y(_0__16_) );
OAI21X1 OAI21X1_69 ( .A(_213_), .B(_210_), .C(_215_), .Y(_14__1_) );
INVX1 INVX1_68 ( .A(_14__3_), .Y(_220_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_221_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_222_) );
NAND3X1 NAND3X1_31 ( .A(_220_), .B(_222_), .C(_221_), .Y(_223_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_217_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_218_) );
OAI21X1 OAI21X1_70 ( .A(_217_), .B(_218_), .C(_14__3_), .Y(_219_) );
NAND2X1 NAND2X1_79 ( .A(_219_), .B(_223_), .Y(_0__19_) );
OAI21X1 OAI21X1_71 ( .A(_220_), .B(_217_), .C(_222_), .Y(_13_) );
INVX1 INVX1_69 ( .A(_14__1_), .Y(_227_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_228_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_229_) );
NAND3X1 NAND3X1_32 ( .A(_227_), .B(_229_), .C(_228_), .Y(_230_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_224_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_225_) );
OAI21X1 OAI21X1_72 ( .A(_224_), .B(_225_), .C(_14__1_), .Y(_226_) );
NAND2X1 NAND2X1_81 ( .A(_226_), .B(_230_), .Y(_0__17_) );
OAI21X1 OAI21X1_73 ( .A(_227_), .B(_224_), .C(_229_), .Y(_14__2_) );
INVX1 INVX1_70 ( .A(_14__2_), .Y(_234_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_235_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_236_) );
NAND3X1 NAND3X1_33 ( .A(_234_), .B(_236_), .C(_235_), .Y(_237_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_231_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_232_) );
OAI21X1 OAI21X1_74 ( .A(_231_), .B(_232_), .C(_14__2_), .Y(_233_) );
NAND2X1 NAND2X1_83 ( .A(_233_), .B(_237_), .Y(_0__18_) );
OAI21X1 OAI21X1_75 ( .A(_234_), .B(_231_), .C(_236_), .Y(_14__3_) );
INVX1 INVX1_71 ( .A(i_add_term1[16]), .Y(_238_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[16]), .B(_238_), .Y(_239_) );
INVX1 INVX1_72 ( .A(i_add_term2[16]), .Y(_240_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term1[16]), .B(_240_), .Y(_241_) );
INVX1 INVX1_73 ( .A(i_add_term1[17]), .Y(_242_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[17]), .B(_242_), .Y(_243_) );
INVX1 INVX1_74 ( .A(i_add_term2[17]), .Y(_244_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term1[17]), .B(_244_), .Y(_245_) );
OAI22X1 OAI22X1_8 ( .A(_239_), .B(_241_), .C(_243_), .D(_245_), .Y(_246_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_247_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_248_) );
NOR2X1 NOR2X1_92 ( .A(_247_), .B(_248_), .Y(_249_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_250_) );
NAND2X1 NAND2X1_84 ( .A(_249_), .B(_250_), .Y(_251_) );
NOR2X1 NOR2X1_93 ( .A(_246_), .B(_251_), .Y(_15_) );
INVX1 INVX1_75 ( .A(_13_), .Y(_252_) );
NAND2X1 NAND2X1_85 ( .A(1'b0), .B(_15_), .Y(_253_) );
OAI21X1 OAI21X1_76 ( .A(_15_), .B(_252_), .C(_253_), .Y(w_cout_5_) );
INVX1 INVX1_76 ( .A(w_cout_5_), .Y(_257_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_258_) );
NAND2X1 NAND2X1_86 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_259_) );
NAND3X1 NAND3X1_34 ( .A(_257_), .B(_259_), .C(_258_), .Y(_260_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_254_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_255_) );
OAI21X1 OAI21X1_77 ( .A(_254_), .B(_255_), .C(w_cout_5_), .Y(_256_) );
NAND2X1 NAND2X1_87 ( .A(_256_), .B(_260_), .Y(_0__20_) );
OAI21X1 OAI21X1_78 ( .A(_257_), .B(_254_), .C(_259_), .Y(_17__1_) );
INVX1 INVX1_77 ( .A(_17__3_), .Y(_264_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_265_) );
NAND2X1 NAND2X1_88 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_266_) );
NAND3X1 NAND3X1_35 ( .A(_264_), .B(_266_), .C(_265_), .Y(_267_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_261_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_262_) );
OAI21X1 OAI21X1_79 ( .A(_261_), .B(_262_), .C(_17__3_), .Y(_263_) );
NAND2X1 NAND2X1_89 ( .A(_263_), .B(_267_), .Y(_0__23_) );
OAI21X1 OAI21X1_80 ( .A(_264_), .B(_261_), .C(_266_), .Y(_16_) );
INVX1 INVX1_78 ( .A(_17__1_), .Y(_271_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_272_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_273_) );
NAND3X1 NAND3X1_36 ( .A(_271_), .B(_273_), .C(_272_), .Y(_274_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_268_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_269_) );
OAI21X1 OAI21X1_81 ( .A(_268_), .B(_269_), .C(_17__1_), .Y(_270_) );
NAND2X1 NAND2X1_91 ( .A(_270_), .B(_274_), .Y(_0__21_) );
OAI21X1 OAI21X1_82 ( .A(_271_), .B(_268_), .C(_273_), .Y(_17__2_) );
INVX1 INVX1_79 ( .A(_17__2_), .Y(_278_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_279_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_280_) );
NAND3X1 NAND3X1_37 ( .A(_278_), .B(_280_), .C(_279_), .Y(_281_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_275_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_276_) );
OAI21X1 OAI21X1_83 ( .A(_275_), .B(_276_), .C(_17__2_), .Y(_277_) );
NAND2X1 NAND2X1_93 ( .A(_277_), .B(_281_), .Y(_0__22_) );
OAI21X1 OAI21X1_84 ( .A(_278_), .B(_275_), .C(_280_), .Y(_17__3_) );
INVX1 INVX1_80 ( .A(i_add_term1[20]), .Y(_282_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[20]), .B(_282_), .Y(_283_) );
INVX1 INVX1_81 ( .A(i_add_term2[20]), .Y(_284_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term1[20]), .B(_284_), .Y(_285_) );
INVX1 INVX1_82 ( .A(i_add_term1[21]), .Y(_286_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[21]), .B(_286_), .Y(_287_) );
INVX1 INVX1_83 ( .A(i_add_term2[21]), .Y(_288_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term1[21]), .B(_288_), .Y(_289_) );
OAI22X1 OAI22X1_9 ( .A(_283_), .B(_285_), .C(_287_), .D(_289_), .Y(_290_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_291_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_292_) );
NOR2X1 NOR2X1_103 ( .A(_291_), .B(_292_), .Y(_293_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_294_) );
NAND2X1 NAND2X1_94 ( .A(_293_), .B(_294_), .Y(_295_) );
NOR2X1 NOR2X1_104 ( .A(_290_), .B(_295_), .Y(_18_) );
INVX1 INVX1_84 ( .A(_16_), .Y(_296_) );
NAND2X1 NAND2X1_95 ( .A(1'b0), .B(_18_), .Y(_297_) );
OAI21X1 OAI21X1_85 ( .A(_18_), .B(_296_), .C(_297_), .Y(w_cout_6_) );
INVX1 INVX1_85 ( .A(w_cout_6_), .Y(_301_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_302_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_303_) );
NAND3X1 NAND3X1_38 ( .A(_301_), .B(_303_), .C(_302_), .Y(_304_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_298_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_299_) );
OAI21X1 OAI21X1_86 ( .A(_298_), .B(_299_), .C(w_cout_6_), .Y(_300_) );
NAND2X1 NAND2X1_97 ( .A(_300_), .B(_304_), .Y(_0__24_) );
OAI21X1 OAI21X1_87 ( .A(_301_), .B(_298_), .C(_303_), .Y(_20__1_) );
INVX1 INVX1_86 ( .A(_20__3_), .Y(_308_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_309_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_310_) );
NAND3X1 NAND3X1_39 ( .A(_308_), .B(_310_), .C(_309_), .Y(_311_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_305_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_306_) );
OAI21X1 OAI21X1_88 ( .A(_305_), .B(_306_), .C(_20__3_), .Y(_307_) );
NAND2X1 NAND2X1_99 ( .A(_307_), .B(_311_), .Y(_0__27_) );
OAI21X1 OAI21X1_89 ( .A(_308_), .B(_305_), .C(_310_), .Y(_19_) );
INVX1 INVX1_87 ( .A(_20__1_), .Y(_315_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_316_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_317_) );
NAND3X1 NAND3X1_40 ( .A(_315_), .B(_317_), .C(_316_), .Y(_318_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_312_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_313_) );
OAI21X1 OAI21X1_90 ( .A(_312_), .B(_313_), .C(_20__1_), .Y(_314_) );
NAND2X1 NAND2X1_101 ( .A(_314_), .B(_318_), .Y(_0__25_) );
OAI21X1 OAI21X1_91 ( .A(_315_), .B(_312_), .C(_317_), .Y(_20__2_) );
INVX1 INVX1_88 ( .A(_20__2_), .Y(_322_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_323_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_324_) );
NAND3X1 NAND3X1_41 ( .A(_322_), .B(_324_), .C(_323_), .Y(_325_) );
NOR2X1 NOR2X1_108 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_319_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_320_) );
OAI21X1 OAI21X1_92 ( .A(_319_), .B(_320_), .C(_20__2_), .Y(_321_) );
NAND2X1 NAND2X1_103 ( .A(_321_), .B(_325_), .Y(_0__26_) );
OAI21X1 OAI21X1_93 ( .A(_322_), .B(_319_), .C(_324_), .Y(_20__3_) );
INVX1 INVX1_89 ( .A(i_add_term1[24]), .Y(_326_) );
NOR2X1 NOR2X1_109 ( .A(i_add_term2[24]), .B(_326_), .Y(_327_) );
INVX1 INVX1_90 ( .A(i_add_term2[24]), .Y(_328_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term1[24]), .B(_328_), .Y(_329_) );
INVX1 INVX1_91 ( .A(i_add_term1[25]), .Y(_330_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term2[25]), .B(_330_), .Y(_331_) );
INVX1 INVX1_92 ( .A(i_add_term2[25]), .Y(_332_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term1[25]), .B(_332_), .Y(_333_) );
OAI22X1 OAI22X1_10 ( .A(_327_), .B(_329_), .C(_331_), .D(_333_), .Y(_334_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_335_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_336_) );
NOR2X1 NOR2X1_114 ( .A(_335_), .B(_336_), .Y(_337_) );
XOR2X1 XOR2X1_11 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_338_) );
NAND2X1 NAND2X1_104 ( .A(_337_), .B(_338_), .Y(_339_) );
NOR2X1 NOR2X1_115 ( .A(_334_), .B(_339_), .Y(_21_) );
INVX1 INVX1_93 ( .A(_19_), .Y(_340_) );
NAND2X1 NAND2X1_105 ( .A(1'b0), .B(_21_), .Y(_341_) );
OAI21X1 OAI21X1_94 ( .A(_21_), .B(_340_), .C(_341_), .Y(w_cout_7_) );
INVX1 INVX1_94 ( .A(w_cout_7_), .Y(_345_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_346_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_347_) );
NAND3X1 NAND3X1_42 ( .A(_345_), .B(_347_), .C(_346_), .Y(_348_) );
NOR2X1 NOR2X1_116 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_342_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_343_) );
OAI21X1 OAI21X1_95 ( .A(_342_), .B(_343_), .C(w_cout_7_), .Y(_344_) );
NAND2X1 NAND2X1_107 ( .A(_344_), .B(_348_), .Y(_0__28_) );
OAI21X1 OAI21X1_96 ( .A(_345_), .B(_342_), .C(_347_), .Y(_23__1_) );
INVX1 INVX1_95 ( .A(_23__3_), .Y(_352_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_353_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_354_) );
NAND3X1 NAND3X1_43 ( .A(_352_), .B(_354_), .C(_353_), .Y(_355_) );
NOR2X1 NOR2X1_117 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_349_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_350_) );
OAI21X1 OAI21X1_97 ( .A(_349_), .B(_350_), .C(_23__3_), .Y(_351_) );
NAND2X1 NAND2X1_109 ( .A(_351_), .B(_355_), .Y(_0__31_) );
OAI21X1 OAI21X1_98 ( .A(_352_), .B(_349_), .C(_354_), .Y(_22_) );
INVX1 INVX1_96 ( .A(_23__1_), .Y(_359_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_360_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_361_) );
NAND3X1 NAND3X1_44 ( .A(_359_), .B(_361_), .C(_360_), .Y(_362_) );
NOR2X1 NOR2X1_118 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_356_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_357_) );
OAI21X1 OAI21X1_99 ( .A(_356_), .B(_357_), .C(_23__1_), .Y(_358_) );
NAND2X1 NAND2X1_111 ( .A(_358_), .B(_362_), .Y(_0__29_) );
OAI21X1 OAI21X1_100 ( .A(_359_), .B(_356_), .C(_361_), .Y(_23__2_) );
INVX1 INVX1_97 ( .A(_23__2_), .Y(_366_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_367_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_368_) );
NAND3X1 NAND3X1_45 ( .A(_366_), .B(_368_), .C(_367_), .Y(_369_) );
NOR2X1 NOR2X1_119 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_363_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_364_) );
OAI21X1 OAI21X1_101 ( .A(_363_), .B(_364_), .C(_23__2_), .Y(_365_) );
NAND2X1 NAND2X1_113 ( .A(_365_), .B(_369_), .Y(_0__30_) );
OAI21X1 OAI21X1_102 ( .A(_366_), .B(_363_), .C(_368_), .Y(_23__3_) );
INVX1 INVX1_98 ( .A(i_add_term1[28]), .Y(_370_) );
NOR2X1 NOR2X1_120 ( .A(i_add_term2[28]), .B(_370_), .Y(_371_) );
INVX1 INVX1_99 ( .A(i_add_term2[28]), .Y(_372_) );
NOR2X1 NOR2X1_121 ( .A(i_add_term1[28]), .B(_372_), .Y(_373_) );
INVX1 INVX1_100 ( .A(i_add_term1[29]), .Y(_374_) );
NOR2X1 NOR2X1_122 ( .A(i_add_term2[29]), .B(_374_), .Y(_375_) );
INVX1 INVX1_101 ( .A(i_add_term2[29]), .Y(_376_) );
NOR2X1 NOR2X1_123 ( .A(i_add_term1[29]), .B(_376_), .Y(_377_) );
OAI22X1 OAI22X1_11 ( .A(_371_), .B(_373_), .C(_375_), .D(_377_), .Y(_378_) );
NOR2X1 NOR2X1_124 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_379_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_380_) );
BUFX2 BUFX2_47 ( .A(cskip1_inst_rca0_fa0_o_sum), .Y(_0__44_) );
BUFX2 BUFX2_48 ( .A(1'b0), .Y(w_cout_0_) );
BUFX2 BUFX2_49 ( .A(cskip1_inst_cin), .Y(w_cout_11_) );
endmodule
