module CSkipA_22bit ( gnd, vdd, i_add_term1, i_add_term2, sum, cout);

input gnd, vdd;
output cout;
input [21:0] i_add_term1;
input [21:0] i_add_term2;
output [21:0] sum;

BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .Y(cout) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_0__21_), .Y(sum[21]) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .Y(_16_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(_16_), .Y(_17_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .Y(_18_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .B(_18_), .Y(_19_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .Y(_20_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(_20_), .Y(_21_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .Y(_22_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .B(_22_), .Y(_23_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_19_), .C(_21_), .D(_23_), .Y(_24_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_25_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_26_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_26_), .Y(_27_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_28_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_28_), .Y(_29_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_29_), .Y(_3_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_30_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_3_), .Y(_31_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_30_), .C(_31_), .Y(w_cout_1_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[4]), .Y(_32_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(_32_), .Y(_33_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .Y(_34_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[4]), .B(_34_), .Y(_35_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[5]), .Y(_36_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(_36_), .Y(_37_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .Y(_38_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[5]), .B(_38_), .Y(_39_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_35_), .C(_37_), .D(_39_), .Y(_40_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_41_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_42_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_42_), .Y(_43_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_44_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_44_), .Y(_45_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_45_), .Y(_6_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(_46_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_6_), .Y(_47_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_46_), .C(_47_), .Y(w_cout_2_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[8]), .Y(_48_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(_48_), .Y(_49_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .Y(_50_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[8]), .B(_50_), .Y(_51_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[9]), .Y(_52_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(_52_), .Y(_53_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .Y(_54_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[9]), .B(_54_), .Y(_55_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_51_), .C(_53_), .D(_55_), .Y(_56_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_57_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_58_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_58_), .Y(_59_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_60_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_60_), .Y(_61_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_61_), .Y(_9_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_62_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_9_), .Y(_63_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_62_), .C(_63_), .Y(w_cout_3_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[12]), .Y(_64_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(_64_), .Y(_65_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .Y(_66_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[12]), .B(_66_), .Y(_67_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[13]), .Y(_68_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(_68_), .Y(_69_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .Y(_70_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[13]), .B(_70_), .Y(_71_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_67_), .C(_69_), .D(_71_), .Y(_72_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_73_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_74_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_74_), .Y(_75_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_76_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_76_), .Y(_77_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_77_), .Y(_12_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(_78_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_12_), .Y(_79_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_78_), .C(_79_), .Y(w_cout_4_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[16]), .Y(_80_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(_80_), .Y(_81_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .Y(_82_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[16]), .B(_82_), .Y(_83_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[17]), .Y(_84_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(_84_), .Y(_85_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .Y(_86_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[17]), .B(_86_), .Y(_87_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_83_), .C(_85_), .D(_87_), .Y(_88_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_89_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_90_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_90_), .Y(_91_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_92_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_92_), .Y(_93_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_93_), .Y(_15_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_94_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_15_), .Y(_95_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_94_), .C(_95_), .Y(cskip2_inst_cin) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_99_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_100_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_101_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_101_), .C(_100_), .Y(_102_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_96_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_97_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_97_), .C(gnd), .Y(_98_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_102_), .Y(_0__0_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_96_), .C(_101_), .Y(_2__1_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_2__1_), .Y(_106_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_107_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_108_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_106_), .B(_108_), .C(_107_), .Y(_109_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_103_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_104_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_104_), .C(_2__1_), .Y(_105_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_109_), .Y(_0__1_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_106_), .B(_103_), .C(_108_), .Y(_2__2_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_2__2_), .Y(_113_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_114_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_115_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_115_), .C(_114_), .Y(_116_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_110_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_111_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_111_), .C(_2__2_), .Y(_112_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_116_), .Y(_0__2_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_110_), .C(_115_), .Y(_2__3_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_2__3_), .Y(_120_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_121_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_122_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_122_), .C(_121_), .Y(_123_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_117_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_118_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_118_), .C(_2__3_), .Y(_119_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_123_), .Y(_0__3_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_117_), .C(_122_), .Y(_1_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .Y(_127_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_128_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_129_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_129_), .C(_128_), .Y(_130_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_124_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_125_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_125_), .C(w_cout_1_), .Y(_126_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_130_), .Y(_0__4_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_124_), .C(_129_), .Y(_5__1_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_5__1_), .Y(_134_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_135_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_136_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_136_), .C(_135_), .Y(_137_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_131_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_132_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_132_), .C(_5__1_), .Y(_133_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_137_), .Y(_0__5_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_131_), .C(_136_), .Y(_5__2_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_5__2_), .Y(_141_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_142_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_143_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_143_), .C(_142_), .Y(_144_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_138_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_139_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_139_), .C(_5__2_), .Y(_140_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_144_), .Y(_0__6_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_138_), .C(_143_), .Y(_5__3_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_5__3_), .Y(_148_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_149_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_150_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_150_), .C(_149_), .Y(_151_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_145_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_146_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_146_), .C(_5__3_), .Y(_147_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_151_), .Y(_0__7_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_145_), .C(_150_), .Y(_4_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .Y(_155_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_156_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_157_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_157_), .C(_156_), .Y(_158_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_152_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_153_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_153_), .C(w_cout_2_), .Y(_154_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_158_), .Y(_0__8_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_152_), .C(_157_), .Y(_8__1_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_8__1_), .Y(_162_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_163_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_164_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_164_), .C(_163_), .Y(_165_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_159_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_160_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_159_), .B(_160_), .C(_8__1_), .Y(_161_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_165_), .Y(_0__9_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_159_), .C(_164_), .Y(_8__2_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_8__2_), .Y(_169_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_170_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_171_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_171_), .C(_170_), .Y(_172_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_166_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_167_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_167_), .C(_8__2_), .Y(_168_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_172_), .Y(_0__10_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_166_), .C(_171_), .Y(_8__3_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_8__3_), .Y(_176_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_177_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_178_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_178_), .C(_177_), .Y(_179_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_173_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_174_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(_174_), .C(_8__3_), .Y(_175_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_175_), .B(_179_), .Y(_0__11_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_173_), .C(_178_), .Y(_7_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .Y(_183_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_184_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_185_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_185_), .C(_184_), .Y(_186_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_180_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_181_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_181_), .C(w_cout_3_), .Y(_182_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_186_), .Y(_0__12_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_180_), .C(_185_), .Y(_11__1_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_11__1_), .Y(_190_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_191_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_192_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_192_), .C(_191_), .Y(_193_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_187_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_188_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(_188_), .C(_11__1_), .Y(_189_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_193_), .Y(_0__13_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_187_), .C(_192_), .Y(_11__2_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_11__2_), .Y(_197_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_198_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_199_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_199_), .C(_198_), .Y(_200_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_194_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_195_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_195_), .C(_11__2_), .Y(_196_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_200_), .Y(_0__14_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_194_), .C(_199_), .Y(_11__3_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_11__3_), .Y(_204_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_205_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_206_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_206_), .C(_205_), .Y(_207_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_201_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_202_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_202_), .C(_11__3_), .Y(_203_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_207_), .Y(_0__15_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_201_), .C(_206_), .Y(_10_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .Y(_211_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_212_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_213_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_213_), .C(_212_), .Y(_214_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_208_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_209_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_209_), .C(w_cout_4_), .Y(_210_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_210_), .B(_214_), .Y(_0__16_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_208_), .C(_213_), .Y(_14__1_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_14__1_), .Y(_218_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_219_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_220_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(_220_), .C(_219_), .Y(_221_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_215_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_216_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_216_), .C(_14__1_), .Y(_217_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_221_), .Y(_0__17_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(_215_), .C(_220_), .Y(_14__2_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_14__2_), .Y(_225_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_226_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_227_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_227_), .C(_226_), .Y(_228_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_222_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_223_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_223_), .C(_14__2_), .Y(_224_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_228_), .Y(_0__18_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_222_), .C(_227_), .Y(_14__3_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_14__3_), .Y(_232_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_233_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_234_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_234_), .C(_233_), .Y(_235_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_229_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_230_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_230_), .C(_14__3_), .Y(_231_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_235_), .Y(_0__19_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_229_), .C(_234_), .Y(_13_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_cin), .Y(_239_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_240_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_241_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_241_), .C(_240_), .Y(_242_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_236_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_237_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_237_), .C(cskip2_inst_cin), .Y(_238_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_238_), .B(_242_), .Y(_0__20_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_236_), .C(_241_), .Y(cskip2_inst_rca0_w_CARRY_1_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_rca0_w_CARRY_1_), .Y(_246_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_247_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_248_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_248_), .C(_247_), .Y(_249_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_243_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_244_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_244_), .C(cskip2_inst_rca0_w_CARRY_1_), .Y(_245_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_249_), .Y(_0__21_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_243_), .C(_248_), .Y(cskip2_inst_rca0_w_CARRY_2_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_rca0_w_CARRY_2_), .Y(_251_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_252_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_250_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_250_), .C(_252_), .Y(cskip2_inst_rca0_w_CARRY_3_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_rca0_w_CARRY_3_), .Y(_254_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_255_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_253_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_253_), .C(_255_), .Y(cskip2_inst_cout0) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[21]), .Y(_260_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(_260_), .Y(_261_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .Y(_262_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[21]), .B(_262_), .Y(_263_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[20]), .Y(_256_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(_256_), .Y(_257_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .Y(_258_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[20]), .B(_258_), .Y(_259_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_263_), .C(_257_), .D(_259_), .Y(cskip2_inst_skip0_P) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_cout0), .Y(_264_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(cskip2_inst_skip0_P), .Y(_265_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_skip0_P), .B(_264_), .C(_265_), .Y(w_cout_6_) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_2__0_) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .Y(_5__0_) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(_5__4_) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .Y(_8__0_) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .Y(_11__0_) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(_11__4_) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .Y(_14__0_) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_cin), .Y(cskip2_inst_rca0_w_CARRY_0_) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_cout0), .Y(cskip2_inst_rca0_w_CARRY_4_) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(cskip2_inst_cin), .Y(w_cout_5_) );
endmodule
