module cla_49bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add1[19], i_add1[20], i_add1[21], i_add1[22], i_add1[23], i_add1[24], i_add1[25], i_add1[26], i_add1[27], i_add1[28], i_add1[29], i_add1[30], i_add1[31], i_add1[32], i_add1[33], i_add1[34], i_add1[35], i_add1[36], i_add1[37], i_add1[38], i_add1[39], i_add1[40], i_add1[41], i_add1[42], i_add1[43], i_add1[44], i_add1[45], i_add1[46], i_add1[47], i_add1[48], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], i_add2[19], i_add2[20], i_add2[21], i_add2[22], i_add2[23], i_add2[24], i_add2[25], i_add2[26], i_add2[27], i_add2[28], i_add2[29], i_add2[30], i_add2[31], i_add2[32], i_add2[33], i_add2[34], i_add2[35], i_add2[36], i_add2[37], i_add2[38], i_add2[39], i_add2[40], i_add2[41], i_add2[42], i_add2[43], i_add2[44], i_add2[45], i_add2[46], i_add2[47], i_add2[48], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21], o_result[22], o_result[23], o_result[24], o_result[25], o_result[26], o_result[27], o_result[28], o_result[29], o_result[30], o_result[31], o_result[32], o_result[33], o_result[34], o_result[35], o_result[36], o_result[37], o_result[38], o_result[39], o_result[40], o_result[41], o_result[42], o_result[43], o_result[44], o_result[45], o_result[46], o_result[47], o_result[48], o_result[49]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add1[19];
input i_add1[20];
input i_add1[21];
input i_add1[22];
input i_add1[23];
input i_add1[24];
input i_add1[25];
input i_add1[26];
input i_add1[27];
input i_add1[28];
input i_add1[29];
input i_add1[30];
input i_add1[31];
input i_add1[32];
input i_add1[33];
input i_add1[34];
input i_add1[35];
input i_add1[36];
input i_add1[37];
input i_add1[38];
input i_add1[39];
input i_add1[40];
input i_add1[41];
input i_add1[42];
input i_add1[43];
input i_add1[44];
input i_add1[45];
input i_add1[46];
input i_add1[47];
input i_add1[48];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
input i_add2[19];
input i_add2[20];
input i_add2[21];
input i_add2[22];
input i_add2[23];
input i_add2[24];
input i_add2[25];
input i_add2[26];
input i_add2[27];
input i_add2[28];
input i_add2[29];
input i_add2[30];
input i_add2[31];
input i_add2[32];
input i_add2[33];
input i_add2[34];
input i_add2[35];
input i_add2[36];
input i_add2[37];
input i_add2[38];
input i_add2[39];
input i_add2[40];
input i_add2[41];
input i_add2[42];
input i_add2[43];
input i_add2[44];
input i_add2[45];
input i_add2[46];
input i_add2[47];
input i_add2[48];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];
output o_result[22];
output o_result[23];
output o_result[24];
output o_result[25];
output o_result[26];
output o_result[27];
output o_result[28];
output o_result[29];
output o_result[30];
output o_result[31];
output o_result[32];
output o_result[33];
output o_result[34];
output o_result[35];
output o_result[36];
output o_result[37];
output o_result[38];
output o_result[39];
output o_result[40];
output o_result[41];
output o_result[42];
output o_result[43];
output o_result[44];
output o_result[45];
output o_result[46];
output o_result[47];
output o_result[48];
output o_result[49];

NAND3X1 NAND3X1_1 ( .A(_281_), .B(_283_), .C(_282_), .Y(_284_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_278_) );
AND2X2 AND2X2_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_279_) );
OAI21X1 OAI21X1_1 ( .A(_278_), .B(_279_), .C(w_C_4_), .Y(_280_) );
NAND2X1 NAND2X1_1 ( .A(_280_), .B(_284_), .Y(_277__4_) );
INVX1 INVX1_1 ( .A(w_C_5_), .Y(_288_) );
OR2X2 OR2X2_1 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_289_) );
NAND2X1 NAND2X1_2 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_290_) );
NAND3X1 NAND3X1_2 ( .A(_288_), .B(_290_), .C(_289_), .Y(_291_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_285_) );
AND2X2 AND2X2_2 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_286_) );
OAI21X1 OAI21X1_2 ( .A(_285_), .B(_286_), .C(w_C_5_), .Y(_287_) );
NAND2X1 NAND2X1_3 ( .A(_287_), .B(_291_), .Y(_277__5_) );
INVX1 INVX1_2 ( .A(w_C_6_), .Y(_295_) );
OR2X2 OR2X2_2 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_296_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_297_) );
NAND3X1 NAND3X1_3 ( .A(_295_), .B(_297_), .C(_296_), .Y(_298_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_292_) );
AND2X2 AND2X2_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_293_) );
OAI21X1 OAI21X1_3 ( .A(_292_), .B(_293_), .C(w_C_6_), .Y(_294_) );
NAND2X1 NAND2X1_5 ( .A(_294_), .B(_298_), .Y(_277__6_) );
INVX1 INVX1_3 ( .A(w_C_7_), .Y(_302_) );
OR2X2 OR2X2_3 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_303_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_304_) );
NAND3X1 NAND3X1_4 ( .A(_302_), .B(_304_), .C(_303_), .Y(_305_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_299_) );
AND2X2 AND2X2_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_300_) );
OAI21X1 OAI21X1_4 ( .A(_299_), .B(_300_), .C(w_C_7_), .Y(_301_) );
NAND2X1 NAND2X1_7 ( .A(_301_), .B(_305_), .Y(_277__7_) );
INVX1 INVX1_4 ( .A(w_C_8_), .Y(_309_) );
OR2X2 OR2X2_4 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_310_) );
NAND2X1 NAND2X1_8 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_311_) );
NAND3X1 NAND3X1_5 ( .A(_309_), .B(_311_), .C(_310_), .Y(_312_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_306_) );
AND2X2 AND2X2_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_307_) );
OAI21X1 OAI21X1_5 ( .A(_306_), .B(_307_), .C(w_C_8_), .Y(_308_) );
NAND2X1 NAND2X1_9 ( .A(_308_), .B(_312_), .Y(_277__8_) );
INVX1 INVX1_5 ( .A(w_C_9_), .Y(_316_) );
OR2X2 OR2X2_5 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_317_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_318_) );
NAND3X1 NAND3X1_6 ( .A(_316_), .B(_318_), .C(_317_), .Y(_319_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_313_) );
AND2X2 AND2X2_6 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_314_) );
OAI21X1 OAI21X1_6 ( .A(_313_), .B(_314_), .C(w_C_9_), .Y(_315_) );
NAND2X1 NAND2X1_11 ( .A(_315_), .B(_319_), .Y(_277__9_) );
INVX1 INVX1_6 ( .A(w_C_10_), .Y(_323_) );
OR2X2 OR2X2_6 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_324_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_325_) );
NAND3X1 NAND3X1_7 ( .A(_323_), .B(_325_), .C(_324_), .Y(_326_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_320_) );
AND2X2 AND2X2_7 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_321_) );
OAI21X1 OAI21X1_7 ( .A(_320_), .B(_321_), .C(w_C_10_), .Y(_322_) );
NAND2X1 NAND2X1_13 ( .A(_322_), .B(_326_), .Y(_277__10_) );
INVX1 INVX1_7 ( .A(w_C_11_), .Y(_330_) );
OR2X2 OR2X2_7 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_331_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_332_) );
NAND3X1 NAND3X1_8 ( .A(_330_), .B(_332_), .C(_331_), .Y(_333_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_327_) );
AND2X2 AND2X2_8 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_328_) );
OAI21X1 OAI21X1_8 ( .A(_327_), .B(_328_), .C(w_C_11_), .Y(_329_) );
NAND2X1 NAND2X1_15 ( .A(_329_), .B(_333_), .Y(_277__11_) );
INVX1 INVX1_8 ( .A(w_C_12_), .Y(_337_) );
OR2X2 OR2X2_8 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_338_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_339_) );
NAND3X1 NAND3X1_9 ( .A(_337_), .B(_339_), .C(_338_), .Y(_340_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_334_) );
AND2X2 AND2X2_9 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_335_) );
OAI21X1 OAI21X1_9 ( .A(_334_), .B(_335_), .C(w_C_12_), .Y(_336_) );
NAND2X1 NAND2X1_17 ( .A(_336_), .B(_340_), .Y(_277__12_) );
INVX1 INVX1_9 ( .A(w_C_13_), .Y(_344_) );
OR2X2 OR2X2_9 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_345_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_346_) );
NAND3X1 NAND3X1_10 ( .A(_344_), .B(_346_), .C(_345_), .Y(_347_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_341_) );
AND2X2 AND2X2_10 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_342_) );
OAI21X1 OAI21X1_10 ( .A(_341_), .B(_342_), .C(w_C_13_), .Y(_343_) );
NAND2X1 NAND2X1_19 ( .A(_343_), .B(_347_), .Y(_277__13_) );
INVX1 INVX1_10 ( .A(w_C_14_), .Y(_351_) );
OR2X2 OR2X2_10 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_352_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_353_) );
NAND3X1 NAND3X1_11 ( .A(_351_), .B(_353_), .C(_352_), .Y(_354_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_348_) );
AND2X2 AND2X2_11 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_349_) );
OAI21X1 OAI21X1_11 ( .A(_348_), .B(_349_), .C(w_C_14_), .Y(_350_) );
NAND2X1 NAND2X1_21 ( .A(_350_), .B(_354_), .Y(_277__14_) );
INVX1 INVX1_11 ( .A(w_C_15_), .Y(_358_) );
OR2X2 OR2X2_11 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_359_) );
NAND2X1 NAND2X1_22 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_360_) );
NAND3X1 NAND3X1_12 ( .A(_358_), .B(_360_), .C(_359_), .Y(_361_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_355_) );
AND2X2 AND2X2_12 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_356_) );
OAI21X1 OAI21X1_12 ( .A(_355_), .B(_356_), .C(w_C_15_), .Y(_357_) );
NAND2X1 NAND2X1_23 ( .A(_357_), .B(_361_), .Y(_277__15_) );
INVX1 INVX1_12 ( .A(w_C_16_), .Y(_365_) );
OR2X2 OR2X2_12 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_366_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_367_) );
NAND3X1 NAND3X1_13 ( .A(_365_), .B(_367_), .C(_366_), .Y(_368_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_362_) );
AND2X2 AND2X2_13 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_363_) );
OAI21X1 OAI21X1_13 ( .A(_362_), .B(_363_), .C(w_C_16_), .Y(_364_) );
NAND2X1 NAND2X1_25 ( .A(_364_), .B(_368_), .Y(_277__16_) );
INVX1 INVX1_13 ( .A(w_C_17_), .Y(_372_) );
OR2X2 OR2X2_13 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_373_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_374_) );
NAND3X1 NAND3X1_14 ( .A(_372_), .B(_374_), .C(_373_), .Y(_375_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_369_) );
AND2X2 AND2X2_14 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_370_) );
OAI21X1 OAI21X1_14 ( .A(_369_), .B(_370_), .C(w_C_17_), .Y(_371_) );
NAND2X1 NAND2X1_27 ( .A(_371_), .B(_375_), .Y(_277__17_) );
INVX1 INVX1_14 ( .A(w_C_18_), .Y(_379_) );
OR2X2 OR2X2_14 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_380_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_381_) );
NAND3X1 NAND3X1_15 ( .A(_379_), .B(_381_), .C(_380_), .Y(_382_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_376_) );
AND2X2 AND2X2_15 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_377_) );
OAI21X1 OAI21X1_15 ( .A(_376_), .B(_377_), .C(w_C_18_), .Y(_378_) );
NAND2X1 NAND2X1_29 ( .A(_378_), .B(_382_), .Y(_277__18_) );
INVX1 INVX1_15 ( .A(w_C_19_), .Y(_386_) );
OR2X2 OR2X2_15 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_387_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_388_) );
NAND3X1 NAND3X1_16 ( .A(_386_), .B(_388_), .C(_387_), .Y(_389_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_383_) );
AND2X2 AND2X2_16 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_384_) );
OAI21X1 OAI21X1_16 ( .A(_383_), .B(_384_), .C(w_C_19_), .Y(_385_) );
NAND2X1 NAND2X1_31 ( .A(_385_), .B(_389_), .Y(_277__19_) );
INVX1 INVX1_16 ( .A(w_C_20_), .Y(_393_) );
OR2X2 OR2X2_16 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_394_) );
NAND2X1 NAND2X1_32 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_395_) );
NAND3X1 NAND3X1_17 ( .A(_393_), .B(_395_), .C(_394_), .Y(_396_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_390_) );
AND2X2 AND2X2_17 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_391_) );
OAI21X1 OAI21X1_17 ( .A(_390_), .B(_391_), .C(w_C_20_), .Y(_392_) );
NAND2X1 NAND2X1_33 ( .A(_392_), .B(_396_), .Y(_277__20_) );
INVX1 INVX1_17 ( .A(w_C_21_), .Y(_400_) );
OR2X2 OR2X2_17 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_401_) );
NAND2X1 NAND2X1_34 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_402_) );
NAND3X1 NAND3X1_18 ( .A(_400_), .B(_402_), .C(_401_), .Y(_403_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_397_) );
AND2X2 AND2X2_18 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_398_) );
OAI21X1 OAI21X1_18 ( .A(_397_), .B(_398_), .C(w_C_21_), .Y(_399_) );
NAND2X1 NAND2X1_35 ( .A(_399_), .B(_403_), .Y(_277__21_) );
INVX1 INVX1_18 ( .A(w_C_22_), .Y(_407_) );
OR2X2 OR2X2_18 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_408_) );
NAND2X1 NAND2X1_36 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_409_) );
NAND3X1 NAND3X1_19 ( .A(_407_), .B(_409_), .C(_408_), .Y(_410_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_404_) );
AND2X2 AND2X2_19 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_405_) );
OAI21X1 OAI21X1_19 ( .A(_404_), .B(_405_), .C(w_C_22_), .Y(_406_) );
NAND2X1 NAND2X1_37 ( .A(_406_), .B(_410_), .Y(_277__22_) );
INVX1 INVX1_19 ( .A(w_C_23_), .Y(_414_) );
OR2X2 OR2X2_19 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_415_) );
NAND2X1 NAND2X1_38 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_416_) );
NAND3X1 NAND3X1_20 ( .A(_414_), .B(_416_), .C(_415_), .Y(_417_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_411_) );
AND2X2 AND2X2_20 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_412_) );
OAI21X1 OAI21X1_20 ( .A(_411_), .B(_412_), .C(w_C_23_), .Y(_413_) );
NAND2X1 NAND2X1_39 ( .A(_413_), .B(_417_), .Y(_277__23_) );
INVX1 INVX1_20 ( .A(w_C_24_), .Y(_421_) );
OR2X2 OR2X2_20 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_422_) );
NAND2X1 NAND2X1_40 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_423_) );
NAND3X1 NAND3X1_21 ( .A(_421_), .B(_423_), .C(_422_), .Y(_424_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_418_) );
AND2X2 AND2X2_21 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_419_) );
OAI21X1 OAI21X1_21 ( .A(_418_), .B(_419_), .C(w_C_24_), .Y(_420_) );
NAND2X1 NAND2X1_41 ( .A(_420_), .B(_424_), .Y(_277__24_) );
INVX1 INVX1_21 ( .A(w_C_25_), .Y(_428_) );
OR2X2 OR2X2_21 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_429_) );
NAND2X1 NAND2X1_42 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_430_) );
NAND3X1 NAND3X1_22 ( .A(_428_), .B(_430_), .C(_429_), .Y(_431_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_425_) );
AND2X2 AND2X2_22 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_426_) );
OAI21X1 OAI21X1_22 ( .A(_425_), .B(_426_), .C(w_C_25_), .Y(_427_) );
NAND2X1 NAND2X1_43 ( .A(_427_), .B(_431_), .Y(_277__25_) );
INVX1 INVX1_22 ( .A(w_C_26_), .Y(_435_) );
OR2X2 OR2X2_22 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_436_) );
NAND2X1 NAND2X1_44 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_437_) );
NAND3X1 NAND3X1_23 ( .A(_435_), .B(_437_), .C(_436_), .Y(_438_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_432_) );
AND2X2 AND2X2_23 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_433_) );
OAI21X1 OAI21X1_23 ( .A(_432_), .B(_433_), .C(w_C_26_), .Y(_434_) );
NAND2X1 NAND2X1_45 ( .A(_434_), .B(_438_), .Y(_277__26_) );
INVX1 INVX1_23 ( .A(w_C_27_), .Y(_442_) );
OR2X2 OR2X2_23 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_443_) );
NAND2X1 NAND2X1_46 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_444_) );
NAND3X1 NAND3X1_24 ( .A(_442_), .B(_444_), .C(_443_), .Y(_445_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_439_) );
AND2X2 AND2X2_24 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_440_) );
OAI21X1 OAI21X1_24 ( .A(_439_), .B(_440_), .C(w_C_27_), .Y(_441_) );
NAND2X1 NAND2X1_47 ( .A(_441_), .B(_445_), .Y(_277__27_) );
INVX1 INVX1_24 ( .A(w_C_28_), .Y(_449_) );
OR2X2 OR2X2_24 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_450_) );
NAND2X1 NAND2X1_48 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_451_) );
NAND3X1 NAND3X1_25 ( .A(_449_), .B(_451_), .C(_450_), .Y(_452_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_446_) );
AND2X2 AND2X2_25 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_447_) );
OAI21X1 OAI21X1_25 ( .A(_446_), .B(_447_), .C(w_C_28_), .Y(_448_) );
NAND2X1 NAND2X1_49 ( .A(_448_), .B(_452_), .Y(_277__28_) );
INVX1 INVX1_25 ( .A(w_C_29_), .Y(_456_) );
OR2X2 OR2X2_25 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_457_) );
NAND2X1 NAND2X1_50 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_458_) );
NAND3X1 NAND3X1_26 ( .A(_456_), .B(_458_), .C(_457_), .Y(_459_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_453_) );
AND2X2 AND2X2_26 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_454_) );
OAI21X1 OAI21X1_26 ( .A(_453_), .B(_454_), .C(w_C_29_), .Y(_455_) );
NAND2X1 NAND2X1_51 ( .A(_455_), .B(_459_), .Y(_277__29_) );
INVX1 INVX1_26 ( .A(w_C_30_), .Y(_463_) );
OR2X2 OR2X2_26 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_464_) );
NAND2X1 NAND2X1_52 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_465_) );
NAND3X1 NAND3X1_27 ( .A(_463_), .B(_465_), .C(_464_), .Y(_466_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_460_) );
AND2X2 AND2X2_27 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_461_) );
OAI21X1 OAI21X1_27 ( .A(_460_), .B(_461_), .C(w_C_30_), .Y(_462_) );
NAND2X1 NAND2X1_53 ( .A(_462_), .B(_466_), .Y(_277__30_) );
INVX1 INVX1_27 ( .A(w_C_31_), .Y(_470_) );
OR2X2 OR2X2_27 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_471_) );
NAND2X1 NAND2X1_54 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_472_) );
NAND3X1 NAND3X1_28 ( .A(_470_), .B(_472_), .C(_471_), .Y(_473_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_467_) );
AND2X2 AND2X2_28 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_468_) );
OAI21X1 OAI21X1_28 ( .A(_467_), .B(_468_), .C(w_C_31_), .Y(_469_) );
NAND2X1 NAND2X1_55 ( .A(_469_), .B(_473_), .Y(_277__31_) );
INVX1 INVX1_28 ( .A(w_C_32_), .Y(_477_) );
OR2X2 OR2X2_28 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_478_) );
NAND2X1 NAND2X1_56 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_479_) );
NAND3X1 NAND3X1_29 ( .A(_477_), .B(_479_), .C(_478_), .Y(_480_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_474_) );
AND2X2 AND2X2_29 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_475_) );
OAI21X1 OAI21X1_29 ( .A(_474_), .B(_475_), .C(w_C_32_), .Y(_476_) );
NAND2X1 NAND2X1_57 ( .A(_476_), .B(_480_), .Y(_277__32_) );
INVX1 INVX1_29 ( .A(w_C_33_), .Y(_484_) );
OR2X2 OR2X2_29 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_485_) );
NAND2X1 NAND2X1_58 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_486_) );
NAND3X1 NAND3X1_30 ( .A(_484_), .B(_486_), .C(_485_), .Y(_487_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_481_) );
AND2X2 AND2X2_30 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_482_) );
OAI21X1 OAI21X1_30 ( .A(_481_), .B(_482_), .C(w_C_33_), .Y(_483_) );
NAND2X1 NAND2X1_59 ( .A(_483_), .B(_487_), .Y(_277__33_) );
INVX1 INVX1_30 ( .A(w_C_34_), .Y(_491_) );
OR2X2 OR2X2_30 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_492_) );
NAND2X1 NAND2X1_60 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_493_) );
NAND3X1 NAND3X1_31 ( .A(_491_), .B(_493_), .C(_492_), .Y(_494_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_488_) );
AND2X2 AND2X2_31 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_489_) );
OAI21X1 OAI21X1_31 ( .A(_488_), .B(_489_), .C(w_C_34_), .Y(_490_) );
NAND2X1 NAND2X1_61 ( .A(_490_), .B(_494_), .Y(_277__34_) );
INVX1 INVX1_31 ( .A(w_C_35_), .Y(_498_) );
OR2X2 OR2X2_31 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_499_) );
NAND2X1 NAND2X1_62 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_500_) );
NAND3X1 NAND3X1_32 ( .A(_498_), .B(_500_), .C(_499_), .Y(_501_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_495_) );
AND2X2 AND2X2_32 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_496_) );
OAI21X1 OAI21X1_32 ( .A(_495_), .B(_496_), .C(w_C_35_), .Y(_497_) );
NAND2X1 NAND2X1_63 ( .A(_497_), .B(_501_), .Y(_277__35_) );
INVX1 INVX1_32 ( .A(w_C_36_), .Y(_505_) );
OR2X2 OR2X2_32 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_506_) );
NAND2X1 NAND2X1_64 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_507_) );
NAND3X1 NAND3X1_33 ( .A(_505_), .B(_507_), .C(_506_), .Y(_508_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_502_) );
AND2X2 AND2X2_33 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_503_) );
OAI21X1 OAI21X1_33 ( .A(_502_), .B(_503_), .C(w_C_36_), .Y(_504_) );
NAND2X1 NAND2X1_65 ( .A(_504_), .B(_508_), .Y(_277__36_) );
INVX1 INVX1_33 ( .A(w_C_37_), .Y(_512_) );
OR2X2 OR2X2_33 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_513_) );
NAND2X1 NAND2X1_66 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_514_) );
NAND3X1 NAND3X1_34 ( .A(_512_), .B(_514_), .C(_513_), .Y(_515_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_509_) );
AND2X2 AND2X2_34 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_510_) );
OAI21X1 OAI21X1_34 ( .A(_509_), .B(_510_), .C(w_C_37_), .Y(_511_) );
NAND2X1 NAND2X1_67 ( .A(_511_), .B(_515_), .Y(_277__37_) );
INVX1 INVX1_34 ( .A(w_C_38_), .Y(_519_) );
OR2X2 OR2X2_34 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_520_) );
NAND2X1 NAND2X1_68 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_521_) );
NAND3X1 NAND3X1_35 ( .A(_519_), .B(_521_), .C(_520_), .Y(_522_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_516_) );
AND2X2 AND2X2_35 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_517_) );
OAI21X1 OAI21X1_35 ( .A(_516_), .B(_517_), .C(w_C_38_), .Y(_518_) );
NAND2X1 NAND2X1_69 ( .A(_518_), .B(_522_), .Y(_277__38_) );
INVX1 INVX1_35 ( .A(w_C_39_), .Y(_526_) );
OR2X2 OR2X2_35 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_527_) );
NAND2X1 NAND2X1_70 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_528_) );
NAND3X1 NAND3X1_36 ( .A(_526_), .B(_528_), .C(_527_), .Y(_529_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_523_) );
AND2X2 AND2X2_36 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_524_) );
OAI21X1 OAI21X1_36 ( .A(_523_), .B(_524_), .C(w_C_39_), .Y(_525_) );
NAND2X1 NAND2X1_71 ( .A(_525_), .B(_529_), .Y(_277__39_) );
INVX1 INVX1_36 ( .A(w_C_40_), .Y(_533_) );
OR2X2 OR2X2_36 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_534_) );
NAND2X1 NAND2X1_72 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_535_) );
NAND3X1 NAND3X1_37 ( .A(_533_), .B(_535_), .C(_534_), .Y(_536_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_530_) );
AND2X2 AND2X2_37 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_531_) );
OAI21X1 OAI21X1_37 ( .A(_530_), .B(_531_), .C(w_C_40_), .Y(_532_) );
NAND2X1 NAND2X1_73 ( .A(_532_), .B(_536_), .Y(_277__40_) );
INVX1 INVX1_37 ( .A(w_C_41_), .Y(_540_) );
OR2X2 OR2X2_37 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_541_) );
NAND2X1 NAND2X1_74 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_542_) );
NAND3X1 NAND3X1_38 ( .A(_540_), .B(_542_), .C(_541_), .Y(_543_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_537_) );
AND2X2 AND2X2_38 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_538_) );
OAI21X1 OAI21X1_38 ( .A(_537_), .B(_538_), .C(w_C_41_), .Y(_539_) );
NAND2X1 NAND2X1_75 ( .A(_539_), .B(_543_), .Y(_277__41_) );
INVX1 INVX1_38 ( .A(w_C_42_), .Y(_547_) );
OR2X2 OR2X2_38 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_548_) );
NAND2X1 NAND2X1_76 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_549_) );
NAND3X1 NAND3X1_39 ( .A(_547_), .B(_549_), .C(_548_), .Y(_550_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_544_) );
AND2X2 AND2X2_39 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_545_) );
OAI21X1 OAI21X1_39 ( .A(_544_), .B(_545_), .C(w_C_42_), .Y(_546_) );
NAND2X1 NAND2X1_77 ( .A(_546_), .B(_550_), .Y(_277__42_) );
INVX1 INVX1_39 ( .A(w_C_43_), .Y(_554_) );
OR2X2 OR2X2_39 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_555_) );
NAND2X1 NAND2X1_78 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_556_) );
NAND3X1 NAND3X1_40 ( .A(_554_), .B(_556_), .C(_555_), .Y(_557_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_551_) );
AND2X2 AND2X2_40 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_552_) );
OAI21X1 OAI21X1_40 ( .A(_551_), .B(_552_), .C(w_C_43_), .Y(_553_) );
NAND2X1 NAND2X1_79 ( .A(_553_), .B(_557_), .Y(_277__43_) );
INVX1 INVX1_40 ( .A(w_C_44_), .Y(_561_) );
OR2X2 OR2X2_40 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_562_) );
NAND2X1 NAND2X1_80 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_563_) );
NAND3X1 NAND3X1_41 ( .A(_561_), .B(_563_), .C(_562_), .Y(_564_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_558_) );
AND2X2 AND2X2_41 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_559_) );
OAI21X1 OAI21X1_41 ( .A(_558_), .B(_559_), .C(w_C_44_), .Y(_560_) );
NAND2X1 NAND2X1_81 ( .A(_560_), .B(_564_), .Y(_277__44_) );
INVX1 INVX1_41 ( .A(w_C_45_), .Y(_568_) );
OR2X2 OR2X2_41 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_569_) );
NAND2X1 NAND2X1_82 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_570_) );
NAND3X1 NAND3X1_42 ( .A(_568_), .B(_570_), .C(_569_), .Y(_571_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_565_) );
AND2X2 AND2X2_42 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_566_) );
OAI21X1 OAI21X1_42 ( .A(_565_), .B(_566_), .C(w_C_45_), .Y(_567_) );
NAND2X1 NAND2X1_83 ( .A(_567_), .B(_571_), .Y(_277__45_) );
INVX1 INVX1_42 ( .A(w_C_46_), .Y(_575_) );
OR2X2 OR2X2_42 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_576_) );
NAND2X1 NAND2X1_84 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_577_) );
NAND3X1 NAND3X1_43 ( .A(_575_), .B(_577_), .C(_576_), .Y(_578_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_572_) );
AND2X2 AND2X2_43 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_573_) );
OAI21X1 OAI21X1_43 ( .A(_572_), .B(_573_), .C(w_C_46_), .Y(_574_) );
NAND2X1 NAND2X1_85 ( .A(_574_), .B(_578_), .Y(_277__46_) );
INVX1 INVX1_43 ( .A(w_C_47_), .Y(_582_) );
OR2X2 OR2X2_43 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_583_) );
NAND2X1 NAND2X1_86 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_584_) );
NAND3X1 NAND3X1_44 ( .A(_582_), .B(_584_), .C(_583_), .Y(_585_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_579_) );
AND2X2 AND2X2_44 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_580_) );
OAI21X1 OAI21X1_44 ( .A(_579_), .B(_580_), .C(w_C_47_), .Y(_581_) );
NAND2X1 NAND2X1_87 ( .A(_581_), .B(_585_), .Y(_277__47_) );
INVX1 INVX1_44 ( .A(w_C_48_), .Y(_589_) );
OR2X2 OR2X2_44 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_590_) );
NAND2X1 NAND2X1_88 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_591_) );
NAND3X1 NAND3X1_45 ( .A(_589_), .B(_591_), .C(_590_), .Y(_592_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_586_) );
AND2X2 AND2X2_45 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_587_) );
OAI21X1 OAI21X1_45 ( .A(_586_), .B(_587_), .C(w_C_48_), .Y(_588_) );
NAND2X1 NAND2X1_89 ( .A(_588_), .B(_592_), .Y(_277__48_) );
INVX1 INVX1_45 ( .A(1'b0), .Y(_596_) );
OR2X2 OR2X2_45 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_597_) );
NAND2X1 NAND2X1_90 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_598_) );
NAND3X1 NAND3X1_46 ( .A(_596_), .B(_598_), .C(_597_), .Y(_599_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_593_) );
AND2X2 AND2X2_46 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_594_) );
OAI21X1 OAI21X1_46 ( .A(_593_), .B(_594_), .C(1'b0), .Y(_595_) );
NAND2X1 NAND2X1_91 ( .A(_595_), .B(_599_), .Y(_277__0_) );
INVX1 INVX1_46 ( .A(w_C_1_), .Y(_603_) );
OR2X2 OR2X2_46 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_604_) );
NAND2X1 NAND2X1_92 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_605_) );
NAND3X1 NAND3X1_47 ( .A(_603_), .B(_605_), .C(_604_), .Y(_606_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_600_) );
AND2X2 AND2X2_47 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_601_) );
OAI21X1 OAI21X1_47 ( .A(_600_), .B(_601_), .C(w_C_1_), .Y(_602_) );
NAND2X1 NAND2X1_93 ( .A(_602_), .B(_606_), .Y(_277__1_) );
INVX1 INVX1_47 ( .A(w_C_2_), .Y(_610_) );
OR2X2 OR2X2_47 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_611_) );
NAND2X1 NAND2X1_94 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_612_) );
NAND3X1 NAND3X1_48 ( .A(_610_), .B(_612_), .C(_611_), .Y(_613_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_607_) );
AND2X2 AND2X2_48 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_608_) );
OAI21X1 OAI21X1_48 ( .A(_607_), .B(_608_), .C(w_C_2_), .Y(_609_) );
NAND2X1 NAND2X1_95 ( .A(_609_), .B(_613_), .Y(_277__2_) );
INVX1 INVX1_48 ( .A(w_C_3_), .Y(_617_) );
OR2X2 OR2X2_48 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_618_) );
NAND2X1 NAND2X1_96 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_619_) );
NAND3X1 NAND3X1_49 ( .A(_617_), .B(_619_), .C(_618_), .Y(_620_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_614_) );
AND2X2 AND2X2_49 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_615_) );
OAI21X1 OAI21X1_49 ( .A(_614_), .B(_615_), .C(w_C_3_), .Y(_616_) );
NAND2X1 NAND2X1_97 ( .A(_616_), .B(_620_), .Y(_277__3_) );
INVX1 INVX1_49 ( .A(_202_), .Y(_203_) );
NAND3X1 NAND3X1_50 ( .A(_201_), .B(_203_), .C(_199_), .Y(_204_) );
OAI21X1 OAI21X1_50 ( .A(i_add2[35]), .B(i_add1[35]), .C(_204_), .Y(_205_) );
INVX1 INVX1_50 ( .A(_205_), .Y(w_C_36_) );
INVX1 INVX1_51 ( .A(i_add2[36]), .Y(_206_) );
INVX1 INVX1_52 ( .A(i_add1[36]), .Y(_207_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_208_) );
INVX1 INVX1_53 ( .A(_208_), .Y(_209_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_210_) );
INVX1 INVX1_54 ( .A(_210_), .Y(_211_) );
NAND3X1 NAND3X1_51 ( .A(_209_), .B(_211_), .C(_204_), .Y(_212_) );
OAI21X1 OAI21X1_51 ( .A(_206_), .B(_207_), .C(_212_), .Y(w_C_37_) );
NOR2X1 NOR2X1_52 ( .A(_206_), .B(_207_), .Y(_213_) );
INVX1 INVX1_55 ( .A(_213_), .Y(_214_) );
AND2X2 AND2X2_50 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_215_) );
INVX1 INVX1_56 ( .A(_215_), .Y(_216_) );
NAND3X1 NAND3X1_52 ( .A(_214_), .B(_216_), .C(_212_), .Y(_217_) );
OAI21X1 OAI21X1_52 ( .A(i_add2[37]), .B(i_add1[37]), .C(_217_), .Y(_218_) );
INVX1 INVX1_57 ( .A(_218_), .Y(w_C_38_) );
INVX1 INVX1_58 ( .A(i_add2[38]), .Y(_219_) );
INVX1 INVX1_59 ( .A(i_add1[38]), .Y(_220_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_221_) );
INVX1 INVX1_60 ( .A(_221_), .Y(_222_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_223_) );
INVX1 INVX1_61 ( .A(_223_), .Y(_224_) );
NAND3X1 NAND3X1_53 ( .A(_222_), .B(_224_), .C(_217_), .Y(_225_) );
OAI21X1 OAI21X1_53 ( .A(_219_), .B(_220_), .C(_225_), .Y(w_C_39_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_226_) );
INVX1 INVX1_62 ( .A(_226_), .Y(_227_) );
NOR2X1 NOR2X1_56 ( .A(_219_), .B(_220_), .Y(_228_) );
INVX1 INVX1_63 ( .A(_228_), .Y(_229_) );
NAND2X1 NAND2X1_98 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_230_) );
NAND3X1 NAND3X1_54 ( .A(_229_), .B(_230_), .C(_225_), .Y(_231_) );
AND2X2 AND2X2_51 ( .A(_231_), .B(_227_), .Y(w_C_40_) );
INVX1 INVX1_64 ( .A(i_add2[40]), .Y(_232_) );
INVX1 INVX1_65 ( .A(i_add1[40]), .Y(_233_) );
NAND2X1 NAND2X1_99 ( .A(_232_), .B(_233_), .Y(_234_) );
NAND3X1 NAND3X1_55 ( .A(_227_), .B(_234_), .C(_231_), .Y(_235_) );
OAI21X1 OAI21X1_54 ( .A(_232_), .B(_233_), .C(_235_), .Y(w_C_41_) );
INVX1 INVX1_66 ( .A(i_add2[41]), .Y(_236_) );
INVX1 INVX1_67 ( .A(i_add1[41]), .Y(_237_) );
OAI21X1 OAI21X1_55 ( .A(i_add2[41]), .B(i_add1[41]), .C(w_C_41_), .Y(_238_) );
OAI21X1 OAI21X1_56 ( .A(_236_), .B(_237_), .C(_238_), .Y(w_C_42_) );
INVX1 INVX1_68 ( .A(i_add2[42]), .Y(_239_) );
INVX1 INVX1_69 ( .A(i_add1[42]), .Y(_240_) );
NOR2X1 NOR2X1_57 ( .A(_239_), .B(_240_), .Y(_241_) );
OR2X2 OR2X2_49 ( .A(w_C_42_), .B(_241_), .Y(_242_) );
OAI21X1 OAI21X1_57 ( .A(i_add2[42]), .B(i_add1[42]), .C(_242_), .Y(_243_) );
INVX1 INVX1_70 ( .A(_243_), .Y(w_C_43_) );
INVX1 INVX1_71 ( .A(_241_), .Y(_244_) );
NAND2X1 NAND2X1_100 ( .A(_236_), .B(_237_), .Y(_245_) );
NAND2X1 NAND2X1_101 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_246_) );
NAND2X1 NAND2X1_102 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_247_) );
NAND3X1 NAND3X1_56 ( .A(_246_), .B(_247_), .C(_235_), .Y(_248_) );
NAND2X1 NAND2X1_103 ( .A(_239_), .B(_240_), .Y(_249_) );
NAND3X1 NAND3X1_57 ( .A(_245_), .B(_249_), .C(_248_), .Y(_250_) );
NAND2X1 NAND2X1_104 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_251_) );
NAND3X1 NAND3X1_58 ( .A(_244_), .B(_251_), .C(_250_), .Y(_252_) );
OAI21X1 OAI21X1_58 ( .A(i_add2[43]), .B(i_add1[43]), .C(_252_), .Y(_253_) );
INVX1 INVX1_72 ( .A(_253_), .Y(w_C_44_) );
INVX1 INVX1_73 ( .A(i_add2[44]), .Y(_254_) );
INVX1 INVX1_74 ( .A(i_add1[44]), .Y(_255_) );
OAI21X1 OAI21X1_59 ( .A(_254_), .B(_255_), .C(_253_), .Y(_256_) );
OAI21X1 OAI21X1_60 ( .A(i_add2[44]), .B(i_add1[44]), .C(_256_), .Y(_257_) );
INVX1 INVX1_75 ( .A(_257_), .Y(w_C_45_) );
NAND2X1 NAND2X1_105 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_258_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_259_) );
OAI21X1 OAI21X1_61 ( .A(_259_), .B(_257_), .C(_258_), .Y(w_C_46_) );
NAND2X1 NAND2X1_106 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_260_) );
INVX1 INVX1_76 ( .A(_259_), .Y(_261_) );
NOR2X1 NOR2X1_59 ( .A(_254_), .B(_255_), .Y(_262_) );
INVX1 INVX1_77 ( .A(_262_), .Y(_263_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_264_) );
INVX1 INVX1_78 ( .A(_264_), .Y(_265_) );
NAND2X1 NAND2X1_107 ( .A(_254_), .B(_255_), .Y(_266_) );
NAND3X1 NAND3X1_59 ( .A(_265_), .B(_266_), .C(_252_), .Y(_267_) );
NAND3X1 NAND3X1_60 ( .A(_263_), .B(_258_), .C(_267_), .Y(_268_) );
OR2X2 OR2X2_50 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_269_) );
NAND3X1 NAND3X1_61 ( .A(_261_), .B(_269_), .C(_268_), .Y(_270_) );
NAND2X1 NAND2X1_108 ( .A(_260_), .B(_270_), .Y(w_C_47_) );
OR2X2 OR2X2_51 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_271_) );
NAND2X1 NAND2X1_109 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_272_) );
NAND3X1 NAND3X1_62 ( .A(_260_), .B(_272_), .C(_270_), .Y(_273_) );
AND2X2 AND2X2_52 ( .A(_273_), .B(_271_), .Y(w_C_48_) );
NAND2X1 NAND2X1_110 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_274_) );
OR2X2 OR2X2_52 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_275_) );
NAND3X1 NAND3X1_63 ( .A(_271_), .B(_275_), .C(_273_), .Y(_276_) );
NAND2X1 NAND2X1_111 ( .A(_274_), .B(_276_), .Y(w_C_49_) );
NAND2X1 NAND2X1_112 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_79 ( .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_113 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_114 ( .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_62 ( .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_80 ( .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_115 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_53 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_54 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_64 ( .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_116 ( .A(_4_), .B(_7_), .Y(w_C_3_) );
OR2X2 OR2X2_55 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
NAND2X1 NAND2X1_117 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_65 ( .A(_4_), .B(_9_), .C(_7_), .Y(_10_) );
AND2X2 AND2X2_53 ( .A(_10_), .B(_8_), .Y(w_C_4_) );
NAND2X1 NAND2X1_118 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
OR2X2 OR2X2_56 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_12_) );
NAND3X1 NAND3X1_66 ( .A(_8_), .B(_12_), .C(_10_), .Y(_13_) );
NAND2X1 NAND2X1_119 ( .A(_11_), .B(_13_), .Y(w_C_5_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_14_) );
INVX1 INVX1_81 ( .A(_14_), .Y(_15_) );
NAND2X1 NAND2X1_120 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_16_) );
NAND3X1 NAND3X1_67 ( .A(_11_), .B(_16_), .C(_13_), .Y(_17_) );
AND2X2 AND2X2_54 ( .A(_17_), .B(_15_), .Y(w_C_6_) );
AND2X2 AND2X2_55 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_18_) );
INVX1 INVX1_82 ( .A(_18_), .Y(_19_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_20_) );
INVX1 INVX1_83 ( .A(_20_), .Y(_21_) );
NAND3X1 NAND3X1_68 ( .A(_15_), .B(_21_), .C(_17_), .Y(_22_) );
AND2X2 AND2X2_56 ( .A(_22_), .B(_19_), .Y(_23_) );
INVX1 INVX1_84 ( .A(_23_), .Y(w_C_7_) );
AND2X2 AND2X2_57 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_24_) );
INVX1 INVX1_85 ( .A(_24_), .Y(_25_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_26_) );
OAI21X1 OAI21X1_63 ( .A(_26_), .B(_23_), .C(_25_), .Y(w_C_8_) );
AND2X2 AND2X2_58 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_27_) );
INVX1 INVX1_86 ( .A(_27_), .Y(_28_) );
INVX1 INVX1_87 ( .A(_26_), .Y(_29_) );
NAND3X1 NAND3X1_69 ( .A(_19_), .B(_25_), .C(_22_), .Y(_30_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_31_) );
INVX1 INVX1_88 ( .A(_31_), .Y(_32_) );
NAND3X1 NAND3X1_70 ( .A(_29_), .B(_32_), .C(_30_), .Y(_33_) );
AND2X2 AND2X2_59 ( .A(_33_), .B(_28_), .Y(_34_) );
INVX1 INVX1_89 ( .A(_34_), .Y(w_C_9_) );
AND2X2 AND2X2_60 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_35_) );
INVX1 INVX1_90 ( .A(_35_), .Y(_36_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_37_) );
OAI21X1 OAI21X1_64 ( .A(_37_), .B(_34_), .C(_36_), .Y(w_C_10_) );
AND2X2 AND2X2_61 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_38_) );
INVX1 INVX1_91 ( .A(_38_), .Y(_39_) );
INVX1 INVX1_92 ( .A(_37_), .Y(_40_) );
NAND3X1 NAND3X1_71 ( .A(_28_), .B(_36_), .C(_33_), .Y(_41_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_42_) );
INVX1 INVX1_93 ( .A(_42_), .Y(_43_) );
NAND3X1 NAND3X1_72 ( .A(_40_), .B(_43_), .C(_41_), .Y(_44_) );
AND2X2 AND2X2_62 ( .A(_44_), .B(_39_), .Y(_45_) );
INVX1 INVX1_94 ( .A(_45_), .Y(w_C_11_) );
AND2X2 AND2X2_63 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_46_) );
INVX1 INVX1_95 ( .A(_46_), .Y(_47_) );
NAND3X1 NAND3X1_73 ( .A(_39_), .B(_47_), .C(_44_), .Y(_48_) );
OAI21X1 OAI21X1_65 ( .A(i_add2[11]), .B(i_add1[11]), .C(_48_), .Y(_49_) );
INVX1 INVX1_96 ( .A(_49_), .Y(w_C_12_) );
INVX1 INVX1_97 ( .A(i_add2[12]), .Y(_50_) );
INVX1 INVX1_98 ( .A(i_add1[12]), .Y(_51_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_52_) );
INVX1 INVX1_99 ( .A(_52_), .Y(_53_) );
NOR2X1 NOR2X1_68 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_54_) );
INVX1 INVX1_100 ( .A(_54_), .Y(_55_) );
NAND3X1 NAND3X1_74 ( .A(_53_), .B(_55_), .C(_48_), .Y(_56_) );
OAI21X1 OAI21X1_66 ( .A(_50_), .B(_51_), .C(_56_), .Y(w_C_13_) );
NOR2X1 NOR2X1_69 ( .A(_50_), .B(_51_), .Y(_57_) );
INVX1 INVX1_101 ( .A(_57_), .Y(_58_) );
AND2X2 AND2X2_64 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_59_) );
INVX1 INVX1_102 ( .A(_59_), .Y(_60_) );
NAND3X1 NAND3X1_75 ( .A(_58_), .B(_60_), .C(_56_), .Y(_61_) );
OAI21X1 OAI21X1_67 ( .A(i_add2[13]), .B(i_add1[13]), .C(_61_), .Y(_62_) );
INVX1 INVX1_103 ( .A(_62_), .Y(w_C_14_) );
INVX1 INVX1_104 ( .A(i_add2[14]), .Y(_63_) );
INVX1 INVX1_105 ( .A(i_add1[14]), .Y(_64_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_65_) );
INVX1 INVX1_106 ( .A(_65_), .Y(_66_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_67_) );
INVX1 INVX1_107 ( .A(_67_), .Y(_68_) );
NAND3X1 NAND3X1_76 ( .A(_66_), .B(_68_), .C(_61_), .Y(_69_) );
OAI21X1 OAI21X1_68 ( .A(_63_), .B(_64_), .C(_69_), .Y(w_C_15_) );
NOR2X1 NOR2X1_72 ( .A(_63_), .B(_64_), .Y(_70_) );
INVX1 INVX1_108 ( .A(_70_), .Y(_71_) );
AND2X2 AND2X2_65 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_72_) );
INVX1 INVX1_109 ( .A(_72_), .Y(_73_) );
NAND3X1 NAND3X1_77 ( .A(_71_), .B(_73_), .C(_69_), .Y(_74_) );
OAI21X1 OAI21X1_69 ( .A(i_add2[15]), .B(i_add1[15]), .C(_74_), .Y(_75_) );
INVX1 INVX1_110 ( .A(_75_), .Y(w_C_16_) );
INVX1 INVX1_111 ( .A(i_add2[16]), .Y(_76_) );
INVX1 INVX1_112 ( .A(i_add1[16]), .Y(_77_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_78_) );
INVX1 INVX1_113 ( .A(_78_), .Y(_79_) );
NOR2X1 NOR2X1_74 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_80_) );
INVX1 INVX1_114 ( .A(_80_), .Y(_81_) );
NAND3X1 NAND3X1_78 ( .A(_79_), .B(_81_), .C(_74_), .Y(_82_) );
OAI21X1 OAI21X1_70 ( .A(_76_), .B(_77_), .C(_82_), .Y(w_C_17_) );
NOR2X1 NOR2X1_75 ( .A(_76_), .B(_77_), .Y(_83_) );
INVX1 INVX1_115 ( .A(_83_), .Y(_84_) );
AND2X2 AND2X2_66 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_85_) );
INVX1 INVX1_116 ( .A(_85_), .Y(_86_) );
NAND3X1 NAND3X1_79 ( .A(_84_), .B(_86_), .C(_82_), .Y(_87_) );
OAI21X1 OAI21X1_71 ( .A(i_add2[17]), .B(i_add1[17]), .C(_87_), .Y(_88_) );
INVX1 INVX1_117 ( .A(_88_), .Y(w_C_18_) );
INVX1 INVX1_118 ( .A(i_add2[18]), .Y(_89_) );
INVX1 INVX1_119 ( .A(i_add1[18]), .Y(_90_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_91_) );
INVX1 INVX1_120 ( .A(_91_), .Y(_92_) );
NOR2X1 NOR2X1_77 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_93_) );
INVX1 INVX1_121 ( .A(_93_), .Y(_94_) );
NAND3X1 NAND3X1_80 ( .A(_92_), .B(_94_), .C(_87_), .Y(_95_) );
OAI21X1 OAI21X1_72 ( .A(_89_), .B(_90_), .C(_95_), .Y(w_C_19_) );
NOR2X1 NOR2X1_78 ( .A(_89_), .B(_90_), .Y(_96_) );
INVX1 INVX1_122 ( .A(_96_), .Y(_97_) );
AND2X2 AND2X2_67 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_98_) );
INVX1 INVX1_123 ( .A(_98_), .Y(_99_) );
NAND3X1 NAND3X1_81 ( .A(_97_), .B(_99_), .C(_95_), .Y(_100_) );
OAI21X1 OAI21X1_73 ( .A(i_add2[19]), .B(i_add1[19]), .C(_100_), .Y(_101_) );
INVX1 INVX1_124 ( .A(_101_), .Y(w_C_20_) );
INVX1 INVX1_125 ( .A(i_add2[20]), .Y(_102_) );
INVX1 INVX1_126 ( .A(i_add1[20]), .Y(_103_) );
NOR2X1 NOR2X1_79 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_104_) );
INVX1 INVX1_127 ( .A(_104_), .Y(_105_) );
NOR2X1 NOR2X1_80 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_106_) );
INVX1 INVX1_128 ( .A(_106_), .Y(_107_) );
NAND3X1 NAND3X1_82 ( .A(_105_), .B(_107_), .C(_100_), .Y(_108_) );
OAI21X1 OAI21X1_74 ( .A(_102_), .B(_103_), .C(_108_), .Y(w_C_21_) );
NOR2X1 NOR2X1_81 ( .A(_102_), .B(_103_), .Y(_109_) );
INVX1 INVX1_129 ( .A(_109_), .Y(_110_) );
AND2X2 AND2X2_68 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_111_) );
INVX1 INVX1_130 ( .A(_111_), .Y(_112_) );
NAND3X1 NAND3X1_83 ( .A(_110_), .B(_112_), .C(_108_), .Y(_113_) );
OAI21X1 OAI21X1_75 ( .A(i_add2[21]), .B(i_add1[21]), .C(_113_), .Y(_114_) );
INVX1 INVX1_131 ( .A(_114_), .Y(w_C_22_) );
INVX1 INVX1_132 ( .A(i_add2[22]), .Y(_115_) );
INVX1 INVX1_133 ( .A(i_add1[22]), .Y(_116_) );
NOR2X1 NOR2X1_82 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_117_) );
INVX1 INVX1_134 ( .A(_117_), .Y(_118_) );
NOR2X1 NOR2X1_83 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_119_) );
INVX1 INVX1_135 ( .A(_119_), .Y(_120_) );
NAND3X1 NAND3X1_84 ( .A(_118_), .B(_120_), .C(_113_), .Y(_121_) );
OAI21X1 OAI21X1_76 ( .A(_115_), .B(_116_), .C(_121_), .Y(w_C_23_) );
NOR2X1 NOR2X1_84 ( .A(_115_), .B(_116_), .Y(_122_) );
INVX1 INVX1_136 ( .A(_122_), .Y(_123_) );
AND2X2 AND2X2_69 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_124_) );
INVX1 INVX1_137 ( .A(_124_), .Y(_125_) );
NAND3X1 NAND3X1_85 ( .A(_123_), .B(_125_), .C(_121_), .Y(_126_) );
OAI21X1 OAI21X1_77 ( .A(i_add2[23]), .B(i_add1[23]), .C(_126_), .Y(_127_) );
INVX1 INVX1_138 ( .A(_127_), .Y(w_C_24_) );
INVX1 INVX1_139 ( .A(i_add2[24]), .Y(_128_) );
INVX1 INVX1_140 ( .A(i_add1[24]), .Y(_129_) );
NOR2X1 NOR2X1_85 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_130_) );
INVX1 INVX1_141 ( .A(_130_), .Y(_131_) );
NOR2X1 NOR2X1_86 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_132_) );
INVX1 INVX1_142 ( .A(_132_), .Y(_133_) );
NAND3X1 NAND3X1_86 ( .A(_131_), .B(_133_), .C(_126_), .Y(_134_) );
OAI21X1 OAI21X1_78 ( .A(_128_), .B(_129_), .C(_134_), .Y(w_C_25_) );
NOR2X1 NOR2X1_87 ( .A(_128_), .B(_129_), .Y(_135_) );
INVX1 INVX1_143 ( .A(_135_), .Y(_136_) );
AND2X2 AND2X2_70 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_137_) );
INVX1 INVX1_144 ( .A(_137_), .Y(_138_) );
NAND3X1 NAND3X1_87 ( .A(_136_), .B(_138_), .C(_134_), .Y(_139_) );
OAI21X1 OAI21X1_79 ( .A(i_add2[25]), .B(i_add1[25]), .C(_139_), .Y(_140_) );
INVX1 INVX1_145 ( .A(_140_), .Y(w_C_26_) );
INVX1 INVX1_146 ( .A(i_add2[26]), .Y(_141_) );
INVX1 INVX1_147 ( .A(i_add1[26]), .Y(_142_) );
NOR2X1 NOR2X1_88 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_143_) );
INVX1 INVX1_148 ( .A(_143_), .Y(_144_) );
NOR2X1 NOR2X1_89 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_145_) );
INVX1 INVX1_149 ( .A(_145_), .Y(_146_) );
NAND3X1 NAND3X1_88 ( .A(_144_), .B(_146_), .C(_139_), .Y(_147_) );
OAI21X1 OAI21X1_80 ( .A(_141_), .B(_142_), .C(_147_), .Y(w_C_27_) );
NOR2X1 NOR2X1_90 ( .A(_141_), .B(_142_), .Y(_148_) );
INVX1 INVX1_150 ( .A(_148_), .Y(_149_) );
AND2X2 AND2X2_71 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_150_) );
INVX1 INVX1_151 ( .A(_150_), .Y(_151_) );
NAND3X1 NAND3X1_89 ( .A(_149_), .B(_151_), .C(_147_), .Y(_152_) );
OAI21X1 OAI21X1_81 ( .A(i_add2[27]), .B(i_add1[27]), .C(_152_), .Y(_153_) );
INVX1 INVX1_152 ( .A(_153_), .Y(w_C_28_) );
INVX1 INVX1_153 ( .A(i_add2[28]), .Y(_154_) );
INVX1 INVX1_154 ( .A(i_add1[28]), .Y(_155_) );
NOR2X1 NOR2X1_91 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_156_) );
INVX1 INVX1_155 ( .A(_156_), .Y(_157_) );
NOR2X1 NOR2X1_92 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_158_) );
INVX1 INVX1_156 ( .A(_158_), .Y(_159_) );
NAND3X1 NAND3X1_90 ( .A(_157_), .B(_159_), .C(_152_), .Y(_160_) );
OAI21X1 OAI21X1_82 ( .A(_154_), .B(_155_), .C(_160_), .Y(w_C_29_) );
NOR2X1 NOR2X1_93 ( .A(_154_), .B(_155_), .Y(_161_) );
INVX1 INVX1_157 ( .A(_161_), .Y(_162_) );
AND2X2 AND2X2_72 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_163_) );
INVX1 INVX1_158 ( .A(_163_), .Y(_164_) );
NAND3X1 NAND3X1_91 ( .A(_162_), .B(_164_), .C(_160_), .Y(_165_) );
OAI21X1 OAI21X1_83 ( .A(i_add2[29]), .B(i_add1[29]), .C(_165_), .Y(_166_) );
INVX1 INVX1_159 ( .A(_166_), .Y(w_C_30_) );
INVX1 INVX1_160 ( .A(i_add2[30]), .Y(_167_) );
INVX1 INVX1_161 ( .A(i_add1[30]), .Y(_168_) );
NOR2X1 NOR2X1_94 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_169_) );
INVX1 INVX1_162 ( .A(_169_), .Y(_170_) );
NOR2X1 NOR2X1_95 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_171_) );
INVX1 INVX1_163 ( .A(_171_), .Y(_172_) );
NAND3X1 NAND3X1_92 ( .A(_170_), .B(_172_), .C(_165_), .Y(_173_) );
OAI21X1 OAI21X1_84 ( .A(_167_), .B(_168_), .C(_173_), .Y(w_C_31_) );
NOR2X1 NOR2X1_96 ( .A(_167_), .B(_168_), .Y(_174_) );
INVX1 INVX1_164 ( .A(_174_), .Y(_175_) );
AND2X2 AND2X2_73 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_176_) );
INVX1 INVX1_165 ( .A(_176_), .Y(_177_) );
NAND3X1 NAND3X1_93 ( .A(_175_), .B(_177_), .C(_173_), .Y(_178_) );
OAI21X1 OAI21X1_85 ( .A(i_add2[31]), .B(i_add1[31]), .C(_178_), .Y(_179_) );
INVX1 INVX1_166 ( .A(_179_), .Y(w_C_32_) );
INVX1 INVX1_167 ( .A(i_add2[32]), .Y(_180_) );
INVX1 INVX1_168 ( .A(i_add1[32]), .Y(_181_) );
NOR2X1 NOR2X1_97 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_182_) );
INVX1 INVX1_169 ( .A(_182_), .Y(_183_) );
NOR2X1 NOR2X1_98 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_184_) );
INVX1 INVX1_170 ( .A(_184_), .Y(_185_) );
NAND3X1 NAND3X1_94 ( .A(_183_), .B(_185_), .C(_178_), .Y(_186_) );
OAI21X1 OAI21X1_86 ( .A(_180_), .B(_181_), .C(_186_), .Y(w_C_33_) );
NOR2X1 NOR2X1_99 ( .A(_180_), .B(_181_), .Y(_187_) );
INVX1 INVX1_171 ( .A(_187_), .Y(_188_) );
AND2X2 AND2X2_74 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_189_) );
INVX1 INVX1_172 ( .A(_189_), .Y(_190_) );
NAND3X1 NAND3X1_95 ( .A(_188_), .B(_190_), .C(_186_), .Y(_191_) );
OAI21X1 OAI21X1_87 ( .A(i_add2[33]), .B(i_add1[33]), .C(_191_), .Y(_192_) );
INVX1 INVX1_173 ( .A(_192_), .Y(w_C_34_) );
INVX1 INVX1_174 ( .A(i_add2[34]), .Y(_193_) );
INVX1 INVX1_175 ( .A(i_add1[34]), .Y(_194_) );
NOR2X1 NOR2X1_100 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_195_) );
INVX1 INVX1_176 ( .A(_195_), .Y(_196_) );
NOR2X1 NOR2X1_101 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_197_) );
INVX1 INVX1_177 ( .A(_197_), .Y(_198_) );
NAND3X1 NAND3X1_96 ( .A(_196_), .B(_198_), .C(_191_), .Y(_199_) );
OAI21X1 OAI21X1_88 ( .A(_193_), .B(_194_), .C(_199_), .Y(w_C_35_) );
NOR2X1 NOR2X1_102 ( .A(_193_), .B(_194_), .Y(_200_) );
INVX1 INVX1_178 ( .A(_200_), .Y(_201_) );
AND2X2 AND2X2_75 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_202_) );
BUFX2 BUFX2_1 ( .A(_277__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_277__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_277__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_277__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_277__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_277__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_277__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_277__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_277__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_277__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_277__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_277__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_277__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_277__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_277__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_277__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_277__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_277__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_277__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_277__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_277__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_277__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_277__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_277__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_277__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_277__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_277__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_277__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_277__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_277__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_277__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_277__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_277__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_277__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_277__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_277__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_277__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(_277__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .A(_277__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .A(_277__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .A(_277__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .A(_277__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .A(_277__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .A(_277__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .A(_277__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .A(_277__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .A(_277__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .A(_277__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .A(_277__48_), .Y(o_result[48]) );
BUFX2 BUFX2_50 ( .A(w_C_49_), .Y(o_result[49]) );
INVX1 INVX1_179 ( .A(w_C_4_), .Y(_281_) );
OR2X2 OR2X2_57 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_282_) );
NAND2X1 NAND2X1_121 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_283_) );
BUFX2 BUFX2_51 ( .A(w_C_49_), .Y(_277__49_) );
BUFX2 BUFX2_52 ( .A(1'b0), .Y(w_C_0_) );
endmodule
