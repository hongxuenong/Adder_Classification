module rca_41bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21], o_result[22], o_result[23], o_result[24], o_result[25], o_result[26], o_result[27], o_result[28], o_result[29], o_result[30], o_result[31], o_result[32], o_result[33], o_result[34], o_result[35], o_result[36], o_result[37], o_result[38], o_result[39], o_result[40], o_result[41]);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];
output o_result[22];
output o_result[23];
output o_result[24];
output o_result[25];
output o_result[26];
output o_result[27];
output o_result[28];
output o_result[29];
output o_result[30];
output o_result[31];
output o_result[32];
output o_result[33];
output o_result[34];
output o_result[35];
output o_result[36];
output o_result[37];
output o_result[38];
output o_result[39];
output o_result[40];
output o_result[41];

BUFX2 BUFX2_1 ( .A(_0__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_0__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_0__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_0__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_0__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_0__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_0__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_0__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_0__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_0__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_0__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_0__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_0__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_0__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_0__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_0__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_0__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_0__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_0__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_0__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_0__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_0__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_0__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_0__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_0__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_0__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_0__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_0__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_0__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_0__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_0__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_0__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_0__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_0__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_0__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_0__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_0__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(_0__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .A(_0__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .A(_0__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .A(_0__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .A(w_CARRY_41_), .Y(o_result[41]) );
INVX1 INVX1_1 ( .A(w_CARRY_4_), .Y(_5_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_6_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_7_) );
OAI21X1 OAI21X1_1 ( .A(_5_), .B(_7_), .C(_6_), .Y(w_CARRY_5_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_1_) );
NAND3X1 NAND3X1_1 ( .A(_5_), .B(_6_), .C(_1_), .Y(_2_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_3_) );
OAI21X1 OAI21X1_2 ( .A(_7_), .B(_3_), .C(w_CARRY_4_), .Y(_4_) );
NAND2X1 NAND2X1_2 ( .A(_4_), .B(_2_), .Y(_0__4_) );
INVX1 INVX1_2 ( .A(w_CARRY_5_), .Y(_12_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_13_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_14_) );
OAI21X1 OAI21X1_3 ( .A(_12_), .B(_14_), .C(_13_), .Y(w_CARRY_6_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_8_) );
NAND3X1 NAND3X1_2 ( .A(_12_), .B(_13_), .C(_8_), .Y(_9_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_10_) );
OAI21X1 OAI21X1_4 ( .A(_14_), .B(_10_), .C(w_CARRY_5_), .Y(_11_) );
NAND2X1 NAND2X1_4 ( .A(_11_), .B(_9_), .Y(_0__5_) );
INVX1 INVX1_3 ( .A(w_CARRY_6_), .Y(_19_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_20_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_21_) );
OAI21X1 OAI21X1_5 ( .A(_19_), .B(_21_), .C(_20_), .Y(w_CARRY_7_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_15_) );
NAND3X1 NAND3X1_3 ( .A(_19_), .B(_20_), .C(_15_), .Y(_16_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_17_) );
OAI21X1 OAI21X1_6 ( .A(_21_), .B(_17_), .C(w_CARRY_6_), .Y(_18_) );
NAND2X1 NAND2X1_6 ( .A(_18_), .B(_16_), .Y(_0__6_) );
INVX1 INVX1_4 ( .A(w_CARRY_7_), .Y(_26_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_27_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_28_) );
OAI21X1 OAI21X1_7 ( .A(_26_), .B(_28_), .C(_27_), .Y(w_CARRY_8_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_22_) );
NAND3X1 NAND3X1_4 ( .A(_26_), .B(_27_), .C(_22_), .Y(_23_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_24_) );
OAI21X1 OAI21X1_8 ( .A(_28_), .B(_24_), .C(w_CARRY_7_), .Y(_25_) );
NAND2X1 NAND2X1_8 ( .A(_25_), .B(_23_), .Y(_0__7_) );
INVX1 INVX1_5 ( .A(w_CARRY_8_), .Y(_33_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_34_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_35_) );
OAI21X1 OAI21X1_9 ( .A(_33_), .B(_35_), .C(_34_), .Y(w_CARRY_9_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_29_) );
NAND3X1 NAND3X1_5 ( .A(_33_), .B(_34_), .C(_29_), .Y(_30_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_31_) );
OAI21X1 OAI21X1_10 ( .A(_35_), .B(_31_), .C(w_CARRY_8_), .Y(_32_) );
NAND2X1 NAND2X1_10 ( .A(_32_), .B(_30_), .Y(_0__8_) );
INVX1 INVX1_6 ( .A(w_CARRY_9_), .Y(_40_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_41_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_42_) );
OAI21X1 OAI21X1_11 ( .A(_40_), .B(_42_), .C(_41_), .Y(w_CARRY_10_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_36_) );
NAND3X1 NAND3X1_6 ( .A(_40_), .B(_41_), .C(_36_), .Y(_37_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_38_) );
OAI21X1 OAI21X1_12 ( .A(_42_), .B(_38_), .C(w_CARRY_9_), .Y(_39_) );
NAND2X1 NAND2X1_12 ( .A(_39_), .B(_37_), .Y(_0__9_) );
INVX1 INVX1_7 ( .A(w_CARRY_10_), .Y(_47_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_48_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_49_) );
OAI21X1 OAI21X1_13 ( .A(_47_), .B(_49_), .C(_48_), .Y(w_CARRY_11_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_43_) );
NAND3X1 NAND3X1_7 ( .A(_47_), .B(_48_), .C(_43_), .Y(_44_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_45_) );
OAI21X1 OAI21X1_14 ( .A(_49_), .B(_45_), .C(w_CARRY_10_), .Y(_46_) );
NAND2X1 NAND2X1_14 ( .A(_46_), .B(_44_), .Y(_0__10_) );
INVX1 INVX1_8 ( .A(w_CARRY_11_), .Y(_54_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_55_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_56_) );
OAI21X1 OAI21X1_15 ( .A(_54_), .B(_56_), .C(_55_), .Y(w_CARRY_12_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_50_) );
NAND3X1 NAND3X1_8 ( .A(_54_), .B(_55_), .C(_50_), .Y(_51_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_52_) );
OAI21X1 OAI21X1_16 ( .A(_56_), .B(_52_), .C(w_CARRY_11_), .Y(_53_) );
NAND2X1 NAND2X1_16 ( .A(_53_), .B(_51_), .Y(_0__11_) );
INVX1 INVX1_9 ( .A(w_CARRY_12_), .Y(_61_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_62_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_63_) );
OAI21X1 OAI21X1_17 ( .A(_61_), .B(_63_), .C(_62_), .Y(w_CARRY_13_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_57_) );
NAND3X1 NAND3X1_9 ( .A(_61_), .B(_62_), .C(_57_), .Y(_58_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_59_) );
OAI21X1 OAI21X1_18 ( .A(_63_), .B(_59_), .C(w_CARRY_12_), .Y(_60_) );
NAND2X1 NAND2X1_18 ( .A(_60_), .B(_58_), .Y(_0__12_) );
INVX1 INVX1_10 ( .A(w_CARRY_13_), .Y(_68_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_69_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_70_) );
OAI21X1 OAI21X1_19 ( .A(_68_), .B(_70_), .C(_69_), .Y(w_CARRY_14_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_64_) );
NAND3X1 NAND3X1_10 ( .A(_68_), .B(_69_), .C(_64_), .Y(_65_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_66_) );
OAI21X1 OAI21X1_20 ( .A(_70_), .B(_66_), .C(w_CARRY_13_), .Y(_67_) );
NAND2X1 NAND2X1_20 ( .A(_67_), .B(_65_), .Y(_0__13_) );
INVX1 INVX1_11 ( .A(w_CARRY_14_), .Y(_75_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_76_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_77_) );
OAI21X1 OAI21X1_21 ( .A(_75_), .B(_77_), .C(_76_), .Y(w_CARRY_15_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_71_) );
NAND3X1 NAND3X1_11 ( .A(_75_), .B(_76_), .C(_71_), .Y(_72_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_73_) );
OAI21X1 OAI21X1_22 ( .A(_77_), .B(_73_), .C(w_CARRY_14_), .Y(_74_) );
NAND2X1 NAND2X1_22 ( .A(_74_), .B(_72_), .Y(_0__14_) );
INVX1 INVX1_12 ( .A(w_CARRY_15_), .Y(_82_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_83_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_84_) );
OAI21X1 OAI21X1_23 ( .A(_82_), .B(_84_), .C(_83_), .Y(w_CARRY_16_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_78_) );
NAND3X1 NAND3X1_12 ( .A(_82_), .B(_83_), .C(_78_), .Y(_79_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_80_) );
OAI21X1 OAI21X1_24 ( .A(_84_), .B(_80_), .C(w_CARRY_15_), .Y(_81_) );
NAND2X1 NAND2X1_24 ( .A(_81_), .B(_79_), .Y(_0__15_) );
INVX1 INVX1_13 ( .A(w_CARRY_16_), .Y(_89_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_90_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_91_) );
OAI21X1 OAI21X1_25 ( .A(_89_), .B(_91_), .C(_90_), .Y(w_CARRY_17_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_85_) );
NAND3X1 NAND3X1_13 ( .A(_89_), .B(_90_), .C(_85_), .Y(_86_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_87_) );
OAI21X1 OAI21X1_26 ( .A(_91_), .B(_87_), .C(w_CARRY_16_), .Y(_88_) );
NAND2X1 NAND2X1_26 ( .A(_88_), .B(_86_), .Y(_0__16_) );
INVX1 INVX1_14 ( .A(w_CARRY_17_), .Y(_96_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_97_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_98_) );
OAI21X1 OAI21X1_27 ( .A(_96_), .B(_98_), .C(_97_), .Y(w_CARRY_18_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_92_) );
NAND3X1 NAND3X1_14 ( .A(_96_), .B(_97_), .C(_92_), .Y(_93_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_94_) );
OAI21X1 OAI21X1_28 ( .A(_98_), .B(_94_), .C(w_CARRY_17_), .Y(_95_) );
NAND2X1 NAND2X1_28 ( .A(_95_), .B(_93_), .Y(_0__17_) );
INVX1 INVX1_15 ( .A(w_CARRY_18_), .Y(_103_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_104_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_105_) );
OAI21X1 OAI21X1_29 ( .A(_103_), .B(_105_), .C(_104_), .Y(w_CARRY_19_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_99_) );
NAND3X1 NAND3X1_15 ( .A(_103_), .B(_104_), .C(_99_), .Y(_100_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_101_) );
OAI21X1 OAI21X1_30 ( .A(_105_), .B(_101_), .C(w_CARRY_18_), .Y(_102_) );
NAND2X1 NAND2X1_30 ( .A(_102_), .B(_100_), .Y(_0__18_) );
INVX1 INVX1_16 ( .A(w_CARRY_19_), .Y(_110_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_111_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_112_) );
OAI21X1 OAI21X1_31 ( .A(_110_), .B(_112_), .C(_111_), .Y(w_CARRY_20_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_106_) );
NAND3X1 NAND3X1_16 ( .A(_110_), .B(_111_), .C(_106_), .Y(_107_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_108_) );
OAI21X1 OAI21X1_32 ( .A(_112_), .B(_108_), .C(w_CARRY_19_), .Y(_109_) );
NAND2X1 NAND2X1_32 ( .A(_109_), .B(_107_), .Y(_0__19_) );
INVX1 INVX1_17 ( .A(w_CARRY_20_), .Y(_117_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_118_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_119_) );
OAI21X1 OAI21X1_33 ( .A(_117_), .B(_119_), .C(_118_), .Y(w_CARRY_21_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_113_) );
NAND3X1 NAND3X1_17 ( .A(_117_), .B(_118_), .C(_113_), .Y(_114_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_115_) );
OAI21X1 OAI21X1_34 ( .A(_119_), .B(_115_), .C(w_CARRY_20_), .Y(_116_) );
NAND2X1 NAND2X1_34 ( .A(_116_), .B(_114_), .Y(_0__20_) );
INVX1 INVX1_18 ( .A(w_CARRY_21_), .Y(_124_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_125_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_126_) );
OAI21X1 OAI21X1_35 ( .A(_124_), .B(_126_), .C(_125_), .Y(w_CARRY_22_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_120_) );
NAND3X1 NAND3X1_18 ( .A(_124_), .B(_125_), .C(_120_), .Y(_121_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_122_) );
OAI21X1 OAI21X1_36 ( .A(_126_), .B(_122_), .C(w_CARRY_21_), .Y(_123_) );
NAND2X1 NAND2X1_36 ( .A(_123_), .B(_121_), .Y(_0__21_) );
INVX1 INVX1_19 ( .A(w_CARRY_22_), .Y(_131_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_132_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_133_) );
OAI21X1 OAI21X1_37 ( .A(_131_), .B(_133_), .C(_132_), .Y(w_CARRY_23_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_127_) );
NAND3X1 NAND3X1_19 ( .A(_131_), .B(_132_), .C(_127_), .Y(_128_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_129_) );
OAI21X1 OAI21X1_38 ( .A(_133_), .B(_129_), .C(w_CARRY_22_), .Y(_130_) );
NAND2X1 NAND2X1_38 ( .A(_130_), .B(_128_), .Y(_0__22_) );
INVX1 INVX1_20 ( .A(w_CARRY_23_), .Y(_138_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_139_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_140_) );
OAI21X1 OAI21X1_39 ( .A(_138_), .B(_140_), .C(_139_), .Y(w_CARRY_24_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_134_) );
NAND3X1 NAND3X1_20 ( .A(_138_), .B(_139_), .C(_134_), .Y(_135_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_136_) );
OAI21X1 OAI21X1_40 ( .A(_140_), .B(_136_), .C(w_CARRY_23_), .Y(_137_) );
NAND2X1 NAND2X1_40 ( .A(_137_), .B(_135_), .Y(_0__23_) );
INVX1 INVX1_21 ( .A(w_CARRY_24_), .Y(_145_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_146_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_147_) );
OAI21X1 OAI21X1_41 ( .A(_145_), .B(_147_), .C(_146_), .Y(w_CARRY_25_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_141_) );
NAND3X1 NAND3X1_21 ( .A(_145_), .B(_146_), .C(_141_), .Y(_142_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_143_) );
OAI21X1 OAI21X1_42 ( .A(_147_), .B(_143_), .C(w_CARRY_24_), .Y(_144_) );
NAND2X1 NAND2X1_42 ( .A(_144_), .B(_142_), .Y(_0__24_) );
INVX1 INVX1_22 ( .A(w_CARRY_25_), .Y(_152_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_153_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_154_) );
OAI21X1 OAI21X1_43 ( .A(_152_), .B(_154_), .C(_153_), .Y(w_CARRY_26_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_148_) );
NAND3X1 NAND3X1_22 ( .A(_152_), .B(_153_), .C(_148_), .Y(_149_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_150_) );
OAI21X1 OAI21X1_44 ( .A(_154_), .B(_150_), .C(w_CARRY_25_), .Y(_151_) );
NAND2X1 NAND2X1_44 ( .A(_151_), .B(_149_), .Y(_0__25_) );
INVX1 INVX1_23 ( .A(w_CARRY_26_), .Y(_159_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_160_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_161_) );
OAI21X1 OAI21X1_45 ( .A(_159_), .B(_161_), .C(_160_), .Y(w_CARRY_27_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_155_) );
NAND3X1 NAND3X1_23 ( .A(_159_), .B(_160_), .C(_155_), .Y(_156_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_157_) );
OAI21X1 OAI21X1_46 ( .A(_161_), .B(_157_), .C(w_CARRY_26_), .Y(_158_) );
NAND2X1 NAND2X1_46 ( .A(_158_), .B(_156_), .Y(_0__26_) );
INVX1 INVX1_24 ( .A(w_CARRY_27_), .Y(_166_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_167_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_168_) );
OAI21X1 OAI21X1_47 ( .A(_166_), .B(_168_), .C(_167_), .Y(w_CARRY_28_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_162_) );
NAND3X1 NAND3X1_24 ( .A(_166_), .B(_167_), .C(_162_), .Y(_163_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_164_) );
OAI21X1 OAI21X1_48 ( .A(_168_), .B(_164_), .C(w_CARRY_27_), .Y(_165_) );
NAND2X1 NAND2X1_48 ( .A(_165_), .B(_163_), .Y(_0__27_) );
INVX1 INVX1_25 ( .A(w_CARRY_28_), .Y(_173_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_174_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_175_) );
OAI21X1 OAI21X1_49 ( .A(_173_), .B(_175_), .C(_174_), .Y(w_CARRY_29_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_169_) );
NAND3X1 NAND3X1_25 ( .A(_173_), .B(_174_), .C(_169_), .Y(_170_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_171_) );
OAI21X1 OAI21X1_50 ( .A(_175_), .B(_171_), .C(w_CARRY_28_), .Y(_172_) );
NAND2X1 NAND2X1_50 ( .A(_172_), .B(_170_), .Y(_0__28_) );
INVX1 INVX1_26 ( .A(w_CARRY_29_), .Y(_180_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_181_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_182_) );
OAI21X1 OAI21X1_51 ( .A(_180_), .B(_182_), .C(_181_), .Y(w_CARRY_30_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_176_) );
NAND3X1 NAND3X1_26 ( .A(_180_), .B(_181_), .C(_176_), .Y(_177_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_178_) );
OAI21X1 OAI21X1_52 ( .A(_182_), .B(_178_), .C(w_CARRY_29_), .Y(_179_) );
NAND2X1 NAND2X1_52 ( .A(_179_), .B(_177_), .Y(_0__29_) );
INVX1 INVX1_27 ( .A(w_CARRY_30_), .Y(_187_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_188_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_189_) );
OAI21X1 OAI21X1_53 ( .A(_187_), .B(_189_), .C(_188_), .Y(w_CARRY_31_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_183_) );
NAND3X1 NAND3X1_27 ( .A(_187_), .B(_188_), .C(_183_), .Y(_184_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_185_) );
OAI21X1 OAI21X1_54 ( .A(_189_), .B(_185_), .C(w_CARRY_30_), .Y(_186_) );
NAND2X1 NAND2X1_54 ( .A(_186_), .B(_184_), .Y(_0__30_) );
INVX1 INVX1_28 ( .A(w_CARRY_31_), .Y(_194_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_195_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_196_) );
OAI21X1 OAI21X1_55 ( .A(_194_), .B(_196_), .C(_195_), .Y(w_CARRY_32_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_190_) );
NAND3X1 NAND3X1_28 ( .A(_194_), .B(_195_), .C(_190_), .Y(_191_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_192_) );
OAI21X1 OAI21X1_56 ( .A(_196_), .B(_192_), .C(w_CARRY_31_), .Y(_193_) );
NAND2X1 NAND2X1_56 ( .A(_193_), .B(_191_), .Y(_0__31_) );
INVX1 INVX1_29 ( .A(w_CARRY_32_), .Y(_201_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_202_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_203_) );
OAI21X1 OAI21X1_57 ( .A(_201_), .B(_203_), .C(_202_), .Y(w_CARRY_33_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_197_) );
NAND3X1 NAND3X1_29 ( .A(_201_), .B(_202_), .C(_197_), .Y(_198_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_199_) );
OAI21X1 OAI21X1_58 ( .A(_203_), .B(_199_), .C(w_CARRY_32_), .Y(_200_) );
NAND2X1 NAND2X1_58 ( .A(_200_), .B(_198_), .Y(_0__32_) );
INVX1 INVX1_30 ( .A(w_CARRY_33_), .Y(_208_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_209_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_210_) );
OAI21X1 OAI21X1_59 ( .A(_208_), .B(_210_), .C(_209_), .Y(w_CARRY_34_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_204_) );
NAND3X1 NAND3X1_30 ( .A(_208_), .B(_209_), .C(_204_), .Y(_205_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_206_) );
OAI21X1 OAI21X1_60 ( .A(_210_), .B(_206_), .C(w_CARRY_33_), .Y(_207_) );
NAND2X1 NAND2X1_60 ( .A(_207_), .B(_205_), .Y(_0__33_) );
INVX1 INVX1_31 ( .A(w_CARRY_34_), .Y(_215_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_216_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_217_) );
OAI21X1 OAI21X1_61 ( .A(_215_), .B(_217_), .C(_216_), .Y(w_CARRY_35_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_211_) );
NAND3X1 NAND3X1_31 ( .A(_215_), .B(_216_), .C(_211_), .Y(_212_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_213_) );
OAI21X1 OAI21X1_62 ( .A(_217_), .B(_213_), .C(w_CARRY_34_), .Y(_214_) );
NAND2X1 NAND2X1_62 ( .A(_214_), .B(_212_), .Y(_0__34_) );
INVX1 INVX1_32 ( .A(w_CARRY_35_), .Y(_222_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_223_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_224_) );
OAI21X1 OAI21X1_63 ( .A(_222_), .B(_224_), .C(_223_), .Y(w_CARRY_36_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_218_) );
NAND3X1 NAND3X1_32 ( .A(_222_), .B(_223_), .C(_218_), .Y(_219_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_220_) );
OAI21X1 OAI21X1_64 ( .A(_224_), .B(_220_), .C(w_CARRY_35_), .Y(_221_) );
NAND2X1 NAND2X1_64 ( .A(_221_), .B(_219_), .Y(_0__35_) );
INVX1 INVX1_33 ( .A(w_CARRY_36_), .Y(_229_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_230_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_231_) );
OAI21X1 OAI21X1_65 ( .A(_229_), .B(_231_), .C(_230_), .Y(w_CARRY_37_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_225_) );
NAND3X1 NAND3X1_33 ( .A(_229_), .B(_230_), .C(_225_), .Y(_226_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_227_) );
OAI21X1 OAI21X1_66 ( .A(_231_), .B(_227_), .C(w_CARRY_36_), .Y(_228_) );
NAND2X1 NAND2X1_66 ( .A(_228_), .B(_226_), .Y(_0__36_) );
INVX1 INVX1_34 ( .A(w_CARRY_37_), .Y(_236_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_237_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_238_) );
OAI21X1 OAI21X1_67 ( .A(_236_), .B(_238_), .C(_237_), .Y(w_CARRY_38_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_232_) );
NAND3X1 NAND3X1_34 ( .A(_236_), .B(_237_), .C(_232_), .Y(_233_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_234_) );
OAI21X1 OAI21X1_68 ( .A(_238_), .B(_234_), .C(w_CARRY_37_), .Y(_235_) );
NAND2X1 NAND2X1_68 ( .A(_235_), .B(_233_), .Y(_0__37_) );
INVX1 INVX1_35 ( .A(w_CARRY_38_), .Y(_243_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_244_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_245_) );
OAI21X1 OAI21X1_69 ( .A(_243_), .B(_245_), .C(_244_), .Y(w_CARRY_39_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_239_) );
NAND3X1 NAND3X1_35 ( .A(_243_), .B(_244_), .C(_239_), .Y(_240_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_241_) );
OAI21X1 OAI21X1_70 ( .A(_245_), .B(_241_), .C(w_CARRY_38_), .Y(_242_) );
NAND2X1 NAND2X1_70 ( .A(_242_), .B(_240_), .Y(_0__38_) );
INVX1 INVX1_36 ( .A(w_CARRY_39_), .Y(_250_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_251_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_252_) );
OAI21X1 OAI21X1_71 ( .A(_250_), .B(_252_), .C(_251_), .Y(w_CARRY_40_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_246_) );
NAND3X1 NAND3X1_36 ( .A(_250_), .B(_251_), .C(_246_), .Y(_247_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_248_) );
OAI21X1 OAI21X1_72 ( .A(_252_), .B(_248_), .C(w_CARRY_39_), .Y(_249_) );
NAND2X1 NAND2X1_72 ( .A(_249_), .B(_247_), .Y(_0__39_) );
INVX1 INVX1_37 ( .A(w_CARRY_40_), .Y(_257_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_258_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_259_) );
OAI21X1 OAI21X1_73 ( .A(_257_), .B(_259_), .C(_258_), .Y(w_CARRY_41_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_253_) );
NAND3X1 NAND3X1_37 ( .A(_257_), .B(_258_), .C(_253_), .Y(_254_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_255_) );
OAI21X1 OAI21X1_74 ( .A(_259_), .B(_255_), .C(w_CARRY_40_), .Y(_256_) );
NAND2X1 NAND2X1_74 ( .A(_256_), .B(_254_), .Y(_0__40_) );
INVX1 INVX1_38 ( .A(1'b0), .Y(_264_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_265_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_266_) );
OAI21X1 OAI21X1_75 ( .A(_264_), .B(_266_), .C(_265_), .Y(w_CARRY_1_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_260_) );
NAND3X1 NAND3X1_38 ( .A(_264_), .B(_265_), .C(_260_), .Y(_261_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_262_) );
OAI21X1 OAI21X1_76 ( .A(_266_), .B(_262_), .C(1'b0), .Y(_263_) );
NAND2X1 NAND2X1_76 ( .A(_263_), .B(_261_), .Y(_0__0_) );
INVX1 INVX1_39 ( .A(w_CARRY_1_), .Y(_271_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_272_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_273_) );
OAI21X1 OAI21X1_77 ( .A(_271_), .B(_273_), .C(_272_), .Y(w_CARRY_2_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_267_) );
NAND3X1 NAND3X1_39 ( .A(_271_), .B(_272_), .C(_267_), .Y(_268_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_269_) );
OAI21X1 OAI21X1_78 ( .A(_273_), .B(_269_), .C(w_CARRY_1_), .Y(_270_) );
NAND2X1 NAND2X1_78 ( .A(_270_), .B(_268_), .Y(_0__1_) );
INVX1 INVX1_40 ( .A(w_CARRY_2_), .Y(_278_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_279_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_280_) );
OAI21X1 OAI21X1_79 ( .A(_278_), .B(_280_), .C(_279_), .Y(w_CARRY_3_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_274_) );
NAND3X1 NAND3X1_40 ( .A(_278_), .B(_279_), .C(_274_), .Y(_275_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_276_) );
OAI21X1 OAI21X1_80 ( .A(_280_), .B(_276_), .C(w_CARRY_2_), .Y(_277_) );
NAND2X1 NAND2X1_80 ( .A(_277_), .B(_275_), .Y(_0__2_) );
INVX1 INVX1_41 ( .A(w_CARRY_3_), .Y(_285_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_286_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_287_) );
OAI21X1 OAI21X1_81 ( .A(_285_), .B(_287_), .C(_286_), .Y(w_CARRY_4_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_281_) );
NAND3X1 NAND3X1_41 ( .A(_285_), .B(_286_), .C(_281_), .Y(_282_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_283_) );
OAI21X1 OAI21X1_82 ( .A(_287_), .B(_283_), .C(w_CARRY_3_), .Y(_284_) );
NAND2X1 NAND2X1_82 ( .A(_284_), .B(_282_), .Y(_0__3_) );
BUFX2 BUFX2_43 ( .A(w_CARRY_41_), .Y(_0__41_) );
BUFX2 BUFX2_44 ( .A(1'b0), .Y(w_CARRY_0_) );
endmodule
