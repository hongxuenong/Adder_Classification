module CSkipA_39bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [38:0] i_add_term1;
input [38:0] i_add_term2;
output [38:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

OR2X2 OR2X2_1 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_442_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_443_) );
NAND3X1 NAND3X1_1 ( .A(_441_), .B(_443_), .C(_442_), .Y(_444_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_438_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_439_) );
OAI21X1 OAI21X1_1 ( .A(_438_), .B(_439_), .C(cskip3_inst_rca0_w_CARRY_2_), .Y(_440_) );
NAND2X1 NAND2X1_2 ( .A(_440_), .B(_444_), .Y(_0__38_) );
OAI21X1 OAI21X1_2 ( .A(_441_), .B(_438_), .C(_443_), .Y(cskip3_inst_rca0_w_CARRY_3_) );
INVX1 INVX1_1 ( .A(cskip3_inst_rca0_w_CARRY_3_), .Y(_446_) );
NAND2X1 NAND2X1_3 ( .A(gnd), .B(gnd), .Y(_447_) );
NOR2X1 NOR2X1_2 ( .A(gnd), .B(gnd), .Y(_445_) );
OAI21X1 OAI21X1_3 ( .A(_446_), .B(_445_), .C(_447_), .Y(cskip3_inst_cout0) );
OR2X2 OR2X2_2 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_451_) );
NAND2X1 NAND2X1_4 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_452_) );
NAND2X1 NAND2X1_5 ( .A(_452_), .B(_451_), .Y(_448_) );
XNOR2X1 XNOR2X1_1 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_449_) );
XNOR2X1 XNOR2X1_2 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_450_) );
NOR3X1 NOR3X1_1 ( .A(_448_), .B(_449_), .C(_450_), .Y(cskip3_inst_skip0_P) );
INVX1 INVX1_2 ( .A(cskip3_inst_cout0), .Y(_453_) );
NAND2X1 NAND2X1_6 ( .A(gnd), .B(cskip3_inst_skip0_P), .Y(_454_) );
OAI21X1 OAI21X1_4 ( .A(cskip3_inst_skip0_P), .B(_453_), .C(_454_), .Y(w_cout_10_) );
BUFX2 BUFX2_1 ( .A(w_cout_10_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
INVX1 INVX1_3 ( .A(i_add_term1[0]), .Y(_28_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[0]), .B(_28_), .Y(_29_) );
INVX1 INVX1_4 ( .A(i_add_term2[0]), .Y(_30_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term1[0]), .B(_30_), .Y(_31_) );
INVX1 INVX1_5 ( .A(i_add_term1[1]), .Y(_32_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[1]), .B(_32_), .Y(_33_) );
INVX1 INVX1_6 ( .A(i_add_term2[1]), .Y(_34_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term1[1]), .B(_34_), .Y(_35_) );
OAI22X1 OAI22X1_1 ( .A(_29_), .B(_31_), .C(_33_), .D(_35_), .Y(_36_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_37_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_38_) );
NOR2X1 NOR2X1_8 ( .A(_37_), .B(_38_), .Y(_39_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_40_) );
NAND2X1 NAND2X1_7 ( .A(_39_), .B(_40_), .Y(_41_) );
NOR2X1 NOR2X1_9 ( .A(_36_), .B(_41_), .Y(_3_) );
INVX1 INVX1_7 ( .A(_1_), .Y(_42_) );
NAND2X1 NAND2X1_8 ( .A(gnd), .B(_3_), .Y(_43_) );
OAI21X1 OAI21X1_5 ( .A(_3_), .B(_42_), .C(_43_), .Y(w_cout_1_) );
INVX1 INVX1_8 ( .A(i_add_term1[4]), .Y(_44_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[4]), .B(_44_), .Y(_45_) );
INVX1 INVX1_9 ( .A(i_add_term2[4]), .Y(_46_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term1[4]), .B(_46_), .Y(_47_) );
INVX1 INVX1_10 ( .A(i_add_term1[5]), .Y(_48_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[5]), .B(_48_), .Y(_49_) );
INVX1 INVX1_11 ( .A(i_add_term2[5]), .Y(_50_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term1[5]), .B(_50_), .Y(_51_) );
OAI22X1 OAI22X1_2 ( .A(_45_), .B(_47_), .C(_49_), .D(_51_), .Y(_52_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_53_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_54_) );
NOR2X1 NOR2X1_15 ( .A(_53_), .B(_54_), .Y(_55_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_56_) );
NAND2X1 NAND2X1_9 ( .A(_55_), .B(_56_), .Y(_57_) );
NOR2X1 NOR2X1_16 ( .A(_52_), .B(_57_), .Y(_6_) );
INVX1 INVX1_12 ( .A(_4_), .Y(_58_) );
NAND2X1 NAND2X1_10 ( .A(gnd), .B(_6_), .Y(_59_) );
OAI21X1 OAI21X1_6 ( .A(_6_), .B(_58_), .C(_59_), .Y(w_cout_2_) );
INVX1 INVX1_13 ( .A(i_add_term1[8]), .Y(_60_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[8]), .B(_60_), .Y(_61_) );
INVX1 INVX1_14 ( .A(i_add_term2[8]), .Y(_62_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term1[8]), .B(_62_), .Y(_63_) );
INVX1 INVX1_15 ( .A(i_add_term1[9]), .Y(_64_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[9]), .B(_64_), .Y(_65_) );
INVX1 INVX1_16 ( .A(i_add_term2[9]), .Y(_66_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term1[9]), .B(_66_), .Y(_67_) );
OAI22X1 OAI22X1_3 ( .A(_61_), .B(_63_), .C(_65_), .D(_67_), .Y(_68_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_69_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_70_) );
NOR2X1 NOR2X1_22 ( .A(_69_), .B(_70_), .Y(_71_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_72_) );
NAND2X1 NAND2X1_11 ( .A(_71_), .B(_72_), .Y(_73_) );
NOR2X1 NOR2X1_23 ( .A(_68_), .B(_73_), .Y(_9_) );
INVX1 INVX1_17 ( .A(_7_), .Y(_74_) );
NAND2X1 NAND2X1_12 ( .A(gnd), .B(_9_), .Y(_75_) );
OAI21X1 OAI21X1_7 ( .A(_9_), .B(_74_), .C(_75_), .Y(w_cout_3_) );
INVX1 INVX1_18 ( .A(i_add_term1[12]), .Y(_76_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[12]), .B(_76_), .Y(_77_) );
INVX1 INVX1_19 ( .A(i_add_term2[12]), .Y(_78_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term1[12]), .B(_78_), .Y(_79_) );
INVX1 INVX1_20 ( .A(i_add_term1[13]), .Y(_80_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[13]), .B(_80_), .Y(_81_) );
INVX1 INVX1_21 ( .A(i_add_term2[13]), .Y(_82_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term1[13]), .B(_82_), .Y(_83_) );
OAI22X1 OAI22X1_4 ( .A(_77_), .B(_79_), .C(_81_), .D(_83_), .Y(_84_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_85_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_86_) );
NOR2X1 NOR2X1_29 ( .A(_85_), .B(_86_), .Y(_87_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_88_) );
NAND2X1 NAND2X1_13 ( .A(_87_), .B(_88_), .Y(_89_) );
NOR2X1 NOR2X1_30 ( .A(_84_), .B(_89_), .Y(_12_) );
INVX1 INVX1_22 ( .A(_10_), .Y(_90_) );
NAND2X1 NAND2X1_14 ( .A(gnd), .B(_12_), .Y(_91_) );
OAI21X1 OAI21X1_8 ( .A(_12_), .B(_90_), .C(_91_), .Y(w_cout_4_) );
INVX1 INVX1_23 ( .A(i_add_term1[16]), .Y(_92_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[16]), .B(_92_), .Y(_93_) );
INVX1 INVX1_24 ( .A(i_add_term2[16]), .Y(_94_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term1[16]), .B(_94_), .Y(_95_) );
INVX1 INVX1_25 ( .A(i_add_term1[17]), .Y(_96_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[17]), .B(_96_), .Y(_97_) );
INVX1 INVX1_26 ( .A(i_add_term2[17]), .Y(_98_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term1[17]), .B(_98_), .Y(_99_) );
OAI22X1 OAI22X1_5 ( .A(_93_), .B(_95_), .C(_97_), .D(_99_), .Y(_100_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_101_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_102_) );
NOR2X1 NOR2X1_36 ( .A(_101_), .B(_102_), .Y(_103_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_104_) );
NAND2X1 NAND2X1_15 ( .A(_103_), .B(_104_), .Y(_105_) );
NOR2X1 NOR2X1_37 ( .A(_100_), .B(_105_), .Y(_15_) );
INVX1 INVX1_27 ( .A(_13_), .Y(_106_) );
NAND2X1 NAND2X1_16 ( .A(gnd), .B(_15_), .Y(_107_) );
OAI21X1 OAI21X1_9 ( .A(_15_), .B(_106_), .C(_107_), .Y(w_cout_5_) );
INVX1 INVX1_28 ( .A(i_add_term1[20]), .Y(_108_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[20]), .B(_108_), .Y(_109_) );
INVX1 INVX1_29 ( .A(i_add_term2[20]), .Y(_110_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term1[20]), .B(_110_), .Y(_111_) );
INVX1 INVX1_30 ( .A(i_add_term1[21]), .Y(_112_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[21]), .B(_112_), .Y(_113_) );
INVX1 INVX1_31 ( .A(i_add_term2[21]), .Y(_114_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term1[21]), .B(_114_), .Y(_115_) );
OAI22X1 OAI22X1_6 ( .A(_109_), .B(_111_), .C(_113_), .D(_115_), .Y(_116_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_117_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_118_) );
NOR2X1 NOR2X1_43 ( .A(_117_), .B(_118_), .Y(_119_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_120_) );
NAND2X1 NAND2X1_17 ( .A(_119_), .B(_120_), .Y(_121_) );
NOR2X1 NOR2X1_44 ( .A(_116_), .B(_121_), .Y(_18_) );
INVX1 INVX1_32 ( .A(_16_), .Y(_122_) );
NAND2X1 NAND2X1_18 ( .A(gnd), .B(_18_), .Y(_123_) );
OAI21X1 OAI21X1_10 ( .A(_18_), .B(_122_), .C(_123_), .Y(w_cout_6_) );
INVX1 INVX1_33 ( .A(i_add_term1[24]), .Y(_124_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[24]), .B(_124_), .Y(_125_) );
INVX1 INVX1_34 ( .A(i_add_term2[24]), .Y(_126_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term1[24]), .B(_126_), .Y(_127_) );
INVX1 INVX1_35 ( .A(i_add_term1[25]), .Y(_128_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[25]), .B(_128_), .Y(_129_) );
INVX1 INVX1_36 ( .A(i_add_term2[25]), .Y(_130_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term1[25]), .B(_130_), .Y(_131_) );
OAI22X1 OAI22X1_7 ( .A(_125_), .B(_127_), .C(_129_), .D(_131_), .Y(_132_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_133_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_134_) );
NOR2X1 NOR2X1_50 ( .A(_133_), .B(_134_), .Y(_135_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_136_) );
NAND2X1 NAND2X1_19 ( .A(_135_), .B(_136_), .Y(_137_) );
NOR2X1 NOR2X1_51 ( .A(_132_), .B(_137_), .Y(_21_) );
INVX1 INVX1_37 ( .A(_19_), .Y(_138_) );
NAND2X1 NAND2X1_20 ( .A(gnd), .B(_21_), .Y(_139_) );
OAI21X1 OAI21X1_11 ( .A(_21_), .B(_138_), .C(_139_), .Y(w_cout_7_) );
INVX1 INVX1_38 ( .A(i_add_term1[28]), .Y(_140_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[28]), .B(_140_), .Y(_141_) );
INVX1 INVX1_39 ( .A(i_add_term2[28]), .Y(_142_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term1[28]), .B(_142_), .Y(_143_) );
INVX1 INVX1_40 ( .A(i_add_term1[29]), .Y(_144_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[29]), .B(_144_), .Y(_145_) );
INVX1 INVX1_41 ( .A(i_add_term2[29]), .Y(_146_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term1[29]), .B(_146_), .Y(_147_) );
OAI22X1 OAI22X1_8 ( .A(_141_), .B(_143_), .C(_145_), .D(_147_), .Y(_148_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_149_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_150_) );
NOR2X1 NOR2X1_57 ( .A(_149_), .B(_150_), .Y(_151_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_152_) );
NAND2X1 NAND2X1_21 ( .A(_151_), .B(_152_), .Y(_153_) );
NOR2X1 NOR2X1_58 ( .A(_148_), .B(_153_), .Y(_24_) );
INVX1 INVX1_42 ( .A(_22_), .Y(_154_) );
NAND2X1 NAND2X1_22 ( .A(gnd), .B(_24_), .Y(_155_) );
OAI21X1 OAI21X1_12 ( .A(_24_), .B(_154_), .C(_155_), .Y(w_cout_8_) );
INVX1 INVX1_43 ( .A(i_add_term1[32]), .Y(_156_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[32]), .B(_156_), .Y(_157_) );
INVX1 INVX1_44 ( .A(i_add_term2[32]), .Y(_158_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term1[32]), .B(_158_), .Y(_159_) );
INVX1 INVX1_45 ( .A(i_add_term1[33]), .Y(_160_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[33]), .B(_160_), .Y(_161_) );
INVX1 INVX1_46 ( .A(i_add_term2[33]), .Y(_162_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term1[33]), .B(_162_), .Y(_163_) );
OAI22X1 OAI22X1_9 ( .A(_157_), .B(_159_), .C(_161_), .D(_163_), .Y(_164_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_165_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_166_) );
NOR2X1 NOR2X1_64 ( .A(_165_), .B(_166_), .Y(_167_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_168_) );
NAND2X1 NAND2X1_23 ( .A(_167_), .B(_168_), .Y(_169_) );
NOR2X1 NOR2X1_65 ( .A(_164_), .B(_169_), .Y(_27_) );
INVX1 INVX1_47 ( .A(_25_), .Y(_170_) );
NAND2X1 NAND2X1_24 ( .A(gnd), .B(_27_), .Y(_171_) );
OAI21X1 OAI21X1_13 ( .A(_27_), .B(_170_), .C(_171_), .Y(cskip3_inst_cin) );
INVX1 INVX1_48 ( .A(gnd), .Y(_175_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_176_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_177_) );
NAND3X1 NAND3X1_2 ( .A(_175_), .B(_177_), .C(_176_), .Y(_178_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_172_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_173_) );
OAI21X1 OAI21X1_14 ( .A(_172_), .B(_173_), .C(gnd), .Y(_174_) );
NAND2X1 NAND2X1_26 ( .A(_174_), .B(_178_), .Y(_0__0_) );
OAI21X1 OAI21X1_15 ( .A(_175_), .B(_172_), .C(_177_), .Y(_2__1_) );
INVX1 INVX1_49 ( .A(_2__1_), .Y(_182_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_183_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_184_) );
NAND3X1 NAND3X1_3 ( .A(_182_), .B(_184_), .C(_183_), .Y(_185_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_179_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_180_) );
OAI21X1 OAI21X1_16 ( .A(_179_), .B(_180_), .C(_2__1_), .Y(_181_) );
NAND2X1 NAND2X1_28 ( .A(_181_), .B(_185_), .Y(_0__1_) );
OAI21X1 OAI21X1_17 ( .A(_182_), .B(_179_), .C(_184_), .Y(_2__2_) );
INVX1 INVX1_50 ( .A(_2__2_), .Y(_189_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_190_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_191_) );
NAND3X1 NAND3X1_4 ( .A(_189_), .B(_191_), .C(_190_), .Y(_192_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_186_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_187_) );
OAI21X1 OAI21X1_18 ( .A(_186_), .B(_187_), .C(_2__2_), .Y(_188_) );
NAND2X1 NAND2X1_30 ( .A(_188_), .B(_192_), .Y(_0__2_) );
OAI21X1 OAI21X1_19 ( .A(_189_), .B(_186_), .C(_191_), .Y(_2__3_) );
INVX1 INVX1_51 ( .A(_2__3_), .Y(_196_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_197_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_198_) );
NAND3X1 NAND3X1_5 ( .A(_196_), .B(_198_), .C(_197_), .Y(_199_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_193_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_194_) );
OAI21X1 OAI21X1_20 ( .A(_193_), .B(_194_), .C(_2__3_), .Y(_195_) );
NAND2X1 NAND2X1_32 ( .A(_195_), .B(_199_), .Y(_0__3_) );
OAI21X1 OAI21X1_21 ( .A(_196_), .B(_193_), .C(_198_), .Y(_1_) );
INVX1 INVX1_52 ( .A(w_cout_1_), .Y(_203_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_204_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_205_) );
NAND3X1 NAND3X1_6 ( .A(_203_), .B(_205_), .C(_204_), .Y(_206_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_200_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_201_) );
OAI21X1 OAI21X1_22 ( .A(_200_), .B(_201_), .C(w_cout_1_), .Y(_202_) );
NAND2X1 NAND2X1_34 ( .A(_202_), .B(_206_), .Y(_0__4_) );
OAI21X1 OAI21X1_23 ( .A(_203_), .B(_200_), .C(_205_), .Y(_5__1_) );
INVX1 INVX1_53 ( .A(_5__1_), .Y(_210_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_211_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_212_) );
NAND3X1 NAND3X1_7 ( .A(_210_), .B(_212_), .C(_211_), .Y(_213_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_207_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_208_) );
OAI21X1 OAI21X1_24 ( .A(_207_), .B(_208_), .C(_5__1_), .Y(_209_) );
NAND2X1 NAND2X1_36 ( .A(_209_), .B(_213_), .Y(_0__5_) );
OAI21X1 OAI21X1_25 ( .A(_210_), .B(_207_), .C(_212_), .Y(_5__2_) );
INVX1 INVX1_54 ( .A(_5__2_), .Y(_217_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_218_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_219_) );
NAND3X1 NAND3X1_8 ( .A(_217_), .B(_219_), .C(_218_), .Y(_220_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_214_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_215_) );
OAI21X1 OAI21X1_26 ( .A(_214_), .B(_215_), .C(_5__2_), .Y(_216_) );
NAND2X1 NAND2X1_38 ( .A(_216_), .B(_220_), .Y(_0__6_) );
OAI21X1 OAI21X1_27 ( .A(_217_), .B(_214_), .C(_219_), .Y(_5__3_) );
INVX1 INVX1_55 ( .A(_5__3_), .Y(_224_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_225_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_226_) );
NAND3X1 NAND3X1_9 ( .A(_224_), .B(_226_), .C(_225_), .Y(_227_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_221_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_222_) );
OAI21X1 OAI21X1_28 ( .A(_221_), .B(_222_), .C(_5__3_), .Y(_223_) );
NAND2X1 NAND2X1_40 ( .A(_223_), .B(_227_), .Y(_0__7_) );
OAI21X1 OAI21X1_29 ( .A(_224_), .B(_221_), .C(_226_), .Y(_4_) );
INVX1 INVX1_56 ( .A(w_cout_2_), .Y(_231_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_232_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_233_) );
NAND3X1 NAND3X1_10 ( .A(_231_), .B(_233_), .C(_232_), .Y(_234_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_228_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_229_) );
OAI21X1 OAI21X1_30 ( .A(_228_), .B(_229_), .C(w_cout_2_), .Y(_230_) );
NAND2X1 NAND2X1_42 ( .A(_230_), .B(_234_), .Y(_0__8_) );
OAI21X1 OAI21X1_31 ( .A(_231_), .B(_228_), .C(_233_), .Y(_8__1_) );
INVX1 INVX1_57 ( .A(_8__1_), .Y(_238_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_239_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_240_) );
NAND3X1 NAND3X1_11 ( .A(_238_), .B(_240_), .C(_239_), .Y(_241_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_235_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_236_) );
OAI21X1 OAI21X1_32 ( .A(_235_), .B(_236_), .C(_8__1_), .Y(_237_) );
NAND2X1 NAND2X1_44 ( .A(_237_), .B(_241_), .Y(_0__9_) );
OAI21X1 OAI21X1_33 ( .A(_238_), .B(_235_), .C(_240_), .Y(_8__2_) );
INVX1 INVX1_58 ( .A(_8__2_), .Y(_245_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_246_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_247_) );
NAND3X1 NAND3X1_12 ( .A(_245_), .B(_247_), .C(_246_), .Y(_248_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_242_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_243_) );
OAI21X1 OAI21X1_34 ( .A(_242_), .B(_243_), .C(_8__2_), .Y(_244_) );
NAND2X1 NAND2X1_46 ( .A(_244_), .B(_248_), .Y(_0__10_) );
OAI21X1 OAI21X1_35 ( .A(_245_), .B(_242_), .C(_247_), .Y(_8__3_) );
INVX1 INVX1_59 ( .A(_8__3_), .Y(_252_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_253_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_254_) );
NAND3X1 NAND3X1_13 ( .A(_252_), .B(_254_), .C(_253_), .Y(_255_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_249_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_250_) );
OAI21X1 OAI21X1_36 ( .A(_249_), .B(_250_), .C(_8__3_), .Y(_251_) );
NAND2X1 NAND2X1_48 ( .A(_251_), .B(_255_), .Y(_0__11_) );
OAI21X1 OAI21X1_37 ( .A(_252_), .B(_249_), .C(_254_), .Y(_7_) );
INVX1 INVX1_60 ( .A(w_cout_3_), .Y(_259_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_260_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_261_) );
NAND3X1 NAND3X1_14 ( .A(_259_), .B(_261_), .C(_260_), .Y(_262_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_256_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_257_) );
OAI21X1 OAI21X1_38 ( .A(_256_), .B(_257_), .C(w_cout_3_), .Y(_258_) );
NAND2X1 NAND2X1_50 ( .A(_258_), .B(_262_), .Y(_0__12_) );
OAI21X1 OAI21X1_39 ( .A(_259_), .B(_256_), .C(_261_), .Y(_11__1_) );
INVX1 INVX1_61 ( .A(_11__1_), .Y(_266_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_267_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_268_) );
NAND3X1 NAND3X1_15 ( .A(_266_), .B(_268_), .C(_267_), .Y(_269_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_263_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_264_) );
OAI21X1 OAI21X1_40 ( .A(_263_), .B(_264_), .C(_11__1_), .Y(_265_) );
NAND2X1 NAND2X1_52 ( .A(_265_), .B(_269_), .Y(_0__13_) );
OAI21X1 OAI21X1_41 ( .A(_266_), .B(_263_), .C(_268_), .Y(_11__2_) );
INVX1 INVX1_62 ( .A(_11__2_), .Y(_273_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_274_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_275_) );
NAND3X1 NAND3X1_16 ( .A(_273_), .B(_275_), .C(_274_), .Y(_276_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_270_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_271_) );
OAI21X1 OAI21X1_42 ( .A(_270_), .B(_271_), .C(_11__2_), .Y(_272_) );
NAND2X1 NAND2X1_54 ( .A(_272_), .B(_276_), .Y(_0__14_) );
OAI21X1 OAI21X1_43 ( .A(_273_), .B(_270_), .C(_275_), .Y(_11__3_) );
INVX1 INVX1_63 ( .A(_11__3_), .Y(_280_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_281_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_282_) );
NAND3X1 NAND3X1_17 ( .A(_280_), .B(_282_), .C(_281_), .Y(_283_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_277_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_278_) );
OAI21X1 OAI21X1_44 ( .A(_277_), .B(_278_), .C(_11__3_), .Y(_279_) );
NAND2X1 NAND2X1_56 ( .A(_279_), .B(_283_), .Y(_0__15_) );
OAI21X1 OAI21X1_45 ( .A(_280_), .B(_277_), .C(_282_), .Y(_10_) );
INVX1 INVX1_64 ( .A(w_cout_4_), .Y(_287_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_288_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_289_) );
NAND3X1 NAND3X1_18 ( .A(_287_), .B(_289_), .C(_288_), .Y(_290_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_284_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_285_) );
OAI21X1 OAI21X1_46 ( .A(_284_), .B(_285_), .C(w_cout_4_), .Y(_286_) );
NAND2X1 NAND2X1_58 ( .A(_286_), .B(_290_), .Y(_0__16_) );
OAI21X1 OAI21X1_47 ( .A(_287_), .B(_284_), .C(_289_), .Y(_14__1_) );
INVX1 INVX1_65 ( .A(_14__1_), .Y(_294_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_295_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_296_) );
NAND3X1 NAND3X1_19 ( .A(_294_), .B(_296_), .C(_295_), .Y(_297_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_291_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_292_) );
OAI21X1 OAI21X1_48 ( .A(_291_), .B(_292_), .C(_14__1_), .Y(_293_) );
NAND2X1 NAND2X1_60 ( .A(_293_), .B(_297_), .Y(_0__17_) );
OAI21X1 OAI21X1_49 ( .A(_294_), .B(_291_), .C(_296_), .Y(_14__2_) );
INVX1 INVX1_66 ( .A(_14__2_), .Y(_301_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_302_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_303_) );
NAND3X1 NAND3X1_20 ( .A(_301_), .B(_303_), .C(_302_), .Y(_304_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_298_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_299_) );
OAI21X1 OAI21X1_50 ( .A(_298_), .B(_299_), .C(_14__2_), .Y(_300_) );
NAND2X1 NAND2X1_62 ( .A(_300_), .B(_304_), .Y(_0__18_) );
OAI21X1 OAI21X1_51 ( .A(_301_), .B(_298_), .C(_303_), .Y(_14__3_) );
INVX1 INVX1_67 ( .A(_14__3_), .Y(_308_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_309_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_310_) );
NAND3X1 NAND3X1_21 ( .A(_308_), .B(_310_), .C(_309_), .Y(_311_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_305_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_306_) );
OAI21X1 OAI21X1_52 ( .A(_305_), .B(_306_), .C(_14__3_), .Y(_307_) );
NAND2X1 NAND2X1_64 ( .A(_307_), .B(_311_), .Y(_0__19_) );
OAI21X1 OAI21X1_53 ( .A(_308_), .B(_305_), .C(_310_), .Y(_13_) );
INVX1 INVX1_68 ( .A(w_cout_5_), .Y(_315_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_316_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_317_) );
NAND3X1 NAND3X1_22 ( .A(_315_), .B(_317_), .C(_316_), .Y(_318_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_312_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_313_) );
OAI21X1 OAI21X1_54 ( .A(_312_), .B(_313_), .C(w_cout_5_), .Y(_314_) );
NAND2X1 NAND2X1_66 ( .A(_314_), .B(_318_), .Y(_0__20_) );
OAI21X1 OAI21X1_55 ( .A(_315_), .B(_312_), .C(_317_), .Y(_17__1_) );
INVX1 INVX1_69 ( .A(_17__1_), .Y(_322_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_323_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_324_) );
NAND3X1 NAND3X1_23 ( .A(_322_), .B(_324_), .C(_323_), .Y(_325_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_319_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_320_) );
OAI21X1 OAI21X1_56 ( .A(_319_), .B(_320_), .C(_17__1_), .Y(_321_) );
NAND2X1 NAND2X1_68 ( .A(_321_), .B(_325_), .Y(_0__21_) );
OAI21X1 OAI21X1_57 ( .A(_322_), .B(_319_), .C(_324_), .Y(_17__2_) );
INVX1 INVX1_70 ( .A(_17__2_), .Y(_329_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_330_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_331_) );
NAND3X1 NAND3X1_24 ( .A(_329_), .B(_331_), .C(_330_), .Y(_332_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_326_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_327_) );
OAI21X1 OAI21X1_58 ( .A(_326_), .B(_327_), .C(_17__2_), .Y(_328_) );
NAND2X1 NAND2X1_70 ( .A(_328_), .B(_332_), .Y(_0__22_) );
OAI21X1 OAI21X1_59 ( .A(_329_), .B(_326_), .C(_331_), .Y(_17__3_) );
INVX1 INVX1_71 ( .A(_17__3_), .Y(_336_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_337_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_338_) );
NAND3X1 NAND3X1_25 ( .A(_336_), .B(_338_), .C(_337_), .Y(_339_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_333_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_334_) );
OAI21X1 OAI21X1_60 ( .A(_333_), .B(_334_), .C(_17__3_), .Y(_335_) );
NAND2X1 NAND2X1_72 ( .A(_335_), .B(_339_), .Y(_0__23_) );
OAI21X1 OAI21X1_61 ( .A(_336_), .B(_333_), .C(_338_), .Y(_16_) );
INVX1 INVX1_72 ( .A(w_cout_6_), .Y(_343_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_344_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_345_) );
NAND3X1 NAND3X1_26 ( .A(_343_), .B(_345_), .C(_344_), .Y(_346_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_340_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_341_) );
OAI21X1 OAI21X1_62 ( .A(_340_), .B(_341_), .C(w_cout_6_), .Y(_342_) );
NAND2X1 NAND2X1_74 ( .A(_342_), .B(_346_), .Y(_0__24_) );
OAI21X1 OAI21X1_63 ( .A(_343_), .B(_340_), .C(_345_), .Y(_20__1_) );
INVX1 INVX1_73 ( .A(_20__1_), .Y(_350_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_351_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_352_) );
NAND3X1 NAND3X1_27 ( .A(_350_), .B(_352_), .C(_351_), .Y(_353_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_347_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_348_) );
OAI21X1 OAI21X1_64 ( .A(_347_), .B(_348_), .C(_20__1_), .Y(_349_) );
NAND2X1 NAND2X1_76 ( .A(_349_), .B(_353_), .Y(_0__25_) );
OAI21X1 OAI21X1_65 ( .A(_350_), .B(_347_), .C(_352_), .Y(_20__2_) );
INVX1 INVX1_74 ( .A(_20__2_), .Y(_357_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_358_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_359_) );
NAND3X1 NAND3X1_28 ( .A(_357_), .B(_359_), .C(_358_), .Y(_360_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_354_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_355_) );
OAI21X1 OAI21X1_66 ( .A(_354_), .B(_355_), .C(_20__2_), .Y(_356_) );
NAND2X1 NAND2X1_78 ( .A(_356_), .B(_360_), .Y(_0__26_) );
OAI21X1 OAI21X1_67 ( .A(_357_), .B(_354_), .C(_359_), .Y(_20__3_) );
INVX1 INVX1_75 ( .A(_20__3_), .Y(_364_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_365_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_366_) );
NAND3X1 NAND3X1_29 ( .A(_364_), .B(_366_), .C(_365_), .Y(_367_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_361_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_362_) );
OAI21X1 OAI21X1_68 ( .A(_361_), .B(_362_), .C(_20__3_), .Y(_363_) );
NAND2X1 NAND2X1_80 ( .A(_363_), .B(_367_), .Y(_0__27_) );
OAI21X1 OAI21X1_69 ( .A(_364_), .B(_361_), .C(_366_), .Y(_19_) );
INVX1 INVX1_76 ( .A(w_cout_7_), .Y(_371_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_372_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_373_) );
NAND3X1 NAND3X1_30 ( .A(_371_), .B(_373_), .C(_372_), .Y(_374_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_368_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_369_) );
OAI21X1 OAI21X1_70 ( .A(_368_), .B(_369_), .C(w_cout_7_), .Y(_370_) );
NAND2X1 NAND2X1_82 ( .A(_370_), .B(_374_), .Y(_0__28_) );
OAI21X1 OAI21X1_71 ( .A(_371_), .B(_368_), .C(_373_), .Y(_23__1_) );
INVX1 INVX1_77 ( .A(_23__1_), .Y(_378_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_379_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_380_) );
NAND3X1 NAND3X1_31 ( .A(_378_), .B(_380_), .C(_379_), .Y(_381_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_375_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_376_) );
OAI21X1 OAI21X1_72 ( .A(_375_), .B(_376_), .C(_23__1_), .Y(_377_) );
NAND2X1 NAND2X1_84 ( .A(_377_), .B(_381_), .Y(_0__29_) );
OAI21X1 OAI21X1_73 ( .A(_378_), .B(_375_), .C(_380_), .Y(_23__2_) );
INVX1 INVX1_78 ( .A(_23__2_), .Y(_385_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_386_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_387_) );
NAND3X1 NAND3X1_32 ( .A(_385_), .B(_387_), .C(_386_), .Y(_388_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_382_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_383_) );
OAI21X1 OAI21X1_74 ( .A(_382_), .B(_383_), .C(_23__2_), .Y(_384_) );
NAND2X1 NAND2X1_86 ( .A(_384_), .B(_388_), .Y(_0__30_) );
OAI21X1 OAI21X1_75 ( .A(_385_), .B(_382_), .C(_387_), .Y(_23__3_) );
INVX1 INVX1_79 ( .A(_23__3_), .Y(_392_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_393_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_394_) );
NAND3X1 NAND3X1_33 ( .A(_392_), .B(_394_), .C(_393_), .Y(_395_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_389_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_390_) );
OAI21X1 OAI21X1_76 ( .A(_389_), .B(_390_), .C(_23__3_), .Y(_391_) );
NAND2X1 NAND2X1_88 ( .A(_391_), .B(_395_), .Y(_0__31_) );
OAI21X1 OAI21X1_77 ( .A(_392_), .B(_389_), .C(_394_), .Y(_22_) );
INVX1 INVX1_80 ( .A(w_cout_8_), .Y(_399_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_400_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_401_) );
NAND3X1 NAND3X1_34 ( .A(_399_), .B(_401_), .C(_400_), .Y(_402_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_396_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_397_) );
OAI21X1 OAI21X1_78 ( .A(_396_), .B(_397_), .C(w_cout_8_), .Y(_398_) );
NAND2X1 NAND2X1_90 ( .A(_398_), .B(_402_), .Y(_0__32_) );
OAI21X1 OAI21X1_79 ( .A(_399_), .B(_396_), .C(_401_), .Y(_26__1_) );
INVX1 INVX1_81 ( .A(_26__1_), .Y(_406_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_407_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_408_) );
NAND3X1 NAND3X1_35 ( .A(_406_), .B(_408_), .C(_407_), .Y(_409_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_403_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_404_) );
OAI21X1 OAI21X1_80 ( .A(_403_), .B(_404_), .C(_26__1_), .Y(_405_) );
NAND2X1 NAND2X1_92 ( .A(_405_), .B(_409_), .Y(_0__33_) );
OAI21X1 OAI21X1_81 ( .A(_406_), .B(_403_), .C(_408_), .Y(_26__2_) );
INVX1 INVX1_82 ( .A(_26__2_), .Y(_413_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_414_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_415_) );
NAND3X1 NAND3X1_36 ( .A(_413_), .B(_415_), .C(_414_), .Y(_416_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_410_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_411_) );
OAI21X1 OAI21X1_82 ( .A(_410_), .B(_411_), .C(_26__2_), .Y(_412_) );
NAND2X1 NAND2X1_94 ( .A(_412_), .B(_416_), .Y(_0__34_) );
OAI21X1 OAI21X1_83 ( .A(_413_), .B(_410_), .C(_415_), .Y(_26__3_) );
INVX1 INVX1_83 ( .A(_26__3_), .Y(_420_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_421_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_422_) );
NAND3X1 NAND3X1_37 ( .A(_420_), .B(_422_), .C(_421_), .Y(_423_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_417_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_418_) );
OAI21X1 OAI21X1_84 ( .A(_417_), .B(_418_), .C(_26__3_), .Y(_419_) );
NAND2X1 NAND2X1_96 ( .A(_419_), .B(_423_), .Y(_0__35_) );
OAI21X1 OAI21X1_85 ( .A(_420_), .B(_417_), .C(_422_), .Y(_25_) );
INVX1 INVX1_84 ( .A(cskip3_inst_cin), .Y(_427_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_428_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_429_) );
NAND3X1 NAND3X1_38 ( .A(_427_), .B(_429_), .C(_428_), .Y(_430_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_424_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_425_) );
OAI21X1 OAI21X1_86 ( .A(_424_), .B(_425_), .C(cskip3_inst_cin), .Y(_426_) );
NAND2X1 NAND2X1_98 ( .A(_426_), .B(_430_), .Y(_0__36_) );
OAI21X1 OAI21X1_87 ( .A(_427_), .B(_424_), .C(_429_), .Y(cskip3_inst_rca0_w_CARRY_1_) );
INVX1 INVX1_85 ( .A(cskip3_inst_rca0_w_CARRY_1_), .Y(_434_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_435_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_436_) );
NAND3X1 NAND3X1_39 ( .A(_434_), .B(_436_), .C(_435_), .Y(_437_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_431_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_432_) );
OAI21X1 OAI21X1_88 ( .A(_431_), .B(_432_), .C(cskip3_inst_rca0_w_CARRY_1_), .Y(_433_) );
NAND2X1 NAND2X1_100 ( .A(_433_), .B(_437_), .Y(_0__37_) );
OAI21X1 OAI21X1_89 ( .A(_434_), .B(_431_), .C(_436_), .Y(cskip3_inst_rca0_w_CARRY_2_) );
INVX1 INVX1_86 ( .A(cskip3_inst_rca0_w_CARRY_2_), .Y(_441_) );
BUFX2 BUFX2_41 ( .A(gnd), .Y(_2__0_) );
BUFX2 BUFX2_42 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_43 ( .A(w_cout_1_), .Y(_5__0_) );
BUFX2 BUFX2_44 ( .A(_4_), .Y(_5__4_) );
BUFX2 BUFX2_45 ( .A(w_cout_2_), .Y(_8__0_) );
BUFX2 BUFX2_46 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_47 ( .A(w_cout_3_), .Y(_11__0_) );
BUFX2 BUFX2_48 ( .A(_10_), .Y(_11__4_) );
BUFX2 BUFX2_49 ( .A(w_cout_4_), .Y(_14__0_) );
BUFX2 BUFX2_50 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_51 ( .A(w_cout_5_), .Y(_17__0_) );
BUFX2 BUFX2_52 ( .A(_16_), .Y(_17__4_) );
BUFX2 BUFX2_53 ( .A(w_cout_6_), .Y(_20__0_) );
BUFX2 BUFX2_54 ( .A(_19_), .Y(_20__4_) );
BUFX2 BUFX2_55 ( .A(w_cout_7_), .Y(_23__0_) );
BUFX2 BUFX2_56 ( .A(_22_), .Y(_23__4_) );
BUFX2 BUFX2_57 ( .A(w_cout_8_), .Y(_26__0_) );
BUFX2 BUFX2_58 ( .A(_25_), .Y(_26__4_) );
BUFX2 BUFX2_59 ( .A(cskip3_inst_cin), .Y(cskip3_inst_rca0_w_CARRY_0_) );
BUFX2 BUFX2_60 ( .A(cskip3_inst_cout0), .Y(cskip3_inst_rca0_w_CARRY_4_) );
BUFX2 BUFX2_61 ( .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_62 ( .A(cskip3_inst_cin), .Y(w_cout_9_) );
endmodule
