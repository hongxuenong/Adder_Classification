module cla_45bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [44:0] i_add1;
input [44:0] i_add2;
output [45:0] o_result;

OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_325_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_326_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_326_), .C(_325_), .Y(_327_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_321_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_322_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_322_), .C(w_C_12_), .Y(_323_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_327_), .Y(_264__12_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(w_C_13_), .Y(_331_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_332_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_333_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_333_), .C(_332_), .Y(_334_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_328_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_329_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_329_), .C(w_C_13_), .Y(_330_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_334_), .Y(_264__13_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(w_C_14_), .Y(_338_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_339_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_340_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_340_), .C(_339_), .Y(_341_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_335_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_336_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_335_), .B(_336_), .C(w_C_14_), .Y(_337_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_341_), .Y(_264__14_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(_345_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_346_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_347_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_347_), .C(_346_), .Y(_348_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_342_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_343_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_343_), .C(w_C_15_), .Y(_344_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_348_), .Y(_264__15_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(w_C_16_), .Y(_352_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_353_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_354_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_354_), .C(_353_), .Y(_355_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_349_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_350_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_350_), .C(w_C_16_), .Y(_351_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_355_), .Y(_264__16_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(w_C_17_), .Y(_359_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_360_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_361_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_361_), .C(_360_), .Y(_362_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_356_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_357_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_357_), .C(w_C_17_), .Y(_358_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_358_), .B(_362_), .Y(_264__17_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(w_C_18_), .Y(_366_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_367_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_368_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_368_), .C(_367_), .Y(_369_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_363_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_364_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_364_), .C(w_C_18_), .Y(_365_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_365_), .B(_369_), .Y(_264__18_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(w_C_19_), .Y(_373_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_374_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_375_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_373_), .B(_375_), .C(_374_), .Y(_376_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_370_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_371_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_371_), .C(w_C_19_), .Y(_372_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_376_), .Y(_264__19_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(w_C_20_), .Y(_380_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_381_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_382_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_382_), .C(_381_), .Y(_383_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_377_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_378_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_378_), .C(w_C_20_), .Y(_379_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_383_), .Y(_264__20_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(w_C_21_), .Y(_387_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_388_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_389_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_389_), .C(_388_), .Y(_390_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_384_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_385_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_385_), .C(w_C_21_), .Y(_386_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_390_), .Y(_264__21_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(w_C_22_), .Y(_394_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_395_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_396_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_396_), .C(_395_), .Y(_397_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_391_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_392_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_392_), .C(w_C_22_), .Y(_393_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_397_), .Y(_264__22_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(w_C_23_), .Y(_401_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_402_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_403_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_403_), .C(_402_), .Y(_404_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_398_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_399_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_399_), .C(w_C_23_), .Y(_400_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_400_), .B(_404_), .Y(_264__23_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(w_C_24_), .Y(_408_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_409_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_410_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_410_), .C(_409_), .Y(_411_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_405_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_406_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_406_), .C(w_C_24_), .Y(_407_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_411_), .Y(_264__24_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(w_C_25_), .Y(_415_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_416_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_417_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_415_), .B(_417_), .C(_416_), .Y(_418_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_412_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_413_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_413_), .C(w_C_25_), .Y(_414_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_414_), .B(_418_), .Y(_264__25_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(w_C_26_), .Y(_422_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_423_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_424_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_422_), .B(_424_), .C(_423_), .Y(_425_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_419_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_420_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_420_), .C(w_C_26_), .Y(_421_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_425_), .Y(_264__26_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(w_C_27_), .Y(_429_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_430_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_431_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(_431_), .C(_430_), .Y(_432_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_426_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_427_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_427_), .C(w_C_27_), .Y(_428_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_432_), .Y(_264__27_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(w_C_28_), .Y(_436_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_437_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_438_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_438_), .C(_437_), .Y(_439_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_433_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_434_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_434_), .C(w_C_28_), .Y(_435_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_439_), .Y(_264__28_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(w_C_29_), .Y(_443_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_444_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_445_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_445_), .C(_444_), .Y(_446_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_440_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_441_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_441_), .C(w_C_29_), .Y(_442_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_446_), .Y(_264__29_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(w_C_30_), .Y(_450_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_451_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_452_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_452_), .C(_451_), .Y(_453_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_447_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_448_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_448_), .C(w_C_30_), .Y(_449_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_453_), .Y(_264__30_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(w_C_31_), .Y(_457_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_458_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_459_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_459_), .C(_458_), .Y(_460_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_454_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_455_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_454_), .B(_455_), .C(w_C_31_), .Y(_456_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_456_), .B(_460_), .Y(_264__31_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(w_C_32_), .Y(_464_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_465_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_466_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_466_), .C(_465_), .Y(_467_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_461_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_462_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_462_), .C(w_C_32_), .Y(_463_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_467_), .Y(_264__32_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(w_C_33_), .Y(_471_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_472_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_473_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_473_), .C(_472_), .Y(_474_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_468_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_469_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_468_), .B(_469_), .C(w_C_33_), .Y(_470_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_470_), .B(_474_), .Y(_264__33_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(w_C_34_), .Y(_478_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_479_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_480_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_480_), .C(_479_), .Y(_481_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_475_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_476_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_476_), .C(w_C_34_), .Y(_477_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_477_), .B(_481_), .Y(_264__34_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(w_C_35_), .Y(_485_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_486_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_487_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_487_), .C(_486_), .Y(_488_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_482_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_483_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_482_), .B(_483_), .C(w_C_35_), .Y(_484_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_484_), .B(_488_), .Y(_264__35_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(w_C_36_), .Y(_492_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_493_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_494_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_492_), .B(_494_), .C(_493_), .Y(_495_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_489_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_490_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_490_), .C(w_C_36_), .Y(_491_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_495_), .Y(_264__36_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(w_C_37_), .Y(_499_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_500_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_501_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_501_), .C(_500_), .Y(_502_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_496_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_497_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_497_), .C(w_C_37_), .Y(_498_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_502_), .Y(_264__37_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(w_C_38_), .Y(_506_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_507_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_508_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_508_), .C(_507_), .Y(_509_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_503_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_504_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_504_), .C(w_C_38_), .Y(_505_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(_509_), .Y(_264__38_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(w_C_39_), .Y(_513_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_514_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_515_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_515_), .C(_514_), .Y(_516_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_510_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_511_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_511_), .C(w_C_39_), .Y(_512_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_516_), .Y(_264__39_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(w_C_40_), .Y(_520_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_521_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_522_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_522_), .C(_521_), .Y(_523_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_517_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_518_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_517_), .B(_518_), .C(w_C_40_), .Y(_519_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_523_), .Y(_264__40_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(w_C_41_), .Y(_527_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_528_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_529_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_529_), .C(_528_), .Y(_530_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_524_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_525_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_525_), .C(w_C_41_), .Y(_526_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_530_), .Y(_264__41_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(w_C_42_), .Y(_534_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_535_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_536_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_536_), .C(_535_), .Y(_537_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_531_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_532_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_532_), .C(w_C_42_), .Y(_533_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_537_), .Y(_264__42_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(w_C_43_), .Y(_541_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_542_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_543_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_541_), .B(_543_), .C(_542_), .Y(_544_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_538_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_539_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_539_), .C(w_C_43_), .Y(_540_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_544_), .Y(_264__43_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(w_C_44_), .Y(_548_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_549_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_550_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_550_), .C(_549_), .Y(_551_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_545_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_546_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_546_), .C(w_C_44_), .Y(_547_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_551_), .Y(_264__44_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_555_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_556_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_557_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_555_), .B(_557_), .C(_556_), .Y(_558_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_552_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_553_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_552_), .B(_553_), .C(gnd), .Y(_554_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_558_), .Y(_264__0_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_562_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_563_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_564_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_562_), .B(_564_), .C(_563_), .Y(_565_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_559_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_560_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_560_), .C(w_C_1_), .Y(_561_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_565_), .Y(_264__1_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_569_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_570_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_571_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_569_), .B(_571_), .C(_570_), .Y(_572_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_566_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_567_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_567_), .C(w_C_2_), .Y(_568_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_572_), .Y(_264__2_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_576_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_577_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_578_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_576_), .B(_578_), .C(_577_), .Y(_579_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_573_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_574_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_574_), .C(w_C_3_), .Y(_575_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_579_), .Y(_264__3_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_253_), .C(_252_), .Y(_254_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_244_), .C(_254_), .Y(_255_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_256_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_256_), .C(_255_), .Y(_257_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_257_), .Y(w_C_43_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_258_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_259_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_259_), .C(_257_), .Y(_260_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_258_), .Y(w_C_44_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_261_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_262_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_262_), .C(_260_), .Y(_263_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_263_), .Y(w_C_45_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_7_), .Y(w_C_3_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .Y(_8_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add1[3]), .Y(_9_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_9_), .Y(_10_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_11_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_11_), .C(_7_), .Y(_12_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_10_), .Y(w_C_4_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_14_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_14_), .C(_12_), .Y(_15_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_15_), .Y(w_C_5_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_16_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_17_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_18_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_18_), .C(_15_), .Y(_19_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_17_), .Y(w_C_6_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .Y(_20_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add1[6]), .Y(_21_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_23_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_23_), .C(_19_), .Y(_24_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .C(_24_), .Y(w_C_7_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .Y(_25_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(_26_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_27_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(_28_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_28_), .C(_24_), .Y(_29_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .C(_29_), .Y(_30_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(w_C_8_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .Y(_31_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add1[8]), .Y(_32_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_33_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_33_), .Y(_34_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_35_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_35_), .Y(_36_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_36_), .C(_29_), .Y(_37_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_32_), .C(_37_), .Y(w_C_9_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_32_), .Y(_38_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_38_), .Y(_39_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_40_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_40_), .Y(_41_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_41_), .C(_37_), .Y(_42_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .C(_42_), .Y(_43_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(w_C_10_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .Y(_44_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add1[10]), .Y(_45_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_46_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_46_), .Y(_47_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_48_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_48_), .Y(_49_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_49_), .C(_42_), .Y(_50_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_45_), .C(_50_), .Y(w_C_11_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_45_), .Y(_51_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_51_), .Y(_52_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_53_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_53_), .Y(_54_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_54_), .C(_50_), .Y(_55_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .C(_55_), .Y(_56_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_56_), .Y(w_C_12_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .Y(_57_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add1[12]), .Y(_58_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_59_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_59_), .Y(_60_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_61_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_61_), .Y(_62_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_62_), .C(_55_), .Y(_63_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_58_), .C(_63_), .Y(w_C_13_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_58_), .Y(_64_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_64_), .Y(_65_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_66_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_66_), .Y(_67_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_67_), .C(_63_), .Y(_68_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .C(_68_), .Y(_69_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(w_C_14_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .Y(_70_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add1[14]), .Y(_71_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_72_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(_72_), .Y(_73_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_74_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_74_), .Y(_75_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_75_), .C(_68_), .Y(_76_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_71_), .C(_76_), .Y(w_C_15_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_71_), .Y(_77_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(_78_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_79_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_79_), .Y(_80_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_80_), .C(_76_), .Y(_81_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .C(_81_), .Y(_82_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_82_), .Y(w_C_16_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .Y(_83_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add1[16]), .Y(_84_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_84_), .Y(_85_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_85_), .Y(_86_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_87_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(_87_), .Y(_88_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_89_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_89_), .Y(_90_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_90_), .C(_81_), .Y(_91_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_86_), .Y(_92_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_92_), .Y(w_C_17_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_93_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_93_), .Y(_94_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_94_), .C(_91_), .Y(_95_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .C(_95_), .Y(_96_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_96_), .Y(w_C_18_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .Y(_97_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add1[18]), .Y(_98_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_98_), .Y(_99_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_99_), .Y(_100_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_101_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(_101_), .Y(_102_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_103_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(_103_), .Y(_104_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_104_), .C(_95_), .Y(_105_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_100_), .Y(_106_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(_106_), .Y(w_C_19_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_107_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_107_), .Y(_108_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_108_), .C(_105_), .Y(_109_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .C(_109_), .Y(_110_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(_110_), .Y(w_C_20_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .Y(_111_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add1[20]), .Y(_112_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_112_), .Y(_113_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_113_), .Y(_114_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_115_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_115_), .Y(_116_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_117_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(_117_), .Y(_118_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_118_), .C(_109_), .Y(_119_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_114_), .Y(_120_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(_120_), .Y(w_C_21_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_121_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(_121_), .Y(_122_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_122_), .C(_119_), .Y(_123_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .C(_123_), .Y(_124_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(_124_), .Y(w_C_22_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .Y(_125_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add1[22]), .Y(_126_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_126_), .Y(_127_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(_127_), .Y(_128_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_129_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_129_), .Y(_130_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_131_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(_131_), .Y(_132_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_132_), .C(_123_), .Y(_133_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_128_), .Y(_134_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_134_), .Y(w_C_23_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_135_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_135_), .Y(_136_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_136_), .C(_133_), .Y(_137_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .C(_137_), .Y(_138_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_138_), .Y(w_C_24_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .Y(_139_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add1[24]), .Y(_140_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_140_), .Y(_141_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(_141_), .Y(_142_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_143_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_143_), .Y(_144_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_145_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(_145_), .Y(_146_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_146_), .C(_137_), .Y(_147_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_142_), .Y(_148_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(_148_), .Y(w_C_25_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_149_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(_149_), .Y(_150_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_150_), .C(_147_), .Y(_151_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .C(_151_), .Y(_152_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(_152_), .Y(w_C_26_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .Y(_153_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add1[26]), .Y(_154_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_154_), .Y(_155_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(_156_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_157_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(_157_), .Y(_158_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_159_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(_159_), .Y(_160_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_160_), .C(_151_), .Y(_161_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_156_), .Y(_162_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(_162_), .Y(w_C_27_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_163_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(_163_), .Y(_164_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_164_), .C(_161_), .Y(_165_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .C(_165_), .Y(_166_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(_166_), .Y(w_C_28_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .Y(_167_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add1[28]), .Y(_168_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_168_), .Y(_169_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(_169_), .Y(_170_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_171_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(_171_), .Y(_172_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_173_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(_173_), .Y(_174_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_174_), .C(_165_), .Y(_175_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_175_), .B(_170_), .Y(_176_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(_176_), .Y(w_C_29_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_177_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(_177_), .Y(_178_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_178_), .C(_175_), .Y(_179_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .C(_179_), .Y(_180_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(_180_), .Y(w_C_30_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .Y(_181_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(i_add1[30]), .Y(_182_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_182_), .Y(_183_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(_183_), .Y(_184_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_185_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(_185_), .Y(_186_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_187_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(_187_), .Y(_188_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_188_), .C(_179_), .Y(_189_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_184_), .Y(_190_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(_190_), .Y(w_C_31_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_191_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(_191_), .Y(_192_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_192_), .C(_189_), .Y(_193_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .C(_193_), .Y(_194_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(_194_), .Y(w_C_32_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .Y(_195_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(i_add1[32]), .Y(_196_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_196_), .Y(_197_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(_197_), .Y(_198_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_199_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(_199_), .Y(_200_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_201_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(_201_), .Y(_202_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_202_), .C(_193_), .Y(_203_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_198_), .Y(_204_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(_204_), .Y(w_C_33_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_205_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(_205_), .Y(_206_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_206_), .C(_203_), .Y(_207_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .C(_207_), .Y(_208_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(_208_), .Y(w_C_34_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .Y(_209_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(i_add1[34]), .Y(_210_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_210_), .Y(_211_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(_211_), .Y(_212_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_213_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(_213_), .Y(_214_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_215_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(_215_), .Y(_216_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_216_), .C(_207_), .Y(_217_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_212_), .Y(_218_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(_218_), .Y(w_C_35_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_219_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(_219_), .Y(_220_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_220_), .C(_217_), .Y(_221_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .C(_221_), .Y(_222_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(_222_), .Y(w_C_36_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_223_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_224_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_222_), .C(_223_), .Y(w_C_37_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_225_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_226_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(_226_), .Y(_227_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(_224_), .Y(_228_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_228_), .C(_221_), .Y(_229_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_230_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_230_), .C(_229_), .Y(_231_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_225_), .Y(w_C_38_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .Y(_232_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(i_add1[38]), .Y(_233_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_233_), .Y(_234_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_234_), .C(_231_), .Y(_235_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_233_), .C(_235_), .Y(w_C_39_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .Y(_236_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(i_add1[39]), .Y(_237_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .C(w_C_39_), .Y(_238_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_237_), .C(_238_), .Y(w_C_40_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .Y(_239_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(i_add1[40]), .Y(_240_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_240_), .Y(_241_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(w_C_40_), .B(_241_), .Y(_242_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .C(_242_), .Y(_243_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(_243_), .Y(w_C_41_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_244_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_245_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_243_), .C(_244_), .Y(w_C_42_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_246_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(_245_), .Y(_247_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(_241_), .Y(_248_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_237_), .Y(_249_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_250_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_251_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_251_), .C(_235_), .Y(_252_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_240_), .Y(_253_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_264__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_264__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_264__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_264__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_264__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_264__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_264__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_264__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_264__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_264__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_264__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_264__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_264__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_264__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_264__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_264__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_264__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_264__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_264__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_264__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_264__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_264__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_264__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_264__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_264__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_264__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_264__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_264__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_264__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_264__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_264__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_264__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_264__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_264__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_264__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_264__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_264__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_264__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_264__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_264__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_264__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_264__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_264__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_264__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_264__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(w_C_45_), .Y(o_result[45]) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_268_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_269_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_270_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_270_), .C(_269_), .Y(_271_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_265_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_266_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_266_), .C(w_C_4_), .Y(_267_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_271_), .Y(_264__4_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_275_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_276_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_277_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_277_), .C(_276_), .Y(_278_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_272_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_273_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_273_), .C(w_C_5_), .Y(_274_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_278_), .Y(_264__5_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_282_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_283_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_284_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_284_), .C(_283_), .Y(_285_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_279_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_280_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_279_), .B(_280_), .C(w_C_6_), .Y(_281_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_285_), .Y(_264__6_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_289_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_290_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_291_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_291_), .C(_290_), .Y(_292_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_286_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_287_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_287_), .C(w_C_7_), .Y(_288_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_292_), .Y(_264__7_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_296_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_297_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_298_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_298_), .C(_297_), .Y(_299_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_293_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_294_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_294_), .C(w_C_8_), .Y(_295_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_299_), .Y(_264__8_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_303_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_304_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_305_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_305_), .C(_304_), .Y(_306_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_300_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_301_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_301_), .C(w_C_9_), .Y(_302_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_306_), .Y(_264__9_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_310_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_311_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_312_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_312_), .C(_311_), .Y(_313_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_307_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_308_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_308_), .C(w_C_10_), .Y(_309_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_313_), .Y(_264__10_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_317_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_318_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_319_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_319_), .C(_318_), .Y(_320_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_314_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_315_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_315_), .C(w_C_11_), .Y(_316_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_316_), .B(_320_), .Y(_264__11_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(w_C_12_), .Y(_324_) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(w_C_45_), .Y(_264__45_) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
