module CSkipA_46bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term1[45], i_add_term1[46], i_add_term1[47], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], i_add_term2[45], i_add_term2[46], i_add_term2[47], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], sum[45], sum[46], sum[47], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term1[45];
input i_add_term1[46];
input i_add_term1[47];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
input i_add_term2[45];
input i_add_term2[46];
input i_add_term2[47];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output sum[45];
output sum[46];
output sum[47];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_11_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_23_) );
OAI21X1 OAI21X1_1 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .C(1'b0), .Y(_24_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_25_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_26_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_27_) );
NAND3X1 NAND3X1_1 ( .A(_25_), .B(_26_), .C(_27_), .Y(_28_) );
OAI21X1 OAI21X1_2 ( .A(_24_), .B(_28_), .C(_23_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3_), .Y(_29_) );
OAI21X1 OAI21X1_3 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .C(1'b0), .Y(_30_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_31_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_32_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_33_) );
NAND3X1 NAND3X1_2 ( .A(_31_), .B(_32_), .C(_33_), .Y(_34_) );
OAI21X1 OAI21X1_4 ( .A(_30_), .B(_34_), .C(_29_), .Y(w_cout_2_) );
INVX1 INVX1_3 ( .A(_5_), .Y(_35_) );
OAI21X1 OAI21X1_5 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .C(1'b0), .Y(_36_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_37_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_38_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_39_) );
NAND3X1 NAND3X1_3 ( .A(_37_), .B(_38_), .C(_39_), .Y(_40_) );
OAI21X1 OAI21X1_6 ( .A(_36_), .B(_40_), .C(_35_), .Y(w_cout_3_) );
INVX1 INVX1_4 ( .A(_7_), .Y(_41_) );
OAI21X1 OAI21X1_7 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .C(1'b0), .Y(_42_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_43_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_44_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_45_) );
NAND3X1 NAND3X1_4 ( .A(_43_), .B(_44_), .C(_45_), .Y(_46_) );
OAI21X1 OAI21X1_8 ( .A(_42_), .B(_46_), .C(_41_), .Y(w_cout_4_) );
INVX1 INVX1_5 ( .A(_9_), .Y(_47_) );
OAI21X1 OAI21X1_9 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .C(1'b0), .Y(_48_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_49_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_50_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_51_) );
NAND3X1 NAND3X1_5 ( .A(_49_), .B(_50_), .C(_51_), .Y(_52_) );
OAI21X1 OAI21X1_10 ( .A(_48_), .B(_52_), .C(_47_), .Y(w_cout_5_) );
INVX1 INVX1_6 ( .A(_11_), .Y(_53_) );
OAI21X1 OAI21X1_11 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .C(1'b0), .Y(_54_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_55_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_56_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_57_) );
NAND3X1 NAND3X1_6 ( .A(_55_), .B(_56_), .C(_57_), .Y(_58_) );
OAI21X1 OAI21X1_12 ( .A(_54_), .B(_58_), .C(_53_), .Y(w_cout_6_) );
INVX1 INVX1_7 ( .A(_13_), .Y(_59_) );
OAI21X1 OAI21X1_13 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .C(1'b0), .Y(_60_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_61_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_62_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_63_) );
NAND3X1 NAND3X1_7 ( .A(_61_), .B(_62_), .C(_63_), .Y(_64_) );
OAI21X1 OAI21X1_14 ( .A(_60_), .B(_64_), .C(_59_), .Y(w_cout_7_) );
INVX1 INVX1_8 ( .A(_15_), .Y(_65_) );
OAI21X1 OAI21X1_15 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .C(1'b0), .Y(_66_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_67_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_68_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_69_) );
NAND3X1 NAND3X1_8 ( .A(_67_), .B(_68_), .C(_69_), .Y(_70_) );
OAI21X1 OAI21X1_16 ( .A(_66_), .B(_70_), .C(_65_), .Y(w_cout_8_) );
INVX1 INVX1_9 ( .A(_17_), .Y(_71_) );
OAI21X1 OAI21X1_17 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .C(1'b0), .Y(_72_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_73_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_74_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_75_) );
NAND3X1 NAND3X1_9 ( .A(_73_), .B(_74_), .C(_75_), .Y(_76_) );
OAI21X1 OAI21X1_18 ( .A(_72_), .B(_76_), .C(_71_), .Y(w_cout_9_) );
INVX1 INVX1_10 ( .A(_19_), .Y(_77_) );
OAI21X1 OAI21X1_19 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .C(1'b0), .Y(_78_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_79_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_80_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_81_) );
NAND3X1 NAND3X1_10 ( .A(_79_), .B(_80_), .C(_81_), .Y(_82_) );
OAI21X1 OAI21X1_20 ( .A(_78_), .B(_82_), .C(_77_), .Y(w_cout_10_) );
INVX1 INVX1_11 ( .A(_21_), .Y(_83_) );
OAI21X1 OAI21X1_21 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .C(1'b0), .Y(_84_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_85_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_86_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_87_) );
NAND3X1 NAND3X1_11 ( .A(_85_), .B(_86_), .C(_87_), .Y(_88_) );
OAI21X1 OAI21X1_22 ( .A(_84_), .B(_88_), .C(_83_), .Y(w_cout_11_) );
INVX1 INVX1_12 ( .A(skip0_cin_next), .Y(_92_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_93_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_94_) );
NAND3X1 NAND3X1_12 ( .A(_92_), .B(_94_), .C(_93_), .Y(_95_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_89_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_90_) );
OAI21X1 OAI21X1_23 ( .A(_89_), .B(_90_), .C(skip0_cin_next), .Y(_91_) );
NAND2X1 NAND2X1_2 ( .A(_91_), .B(_95_), .Y(_0__4_) );
OAI21X1 OAI21X1_24 ( .A(_92_), .B(_89_), .C(_94_), .Y(_2__1_) );
INVX1 INVX1_13 ( .A(_2__1_), .Y(_99_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_100_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_101_) );
NAND3X1 NAND3X1_13 ( .A(_99_), .B(_101_), .C(_100_), .Y(_102_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_96_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_97_) );
OAI21X1 OAI21X1_25 ( .A(_96_), .B(_97_), .C(_2__1_), .Y(_98_) );
NAND2X1 NAND2X1_4 ( .A(_98_), .B(_102_), .Y(_0__5_) );
OAI21X1 OAI21X1_26 ( .A(_99_), .B(_96_), .C(_101_), .Y(_2__2_) );
INVX1 INVX1_14 ( .A(_2__2_), .Y(_106_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_107_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_108_) );
NAND3X1 NAND3X1_14 ( .A(_106_), .B(_108_), .C(_107_), .Y(_109_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_103_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_104_) );
OAI21X1 OAI21X1_27 ( .A(_103_), .B(_104_), .C(_2__2_), .Y(_105_) );
NAND2X1 NAND2X1_6 ( .A(_105_), .B(_109_), .Y(_0__6_) );
OAI21X1 OAI21X1_28 ( .A(_106_), .B(_103_), .C(_108_), .Y(_2__3_) );
INVX1 INVX1_15 ( .A(_2__3_), .Y(_113_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_114_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_115_) );
NAND3X1 NAND3X1_15 ( .A(_113_), .B(_115_), .C(_114_), .Y(_116_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_110_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_111_) );
OAI21X1 OAI21X1_29 ( .A(_110_), .B(_111_), .C(_2__3_), .Y(_112_) );
NAND2X1 NAND2X1_8 ( .A(_112_), .B(_116_), .Y(_0__7_) );
OAI21X1 OAI21X1_30 ( .A(_113_), .B(_110_), .C(_115_), .Y(_1_) );
INVX1 INVX1_16 ( .A(w_cout_1_), .Y(_120_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_121_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_122_) );
NAND3X1 NAND3X1_16 ( .A(_120_), .B(_122_), .C(_121_), .Y(_123_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_117_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_118_) );
OAI21X1 OAI21X1_31 ( .A(_117_), .B(_118_), .C(w_cout_1_), .Y(_119_) );
NAND2X1 NAND2X1_10 ( .A(_119_), .B(_123_), .Y(_0__8_) );
OAI21X1 OAI21X1_32 ( .A(_120_), .B(_117_), .C(_122_), .Y(_4__1_) );
INVX1 INVX1_17 ( .A(_4__1_), .Y(_127_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_128_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_129_) );
NAND3X1 NAND3X1_17 ( .A(_127_), .B(_129_), .C(_128_), .Y(_130_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_124_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_125_) );
OAI21X1 OAI21X1_33 ( .A(_124_), .B(_125_), .C(_4__1_), .Y(_126_) );
NAND2X1 NAND2X1_12 ( .A(_126_), .B(_130_), .Y(_0__9_) );
OAI21X1 OAI21X1_34 ( .A(_127_), .B(_124_), .C(_129_), .Y(_4__2_) );
INVX1 INVX1_18 ( .A(_4__2_), .Y(_134_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_135_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_136_) );
NAND3X1 NAND3X1_18 ( .A(_134_), .B(_136_), .C(_135_), .Y(_137_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_131_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_132_) );
OAI21X1 OAI21X1_35 ( .A(_131_), .B(_132_), .C(_4__2_), .Y(_133_) );
NAND2X1 NAND2X1_14 ( .A(_133_), .B(_137_), .Y(_0__10_) );
OAI21X1 OAI21X1_36 ( .A(_134_), .B(_131_), .C(_136_), .Y(_4__3_) );
INVX1 INVX1_19 ( .A(_4__3_), .Y(_141_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_142_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_143_) );
NAND3X1 NAND3X1_19 ( .A(_141_), .B(_143_), .C(_142_), .Y(_144_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_138_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_139_) );
OAI21X1 OAI21X1_37 ( .A(_138_), .B(_139_), .C(_4__3_), .Y(_140_) );
NAND2X1 NAND2X1_16 ( .A(_140_), .B(_144_), .Y(_0__11_) );
OAI21X1 OAI21X1_38 ( .A(_141_), .B(_138_), .C(_143_), .Y(_3_) );
INVX1 INVX1_20 ( .A(w_cout_2_), .Y(_148_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_149_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_150_) );
NAND3X1 NAND3X1_20 ( .A(_148_), .B(_150_), .C(_149_), .Y(_151_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_145_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_146_) );
OAI21X1 OAI21X1_39 ( .A(_145_), .B(_146_), .C(w_cout_2_), .Y(_147_) );
NAND2X1 NAND2X1_18 ( .A(_147_), .B(_151_), .Y(_0__12_) );
OAI21X1 OAI21X1_40 ( .A(_148_), .B(_145_), .C(_150_), .Y(_6__1_) );
INVX1 INVX1_21 ( .A(_6__1_), .Y(_155_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_156_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_157_) );
NAND3X1 NAND3X1_21 ( .A(_155_), .B(_157_), .C(_156_), .Y(_158_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_152_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_153_) );
OAI21X1 OAI21X1_41 ( .A(_152_), .B(_153_), .C(_6__1_), .Y(_154_) );
NAND2X1 NAND2X1_20 ( .A(_154_), .B(_158_), .Y(_0__13_) );
OAI21X1 OAI21X1_42 ( .A(_155_), .B(_152_), .C(_157_), .Y(_6__2_) );
INVX1 INVX1_22 ( .A(_6__2_), .Y(_162_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_163_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_164_) );
NAND3X1 NAND3X1_22 ( .A(_162_), .B(_164_), .C(_163_), .Y(_165_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_159_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_160_) );
OAI21X1 OAI21X1_43 ( .A(_159_), .B(_160_), .C(_6__2_), .Y(_161_) );
NAND2X1 NAND2X1_22 ( .A(_161_), .B(_165_), .Y(_0__14_) );
OAI21X1 OAI21X1_44 ( .A(_162_), .B(_159_), .C(_164_), .Y(_6__3_) );
INVX1 INVX1_23 ( .A(_6__3_), .Y(_169_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_170_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_171_) );
NAND3X1 NAND3X1_23 ( .A(_169_), .B(_171_), .C(_170_), .Y(_172_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_166_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_167_) );
OAI21X1 OAI21X1_45 ( .A(_166_), .B(_167_), .C(_6__3_), .Y(_168_) );
NAND2X1 NAND2X1_24 ( .A(_168_), .B(_172_), .Y(_0__15_) );
OAI21X1 OAI21X1_46 ( .A(_169_), .B(_166_), .C(_171_), .Y(_5_) );
INVX1 INVX1_24 ( .A(w_cout_3_), .Y(_176_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_177_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_178_) );
NAND3X1 NAND3X1_24 ( .A(_176_), .B(_178_), .C(_177_), .Y(_179_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_173_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_174_) );
OAI21X1 OAI21X1_47 ( .A(_173_), .B(_174_), .C(w_cout_3_), .Y(_175_) );
NAND2X1 NAND2X1_26 ( .A(_175_), .B(_179_), .Y(_0__16_) );
OAI21X1 OAI21X1_48 ( .A(_176_), .B(_173_), .C(_178_), .Y(_8__1_) );
INVX1 INVX1_25 ( .A(_8__1_), .Y(_183_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_184_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_185_) );
NAND3X1 NAND3X1_25 ( .A(_183_), .B(_185_), .C(_184_), .Y(_186_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_180_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_181_) );
OAI21X1 OAI21X1_49 ( .A(_180_), .B(_181_), .C(_8__1_), .Y(_182_) );
NAND2X1 NAND2X1_28 ( .A(_182_), .B(_186_), .Y(_0__17_) );
OAI21X1 OAI21X1_50 ( .A(_183_), .B(_180_), .C(_185_), .Y(_8__2_) );
INVX1 INVX1_26 ( .A(_8__2_), .Y(_190_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_191_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_192_) );
NAND3X1 NAND3X1_26 ( .A(_190_), .B(_192_), .C(_191_), .Y(_193_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_187_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_188_) );
OAI21X1 OAI21X1_51 ( .A(_187_), .B(_188_), .C(_8__2_), .Y(_189_) );
NAND2X1 NAND2X1_30 ( .A(_189_), .B(_193_), .Y(_0__18_) );
OAI21X1 OAI21X1_52 ( .A(_190_), .B(_187_), .C(_192_), .Y(_8__3_) );
INVX1 INVX1_27 ( .A(_8__3_), .Y(_197_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_198_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_199_) );
NAND3X1 NAND3X1_27 ( .A(_197_), .B(_199_), .C(_198_), .Y(_200_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_194_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_195_) );
OAI21X1 OAI21X1_53 ( .A(_194_), .B(_195_), .C(_8__3_), .Y(_196_) );
NAND2X1 NAND2X1_32 ( .A(_196_), .B(_200_), .Y(_0__19_) );
OAI21X1 OAI21X1_54 ( .A(_197_), .B(_194_), .C(_199_), .Y(_7_) );
INVX1 INVX1_28 ( .A(w_cout_4_), .Y(_204_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_205_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_206_) );
NAND3X1 NAND3X1_28 ( .A(_204_), .B(_206_), .C(_205_), .Y(_207_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_201_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_202_) );
OAI21X1 OAI21X1_55 ( .A(_201_), .B(_202_), .C(w_cout_4_), .Y(_203_) );
NAND2X1 NAND2X1_34 ( .A(_203_), .B(_207_), .Y(_0__20_) );
OAI21X1 OAI21X1_56 ( .A(_204_), .B(_201_), .C(_206_), .Y(_10__1_) );
INVX1 INVX1_29 ( .A(_10__1_), .Y(_211_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_212_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_213_) );
NAND3X1 NAND3X1_29 ( .A(_211_), .B(_213_), .C(_212_), .Y(_214_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_208_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_209_) );
OAI21X1 OAI21X1_57 ( .A(_208_), .B(_209_), .C(_10__1_), .Y(_210_) );
NAND2X1 NAND2X1_36 ( .A(_210_), .B(_214_), .Y(_0__21_) );
OAI21X1 OAI21X1_58 ( .A(_211_), .B(_208_), .C(_213_), .Y(_10__2_) );
INVX1 INVX1_30 ( .A(_10__2_), .Y(_218_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_219_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_220_) );
NAND3X1 NAND3X1_30 ( .A(_218_), .B(_220_), .C(_219_), .Y(_221_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_215_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_216_) );
OAI21X1 OAI21X1_59 ( .A(_215_), .B(_216_), .C(_10__2_), .Y(_217_) );
NAND2X1 NAND2X1_38 ( .A(_217_), .B(_221_), .Y(_0__22_) );
OAI21X1 OAI21X1_60 ( .A(_218_), .B(_215_), .C(_220_), .Y(_10__3_) );
INVX1 INVX1_31 ( .A(_10__3_), .Y(_225_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_226_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_227_) );
NAND3X1 NAND3X1_31 ( .A(_225_), .B(_227_), .C(_226_), .Y(_228_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_222_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_223_) );
OAI21X1 OAI21X1_61 ( .A(_222_), .B(_223_), .C(_10__3_), .Y(_224_) );
NAND2X1 NAND2X1_40 ( .A(_224_), .B(_228_), .Y(_0__23_) );
OAI21X1 OAI21X1_62 ( .A(_225_), .B(_222_), .C(_227_), .Y(_9_) );
INVX1 INVX1_32 ( .A(w_cout_5_), .Y(_232_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_233_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_234_) );
NAND3X1 NAND3X1_32 ( .A(_232_), .B(_234_), .C(_233_), .Y(_235_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_229_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_230_) );
OAI21X1 OAI21X1_63 ( .A(_229_), .B(_230_), .C(w_cout_5_), .Y(_231_) );
NAND2X1 NAND2X1_42 ( .A(_231_), .B(_235_), .Y(_0__24_) );
OAI21X1 OAI21X1_64 ( .A(_232_), .B(_229_), .C(_234_), .Y(_12__1_) );
INVX1 INVX1_33 ( .A(_12__1_), .Y(_239_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_240_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_241_) );
NAND3X1 NAND3X1_33 ( .A(_239_), .B(_241_), .C(_240_), .Y(_242_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_236_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_237_) );
OAI21X1 OAI21X1_65 ( .A(_236_), .B(_237_), .C(_12__1_), .Y(_238_) );
NAND2X1 NAND2X1_44 ( .A(_238_), .B(_242_), .Y(_0__25_) );
OAI21X1 OAI21X1_66 ( .A(_239_), .B(_236_), .C(_241_), .Y(_12__2_) );
INVX1 INVX1_34 ( .A(_12__2_), .Y(_246_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_247_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_248_) );
NAND3X1 NAND3X1_34 ( .A(_246_), .B(_248_), .C(_247_), .Y(_249_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_243_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_244_) );
OAI21X1 OAI21X1_67 ( .A(_243_), .B(_244_), .C(_12__2_), .Y(_245_) );
NAND2X1 NAND2X1_46 ( .A(_245_), .B(_249_), .Y(_0__26_) );
OAI21X1 OAI21X1_68 ( .A(_246_), .B(_243_), .C(_248_), .Y(_12__3_) );
INVX1 INVX1_35 ( .A(_12__3_), .Y(_253_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_254_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_255_) );
NAND3X1 NAND3X1_35 ( .A(_253_), .B(_255_), .C(_254_), .Y(_256_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_250_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_251_) );
OAI21X1 OAI21X1_69 ( .A(_250_), .B(_251_), .C(_12__3_), .Y(_252_) );
NAND2X1 NAND2X1_48 ( .A(_252_), .B(_256_), .Y(_0__27_) );
OAI21X1 OAI21X1_70 ( .A(_253_), .B(_250_), .C(_255_), .Y(_11_) );
INVX1 INVX1_36 ( .A(w_cout_6_), .Y(_260_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_261_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_262_) );
NAND3X1 NAND3X1_36 ( .A(_260_), .B(_262_), .C(_261_), .Y(_263_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_257_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_258_) );
OAI21X1 OAI21X1_71 ( .A(_257_), .B(_258_), .C(w_cout_6_), .Y(_259_) );
NAND2X1 NAND2X1_50 ( .A(_259_), .B(_263_), .Y(_0__28_) );
OAI21X1 OAI21X1_72 ( .A(_260_), .B(_257_), .C(_262_), .Y(_14__1_) );
INVX1 INVX1_37 ( .A(_14__1_), .Y(_267_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_268_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_269_) );
NAND3X1 NAND3X1_37 ( .A(_267_), .B(_269_), .C(_268_), .Y(_270_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_264_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_265_) );
OAI21X1 OAI21X1_73 ( .A(_264_), .B(_265_), .C(_14__1_), .Y(_266_) );
NAND2X1 NAND2X1_52 ( .A(_266_), .B(_270_), .Y(_0__29_) );
OAI21X1 OAI21X1_74 ( .A(_267_), .B(_264_), .C(_269_), .Y(_14__2_) );
INVX1 INVX1_38 ( .A(_14__2_), .Y(_274_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_275_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_276_) );
NAND3X1 NAND3X1_38 ( .A(_274_), .B(_276_), .C(_275_), .Y(_277_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_271_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_272_) );
OAI21X1 OAI21X1_75 ( .A(_271_), .B(_272_), .C(_14__2_), .Y(_273_) );
NAND2X1 NAND2X1_54 ( .A(_273_), .B(_277_), .Y(_0__30_) );
OAI21X1 OAI21X1_76 ( .A(_274_), .B(_271_), .C(_276_), .Y(_14__3_) );
INVX1 INVX1_39 ( .A(_14__3_), .Y(_281_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_282_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_283_) );
NAND3X1 NAND3X1_39 ( .A(_281_), .B(_283_), .C(_282_), .Y(_284_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_278_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_279_) );
OAI21X1 OAI21X1_77 ( .A(_278_), .B(_279_), .C(_14__3_), .Y(_280_) );
NAND2X1 NAND2X1_56 ( .A(_280_), .B(_284_), .Y(_0__31_) );
OAI21X1 OAI21X1_78 ( .A(_281_), .B(_278_), .C(_283_), .Y(_13_) );
INVX1 INVX1_40 ( .A(w_cout_7_), .Y(_288_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_289_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_290_) );
NAND3X1 NAND3X1_40 ( .A(_288_), .B(_290_), .C(_289_), .Y(_291_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_285_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_286_) );
OAI21X1 OAI21X1_79 ( .A(_285_), .B(_286_), .C(w_cout_7_), .Y(_287_) );
NAND2X1 NAND2X1_58 ( .A(_287_), .B(_291_), .Y(_0__32_) );
OAI21X1 OAI21X1_80 ( .A(_288_), .B(_285_), .C(_290_), .Y(_16__1_) );
INVX1 INVX1_41 ( .A(_16__1_), .Y(_295_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_296_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_297_) );
NAND3X1 NAND3X1_41 ( .A(_295_), .B(_297_), .C(_296_), .Y(_298_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_292_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_293_) );
OAI21X1 OAI21X1_81 ( .A(_292_), .B(_293_), .C(_16__1_), .Y(_294_) );
NAND2X1 NAND2X1_60 ( .A(_294_), .B(_298_), .Y(_0__33_) );
OAI21X1 OAI21X1_82 ( .A(_295_), .B(_292_), .C(_297_), .Y(_16__2_) );
INVX1 INVX1_42 ( .A(_16__2_), .Y(_302_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_303_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_304_) );
NAND3X1 NAND3X1_42 ( .A(_302_), .B(_304_), .C(_303_), .Y(_305_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_299_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_300_) );
OAI21X1 OAI21X1_83 ( .A(_299_), .B(_300_), .C(_16__2_), .Y(_301_) );
NAND2X1 NAND2X1_62 ( .A(_301_), .B(_305_), .Y(_0__34_) );
OAI21X1 OAI21X1_84 ( .A(_302_), .B(_299_), .C(_304_), .Y(_16__3_) );
INVX1 INVX1_43 ( .A(_16__3_), .Y(_309_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_310_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_311_) );
NAND3X1 NAND3X1_43 ( .A(_309_), .B(_311_), .C(_310_), .Y(_312_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_306_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_307_) );
OAI21X1 OAI21X1_85 ( .A(_306_), .B(_307_), .C(_16__3_), .Y(_308_) );
NAND2X1 NAND2X1_64 ( .A(_308_), .B(_312_), .Y(_0__35_) );
OAI21X1 OAI21X1_86 ( .A(_309_), .B(_306_), .C(_311_), .Y(_15_) );
INVX1 INVX1_44 ( .A(w_cout_8_), .Y(_316_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_317_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_318_) );
NAND3X1 NAND3X1_44 ( .A(_316_), .B(_318_), .C(_317_), .Y(_319_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_313_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_314_) );
OAI21X1 OAI21X1_87 ( .A(_313_), .B(_314_), .C(w_cout_8_), .Y(_315_) );
NAND2X1 NAND2X1_66 ( .A(_315_), .B(_319_), .Y(_0__36_) );
OAI21X1 OAI21X1_88 ( .A(_316_), .B(_313_), .C(_318_), .Y(_18__1_) );
INVX1 INVX1_45 ( .A(_18__1_), .Y(_323_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_324_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_325_) );
NAND3X1 NAND3X1_45 ( .A(_323_), .B(_325_), .C(_324_), .Y(_326_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_320_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_321_) );
OAI21X1 OAI21X1_89 ( .A(_320_), .B(_321_), .C(_18__1_), .Y(_322_) );
NAND2X1 NAND2X1_68 ( .A(_322_), .B(_326_), .Y(_0__37_) );
OAI21X1 OAI21X1_90 ( .A(_323_), .B(_320_), .C(_325_), .Y(_18__2_) );
INVX1 INVX1_46 ( .A(_18__2_), .Y(_330_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_331_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_332_) );
NAND3X1 NAND3X1_46 ( .A(_330_), .B(_332_), .C(_331_), .Y(_333_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_327_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_328_) );
OAI21X1 OAI21X1_91 ( .A(_327_), .B(_328_), .C(_18__2_), .Y(_329_) );
NAND2X1 NAND2X1_70 ( .A(_329_), .B(_333_), .Y(_0__38_) );
OAI21X1 OAI21X1_92 ( .A(_330_), .B(_327_), .C(_332_), .Y(_18__3_) );
INVX1 INVX1_47 ( .A(_18__3_), .Y(_337_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_338_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_339_) );
NAND3X1 NAND3X1_47 ( .A(_337_), .B(_339_), .C(_338_), .Y(_340_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_334_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_335_) );
OAI21X1 OAI21X1_93 ( .A(_334_), .B(_335_), .C(_18__3_), .Y(_336_) );
NAND2X1 NAND2X1_72 ( .A(_336_), .B(_340_), .Y(_0__39_) );
OAI21X1 OAI21X1_94 ( .A(_337_), .B(_334_), .C(_339_), .Y(_17_) );
INVX1 INVX1_48 ( .A(w_cout_9_), .Y(_344_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_345_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_346_) );
NAND3X1 NAND3X1_48 ( .A(_344_), .B(_346_), .C(_345_), .Y(_347_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_341_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_342_) );
OAI21X1 OAI21X1_95 ( .A(_341_), .B(_342_), .C(w_cout_9_), .Y(_343_) );
NAND2X1 NAND2X1_74 ( .A(_343_), .B(_347_), .Y(_0__40_) );
OAI21X1 OAI21X1_96 ( .A(_344_), .B(_341_), .C(_346_), .Y(_20__1_) );
INVX1 INVX1_49 ( .A(_20__1_), .Y(_351_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_352_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_353_) );
NAND3X1 NAND3X1_49 ( .A(_351_), .B(_353_), .C(_352_), .Y(_354_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_348_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_349_) );
OAI21X1 OAI21X1_97 ( .A(_348_), .B(_349_), .C(_20__1_), .Y(_350_) );
NAND2X1 NAND2X1_76 ( .A(_350_), .B(_354_), .Y(_0__41_) );
OAI21X1 OAI21X1_98 ( .A(_351_), .B(_348_), .C(_353_), .Y(_20__2_) );
INVX1 INVX1_50 ( .A(_20__2_), .Y(_358_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_359_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_360_) );
NAND3X1 NAND3X1_50 ( .A(_358_), .B(_360_), .C(_359_), .Y(_361_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_355_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_356_) );
OAI21X1 OAI21X1_99 ( .A(_355_), .B(_356_), .C(_20__2_), .Y(_357_) );
NAND2X1 NAND2X1_78 ( .A(_357_), .B(_361_), .Y(_0__42_) );
OAI21X1 OAI21X1_100 ( .A(_358_), .B(_355_), .C(_360_), .Y(_20__3_) );
INVX1 INVX1_51 ( .A(_20__3_), .Y(_365_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_366_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_367_) );
NAND3X1 NAND3X1_51 ( .A(_365_), .B(_367_), .C(_366_), .Y(_368_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_362_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_363_) );
OAI21X1 OAI21X1_101 ( .A(_362_), .B(_363_), .C(_20__3_), .Y(_364_) );
NAND2X1 NAND2X1_80 ( .A(_364_), .B(_368_), .Y(_0__43_) );
OAI21X1 OAI21X1_102 ( .A(_365_), .B(_362_), .C(_367_), .Y(_19_) );
INVX1 INVX1_52 ( .A(w_cout_10_), .Y(_372_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_373_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_374_) );
NAND3X1 NAND3X1_52 ( .A(_372_), .B(_374_), .C(_373_), .Y(_375_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_369_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_370_) );
OAI21X1 OAI21X1_103 ( .A(_369_), .B(_370_), .C(w_cout_10_), .Y(_371_) );
NAND2X1 NAND2X1_82 ( .A(_371_), .B(_375_), .Y(_0__44_) );
OAI21X1 OAI21X1_104 ( .A(_372_), .B(_369_), .C(_374_), .Y(_22__1_) );
INVX1 INVX1_53 ( .A(_22__1_), .Y(_379_) );
OR2X2 OR2X2_75 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_380_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_381_) );
NAND3X1 NAND3X1_53 ( .A(_379_), .B(_381_), .C(_380_), .Y(_382_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_376_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_377_) );
OAI21X1 OAI21X1_105 ( .A(_376_), .B(_377_), .C(_22__1_), .Y(_378_) );
NAND2X1 NAND2X1_84 ( .A(_378_), .B(_382_), .Y(_0__45_) );
OAI21X1 OAI21X1_106 ( .A(_379_), .B(_376_), .C(_381_), .Y(_22__2_) );
INVX1 INVX1_54 ( .A(_22__2_), .Y(_386_) );
OR2X2 OR2X2_76 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_387_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_388_) );
NAND3X1 NAND3X1_54 ( .A(_386_), .B(_388_), .C(_387_), .Y(_389_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_383_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_384_) );
OAI21X1 OAI21X1_107 ( .A(_383_), .B(_384_), .C(_22__2_), .Y(_385_) );
NAND2X1 NAND2X1_86 ( .A(_385_), .B(_389_), .Y(_0__46_) );
OAI21X1 OAI21X1_108 ( .A(_386_), .B(_383_), .C(_388_), .Y(_22__3_) );
INVX1 INVX1_55 ( .A(_22__3_), .Y(_393_) );
OR2X2 OR2X2_77 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_394_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_395_) );
NAND3X1 NAND3X1_55 ( .A(_393_), .B(_395_), .C(_394_), .Y(_396_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_390_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_391_) );
OAI21X1 OAI21X1_109 ( .A(_390_), .B(_391_), .C(_22__3_), .Y(_392_) );
NAND2X1 NAND2X1_88 ( .A(_392_), .B(_396_), .Y(_0__47_) );
OAI21X1 OAI21X1_110 ( .A(_393_), .B(_390_), .C(_395_), .Y(_21_) );
INVX1 INVX1_56 ( .A(1'b0), .Y(_400_) );
OR2X2 OR2X2_78 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_401_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_402_) );
NAND3X1 NAND3X1_56 ( .A(_400_), .B(_402_), .C(_401_), .Y(_403_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_397_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_398_) );
OAI21X1 OAI21X1_111 ( .A(_397_), .B(_398_), .C(1'b0), .Y(_399_) );
NAND2X1 NAND2X1_90 ( .A(_399_), .B(_403_), .Y(_0__0_) );
OAI21X1 OAI21X1_112 ( .A(_400_), .B(_397_), .C(_402_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_57 ( .A(rca_inst_w_CARRY_1_), .Y(_407_) );
OR2X2 OR2X2_79 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_408_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_409_) );
NAND3X1 NAND3X1_57 ( .A(_407_), .B(_409_), .C(_408_), .Y(_410_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_404_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_405_) );
OAI21X1 OAI21X1_113 ( .A(_404_), .B(_405_), .C(rca_inst_w_CARRY_1_), .Y(_406_) );
NAND2X1 NAND2X1_92 ( .A(_406_), .B(_410_), .Y(_0__1_) );
OAI21X1 OAI21X1_114 ( .A(_407_), .B(_404_), .C(_409_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_58 ( .A(rca_inst_w_CARRY_2_), .Y(_414_) );
OR2X2 OR2X2_80 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_415_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_416_) );
NAND3X1 NAND3X1_58 ( .A(_414_), .B(_416_), .C(_415_), .Y(_417_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_411_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_412_) );
OAI21X1 OAI21X1_115 ( .A(_411_), .B(_412_), .C(rca_inst_w_CARRY_2_), .Y(_413_) );
NAND2X1 NAND2X1_94 ( .A(_413_), .B(_417_), .Y(_0__2_) );
OAI21X1 OAI21X1_116 ( .A(_414_), .B(_411_), .C(_416_), .Y(rca_inst_w_CARRY_3_) );
INVX1 INVX1_59 ( .A(rca_inst_w_CARRY_3_), .Y(_421_) );
OR2X2 OR2X2_81 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_422_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_423_) );
NAND3X1 NAND3X1_59 ( .A(_421_), .B(_423_), .C(_422_), .Y(_424_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_418_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_419_) );
OAI21X1 OAI21X1_117 ( .A(_418_), .B(_419_), .C(rca_inst_w_CARRY_3_), .Y(_420_) );
NAND2X1 NAND2X1_96 ( .A(_420_), .B(_424_), .Y(_0__3_) );
OAI21X1 OAI21X1_118 ( .A(_421_), .B(_418_), .C(_423_), .Y(cout0) );
INVX1 INVX1_60 ( .A(cout0), .Y(_425_) );
OAI21X1 OAI21X1_119 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .C(1'b0), .Y(_426_) );
OR2X2 OR2X2_82 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_427_) );
OR2X2 OR2X2_83 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_428_) );
OR2X2 OR2X2_84 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_429_) );
NAND3X1 NAND3X1_60 ( .A(_427_), .B(_428_), .C(_429_), .Y(_430_) );
OAI21X1 OAI21X1_120 ( .A(_426_), .B(_430_), .C(_425_), .Y(skip0_cin_next) );
BUFX2 BUFX2_50 ( .A(skip0_cin_next), .Y(_2__0_) );
BUFX2 BUFX2_51 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_52 ( .A(w_cout_1_), .Y(_4__0_) );
BUFX2 BUFX2_53 ( .A(_3_), .Y(_4__4_) );
BUFX2 BUFX2_54 ( .A(w_cout_2_), .Y(_6__0_) );
BUFX2 BUFX2_55 ( .A(_5_), .Y(_6__4_) );
BUFX2 BUFX2_56 ( .A(w_cout_3_), .Y(_8__0_) );
BUFX2 BUFX2_57 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_58 ( .A(w_cout_4_), .Y(_10__0_) );
BUFX2 BUFX2_59 ( .A(_9_), .Y(_10__4_) );
BUFX2 BUFX2_60 ( .A(w_cout_5_), .Y(_12__0_) );
BUFX2 BUFX2_61 ( .A(_11_), .Y(_12__4_) );
BUFX2 BUFX2_62 ( .A(w_cout_6_), .Y(_14__0_) );
BUFX2 BUFX2_63 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_64 ( .A(w_cout_7_), .Y(_16__0_) );
BUFX2 BUFX2_65 ( .A(_15_), .Y(_16__4_) );
BUFX2 BUFX2_66 ( .A(w_cout_8_), .Y(_18__0_) );
BUFX2 BUFX2_67 ( .A(_17_), .Y(_18__4_) );
BUFX2 BUFX2_68 ( .A(w_cout_9_), .Y(_20__0_) );
BUFX2 BUFX2_69 ( .A(_19_), .Y(_20__4_) );
BUFX2 BUFX2_70 ( .A(w_cout_10_), .Y(_22__0_) );
BUFX2 BUFX2_71 ( .A(_21_), .Y(_22__4_) );
BUFX2 BUFX2_72 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_73 ( .A(cout0), .Y(rca_inst_w_CARRY_4_) );
BUFX2 BUFX2_74 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
