module cla_61bit (i_add1, i_add2, o_result);

input [60:0] i_add1;
input [60:0] i_add2;
output [61:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

NOR2X1 NOR2X1_1 ( .A(_233_), .B(_234_), .Y(_240_) );
INVX1 INVX1_1 ( .A(_240_), .Y(_241_) );
AND2X2 AND2X2_1 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_242_) );
INVX1 INVX1_2 ( .A(_242_), .Y(_243_) );
NAND3X1 NAND3X1_1 ( .A(_241_), .B(_243_), .C(_239_), .Y(_244_) );
OAI21X1 OAI21X1_1 ( .A(i_add2[41]), .B(i_add1[41]), .C(_244_), .Y(_245_) );
INVX1 INVX1_3 ( .A(_245_), .Y(w_C_42_) );
INVX1 INVX1_4 ( .A(i_add2[42]), .Y(_246_) );
INVX1 INVX1_5 ( .A(i_add1[42]), .Y(_247_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_248_) );
INVX1 INVX1_6 ( .A(_248_), .Y(_249_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_250_) );
INVX1 INVX1_7 ( .A(_250_), .Y(_251_) );
NAND3X1 NAND3X1_2 ( .A(_249_), .B(_251_), .C(_244_), .Y(_252_) );
OAI21X1 OAI21X1_2 ( .A(_246_), .B(_247_), .C(_252_), .Y(w_C_43_) );
NOR2X1 NOR2X1_4 ( .A(_246_), .B(_247_), .Y(_253_) );
INVX1 INVX1_8 ( .A(_253_), .Y(_254_) );
AND2X2 AND2X2_2 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_255_) );
INVX1 INVX1_9 ( .A(_255_), .Y(_256_) );
NAND3X1 NAND3X1_3 ( .A(_254_), .B(_256_), .C(_252_), .Y(_257_) );
OAI21X1 OAI21X1_3 ( .A(i_add2[43]), .B(i_add1[43]), .C(_257_), .Y(_258_) );
INVX1 INVX1_10 ( .A(_258_), .Y(w_C_44_) );
INVX1 INVX1_11 ( .A(i_add2[44]), .Y(_259_) );
INVX1 INVX1_12 ( .A(i_add1[44]), .Y(_260_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_261_) );
INVX1 INVX1_13 ( .A(_261_), .Y(_262_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_263_) );
INVX1 INVX1_14 ( .A(_263_), .Y(_264_) );
NAND3X1 NAND3X1_4 ( .A(_262_), .B(_264_), .C(_257_), .Y(_265_) );
OAI21X1 OAI21X1_4 ( .A(_259_), .B(_260_), .C(_265_), .Y(w_C_45_) );
NOR2X1 NOR2X1_7 ( .A(_259_), .B(_260_), .Y(_266_) );
INVX1 INVX1_15 ( .A(_266_), .Y(_267_) );
AND2X2 AND2X2_3 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_268_) );
INVX1 INVX1_16 ( .A(_268_), .Y(_269_) );
NAND3X1 NAND3X1_5 ( .A(_267_), .B(_269_), .C(_265_), .Y(_270_) );
OAI21X1 OAI21X1_5 ( .A(i_add2[45]), .B(i_add1[45]), .C(_270_), .Y(_271_) );
INVX1 INVX1_17 ( .A(_271_), .Y(w_C_46_) );
INVX1 INVX1_18 ( .A(i_add2[46]), .Y(_272_) );
INVX1 INVX1_19 ( .A(i_add1[46]), .Y(_273_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_274_) );
INVX1 INVX1_20 ( .A(_274_), .Y(_275_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_276_) );
INVX1 INVX1_21 ( .A(_276_), .Y(_277_) );
NAND3X1 NAND3X1_6 ( .A(_275_), .B(_277_), .C(_270_), .Y(_278_) );
OAI21X1 OAI21X1_6 ( .A(_272_), .B(_273_), .C(_278_), .Y(w_C_47_) );
NOR2X1 NOR2X1_10 ( .A(_272_), .B(_273_), .Y(_279_) );
INVX1 INVX1_22 ( .A(_279_), .Y(_280_) );
AND2X2 AND2X2_4 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_281_) );
INVX1 INVX1_23 ( .A(_281_), .Y(_282_) );
NAND3X1 NAND3X1_7 ( .A(_280_), .B(_282_), .C(_278_), .Y(_283_) );
OAI21X1 OAI21X1_7 ( .A(i_add2[47]), .B(i_add1[47]), .C(_283_), .Y(_284_) );
INVX1 INVX1_24 ( .A(_284_), .Y(w_C_48_) );
INVX1 INVX1_25 ( .A(i_add2[48]), .Y(_285_) );
INVX1 INVX1_26 ( .A(i_add1[48]), .Y(_286_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_287_) );
INVX1 INVX1_27 ( .A(_287_), .Y(_288_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_289_) );
INVX1 INVX1_28 ( .A(_289_), .Y(_290_) );
NAND3X1 NAND3X1_8 ( .A(_288_), .B(_290_), .C(_283_), .Y(_291_) );
OAI21X1 OAI21X1_8 ( .A(_285_), .B(_286_), .C(_291_), .Y(w_C_49_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_292_) );
INVX1 INVX1_29 ( .A(_292_), .Y(_293_) );
NOR2X1 NOR2X1_14 ( .A(_285_), .B(_286_), .Y(_294_) );
INVX1 INVX1_30 ( .A(_294_), .Y(_295_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_296_) );
NAND3X1 NAND3X1_9 ( .A(_295_), .B(_296_), .C(_291_), .Y(_297_) );
AND2X2 AND2X2_5 ( .A(_297_), .B(_293_), .Y(w_C_50_) );
INVX1 INVX1_31 ( .A(i_add2[50]), .Y(_298_) );
INVX1 INVX1_32 ( .A(i_add1[50]), .Y(_299_) );
NAND2X1 NAND2X1_2 ( .A(_298_), .B(_299_), .Y(_300_) );
NAND3X1 NAND3X1_10 ( .A(_293_), .B(_300_), .C(_297_), .Y(_301_) );
OAI21X1 OAI21X1_9 ( .A(_298_), .B(_299_), .C(_301_), .Y(w_C_51_) );
INVX1 INVX1_33 ( .A(i_add2[51]), .Y(_302_) );
INVX1 INVX1_34 ( .A(i_add1[51]), .Y(_303_) );
OAI21X1 OAI21X1_10 ( .A(i_add2[51]), .B(i_add1[51]), .C(w_C_51_), .Y(_304_) );
OAI21X1 OAI21X1_11 ( .A(_302_), .B(_303_), .C(_304_), .Y(w_C_52_) );
INVX1 INVX1_35 ( .A(i_add2[52]), .Y(_305_) );
INVX1 INVX1_36 ( .A(i_add1[52]), .Y(_306_) );
NOR2X1 NOR2X1_15 ( .A(_305_), .B(_306_), .Y(_307_) );
OR2X2 OR2X2_1 ( .A(w_C_52_), .B(_307_), .Y(_308_) );
OAI21X1 OAI21X1_12 ( .A(i_add2[52]), .B(i_add1[52]), .C(_308_), .Y(_309_) );
INVX1 INVX1_37 ( .A(_309_), .Y(w_C_53_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_310_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_311_) );
OAI21X1 OAI21X1_13 ( .A(_311_), .B(_309_), .C(_310_), .Y(w_C_54_) );
INVX1 INVX1_38 ( .A(i_add2[54]), .Y(_312_) );
INVX1 INVX1_39 ( .A(i_add1[54]), .Y(_313_) );
INVX1 INVX1_40 ( .A(_311_), .Y(_314_) );
INVX1 INVX1_41 ( .A(_307_), .Y(_315_) );
NAND2X1 NAND2X1_4 ( .A(_302_), .B(_303_), .Y(_316_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_317_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_318_) );
NAND3X1 NAND3X1_11 ( .A(_317_), .B(_318_), .C(_301_), .Y(_319_) );
NAND2X1 NAND2X1_7 ( .A(_305_), .B(_306_), .Y(_320_) );
NAND3X1 NAND3X1_12 ( .A(_316_), .B(_320_), .C(_319_), .Y(_321_) );
NAND3X1 NAND3X1_13 ( .A(_315_), .B(_310_), .C(_321_), .Y(_322_) );
NAND2X1 NAND2X1_8 ( .A(_312_), .B(_313_), .Y(_323_) );
NAND3X1 NAND3X1_14 ( .A(_314_), .B(_323_), .C(_322_), .Y(_324_) );
OAI21X1 OAI21X1_14 ( .A(_312_), .B(_313_), .C(_324_), .Y(w_C_55_) );
INVX1 INVX1_42 ( .A(i_add2[55]), .Y(_325_) );
INVX1 INVX1_43 ( .A(i_add1[55]), .Y(_326_) );
OAI21X1 OAI21X1_15 ( .A(i_add2[55]), .B(i_add1[55]), .C(w_C_55_), .Y(_327_) );
OAI21X1 OAI21X1_16 ( .A(_325_), .B(_326_), .C(_327_), .Y(w_C_56_) );
NOR2X1 NOR2X1_17 ( .A(_325_), .B(_326_), .Y(_328_) );
INVX1 INVX1_44 ( .A(_328_), .Y(_329_) );
AND2X2 AND2X2_6 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_330_) );
INVX1 INVX1_45 ( .A(_330_), .Y(_331_) );
NAND3X1 NAND3X1_15 ( .A(_329_), .B(_331_), .C(_327_), .Y(_332_) );
OAI21X1 OAI21X1_17 ( .A(i_add2[56]), .B(i_add1[56]), .C(_332_), .Y(_333_) );
INVX1 INVX1_46 ( .A(_333_), .Y(w_C_57_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_334_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_335_) );
OAI21X1 OAI21X1_18 ( .A(_335_), .B(_333_), .C(_334_), .Y(w_C_58_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[58]), .B(i_add1[58]), .Y(_336_) );
INVX1 INVX1_47 ( .A(_335_), .Y(_337_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_338_) );
INVX1 INVX1_48 ( .A(_338_), .Y(_339_) );
NOR2X1 NOR2X1_20 ( .A(_312_), .B(_313_), .Y(_340_) );
INVX1 INVX1_49 ( .A(_340_), .Y(_341_) );
NAND3X1 NAND3X1_16 ( .A(_341_), .B(_329_), .C(_324_), .Y(_342_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_343_) );
INVX1 INVX1_50 ( .A(_343_), .Y(_344_) );
NAND3X1 NAND3X1_17 ( .A(_339_), .B(_344_), .C(_342_), .Y(_345_) );
NAND3X1 NAND3X1_18 ( .A(_331_), .B(_334_), .C(_345_), .Y(_346_) );
OR2X2 OR2X2_2 ( .A(i_add2[58]), .B(i_add1[58]), .Y(_347_) );
NAND3X1 NAND3X1_19 ( .A(_337_), .B(_347_), .C(_346_), .Y(_348_) );
NAND2X1 NAND2X1_11 ( .A(_336_), .B(_348_), .Y(w_C_59_) );
OR2X2 OR2X2_3 ( .A(i_add2[59]), .B(i_add1[59]), .Y(_349_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[59]), .B(i_add1[59]), .Y(_350_) );
NAND3X1 NAND3X1_20 ( .A(_336_), .B(_350_), .C(_348_), .Y(_351_) );
AND2X2 AND2X2_7 ( .A(_351_), .B(_349_), .Y(w_C_60_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[60]), .B(i_add1[60]), .Y(_352_) );
OR2X2 OR2X2_4 ( .A(i_add2[60]), .B(i_add1[60]), .Y(_353_) );
NAND3X1 NAND3X1_21 ( .A(_349_), .B(_353_), .C(_351_), .Y(_354_) );
NAND2X1 NAND2X1_14 ( .A(_352_), .B(_354_), .Y(w_C_61_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_51 ( .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_17 ( .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_19 ( .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_52 ( .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_5 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_6 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_22 ( .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_19 ( .A(_4_), .B(_7_), .Y(w_C_3_) );
OR2X2 OR2X2_7 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_23 ( .A(_4_), .B(_9_), .C(_7_), .Y(_10_) );
AND2X2 AND2X2_8 ( .A(_10_), .B(_8_), .Y(w_C_4_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
OR2X2 OR2X2_8 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_12_) );
NAND3X1 NAND3X1_24 ( .A(_8_), .B(_12_), .C(_10_), .Y(_13_) );
NAND2X1 NAND2X1_22 ( .A(_11_), .B(_13_), .Y(w_C_5_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_14_) );
INVX1 INVX1_53 ( .A(_14_), .Y(_15_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_16_) );
NAND3X1 NAND3X1_25 ( .A(_11_), .B(_16_), .C(_13_), .Y(_17_) );
AND2X2 AND2X2_9 ( .A(_17_), .B(_15_), .Y(w_C_6_) );
INVX1 INVX1_54 ( .A(i_add2[6]), .Y(_18_) );
INVX1 INVX1_55 ( .A(i_add1[6]), .Y(_19_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_20_) );
INVX1 INVX1_56 ( .A(_20_), .Y(_21_) );
NAND3X1 NAND3X1_26 ( .A(_15_), .B(_21_), .C(_17_), .Y(_22_) );
OAI21X1 OAI21X1_20 ( .A(_18_), .B(_19_), .C(_22_), .Y(w_C_7_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_23_) );
INVX1 INVX1_57 ( .A(_23_), .Y(_24_) );
NOR2X1 NOR2X1_25 ( .A(_18_), .B(_19_), .Y(_25_) );
INVX1 INVX1_58 ( .A(_25_), .Y(_26_) );
AND2X2 AND2X2_10 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_27_) );
INVX1 INVX1_59 ( .A(_27_), .Y(_28_) );
NAND3X1 NAND3X1_27 ( .A(_26_), .B(_28_), .C(_22_), .Y(_29_) );
AND2X2 AND2X2_11 ( .A(_29_), .B(_24_), .Y(w_C_8_) );
AND2X2 AND2X2_12 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_30_) );
INVX1 INVX1_60 ( .A(_30_), .Y(_31_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_32_) );
INVX1 INVX1_61 ( .A(_32_), .Y(_33_) );
NAND3X1 NAND3X1_28 ( .A(_24_), .B(_33_), .C(_29_), .Y(_34_) );
AND2X2 AND2X2_13 ( .A(_34_), .B(_31_), .Y(_35_) );
INVX1 INVX1_62 ( .A(_35_), .Y(w_C_9_) );
AND2X2 AND2X2_14 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_36_) );
INVX1 INVX1_63 ( .A(_36_), .Y(_37_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_38_) );
OAI21X1 OAI21X1_21 ( .A(_38_), .B(_35_), .C(_37_), .Y(w_C_10_) );
AND2X2 AND2X2_15 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_39_) );
INVX1 INVX1_64 ( .A(_39_), .Y(_40_) );
INVX1 INVX1_65 ( .A(_38_), .Y(_41_) );
NAND3X1 NAND3X1_29 ( .A(_31_), .B(_37_), .C(_34_), .Y(_42_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_43_) );
INVX1 INVX1_66 ( .A(_43_), .Y(_44_) );
NAND3X1 NAND3X1_30 ( .A(_41_), .B(_44_), .C(_42_), .Y(_45_) );
AND2X2 AND2X2_16 ( .A(_45_), .B(_40_), .Y(_46_) );
INVX1 INVX1_67 ( .A(_46_), .Y(w_C_11_) );
AND2X2 AND2X2_17 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_47_) );
INVX1 INVX1_68 ( .A(_47_), .Y(_48_) );
NAND3X1 NAND3X1_31 ( .A(_40_), .B(_48_), .C(_45_), .Y(_49_) );
OAI21X1 OAI21X1_22 ( .A(i_add2[11]), .B(i_add1[11]), .C(_49_), .Y(_50_) );
INVX1 INVX1_69 ( .A(_50_), .Y(w_C_12_) );
INVX1 INVX1_70 ( .A(i_add2[12]), .Y(_51_) );
BUFX2 BUFX2_1 ( .A(_355__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_355__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_355__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_355__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_355__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_355__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_355__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_355__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_355__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_355__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_355__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_355__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_355__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_355__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_355__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_355__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_355__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_355__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_355__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_355__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_355__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_355__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_355__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_355__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_355__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_355__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_355__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_355__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_355__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_355__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_355__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_355__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_355__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_355__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_355__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_355__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_355__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(_355__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .A(_355__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .A(_355__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .A(_355__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .A(_355__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .A(_355__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .A(_355__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .A(_355__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .A(_355__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .A(_355__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .A(_355__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .A(_355__48_), .Y(o_result[48]) );
BUFX2 BUFX2_50 ( .A(_355__49_), .Y(o_result[49]) );
BUFX2 BUFX2_51 ( .A(_355__50_), .Y(o_result[50]) );
BUFX2 BUFX2_52 ( .A(_355__51_), .Y(o_result[51]) );
BUFX2 BUFX2_53 ( .A(_355__52_), .Y(o_result[52]) );
BUFX2 BUFX2_54 ( .A(_355__53_), .Y(o_result[53]) );
BUFX2 BUFX2_55 ( .A(_355__54_), .Y(o_result[54]) );
BUFX2 BUFX2_56 ( .A(_355__55_), .Y(o_result[55]) );
BUFX2 BUFX2_57 ( .A(_355__56_), .Y(o_result[56]) );
BUFX2 BUFX2_58 ( .A(_355__57_), .Y(o_result[57]) );
BUFX2 BUFX2_59 ( .A(_355__58_), .Y(o_result[58]) );
BUFX2 BUFX2_60 ( .A(_355__59_), .Y(o_result[59]) );
BUFX2 BUFX2_61 ( .A(_355__60_), .Y(o_result[60]) );
BUFX2 BUFX2_62 ( .A(w_C_61_), .Y(o_result[61]) );
INVX1 INVX1_71 ( .A(w_C_4_), .Y(_359_) );
OR2X2 OR2X2_9 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_360_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_361_) );
NAND3X1 NAND3X1_32 ( .A(_359_), .B(_361_), .C(_360_), .Y(_362_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_356_) );
AND2X2 AND2X2_18 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_357_) );
OAI21X1 OAI21X1_23 ( .A(_356_), .B(_357_), .C(w_C_4_), .Y(_358_) );
NAND2X1 NAND2X1_25 ( .A(_358_), .B(_362_), .Y(_355__4_) );
INVX1 INVX1_72 ( .A(w_C_5_), .Y(_366_) );
OR2X2 OR2X2_10 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_367_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_368_) );
NAND3X1 NAND3X1_33 ( .A(_366_), .B(_368_), .C(_367_), .Y(_369_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_363_) );
AND2X2 AND2X2_19 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_364_) );
OAI21X1 OAI21X1_24 ( .A(_363_), .B(_364_), .C(w_C_5_), .Y(_365_) );
NAND2X1 NAND2X1_27 ( .A(_365_), .B(_369_), .Y(_355__5_) );
INVX1 INVX1_73 ( .A(w_C_6_), .Y(_373_) );
OR2X2 OR2X2_11 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_374_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_375_) );
NAND3X1 NAND3X1_34 ( .A(_373_), .B(_375_), .C(_374_), .Y(_376_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_370_) );
AND2X2 AND2X2_20 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_371_) );
OAI21X1 OAI21X1_25 ( .A(_370_), .B(_371_), .C(w_C_6_), .Y(_372_) );
NAND2X1 NAND2X1_29 ( .A(_372_), .B(_376_), .Y(_355__6_) );
INVX1 INVX1_74 ( .A(w_C_7_), .Y(_380_) );
OR2X2 OR2X2_12 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_381_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_382_) );
NAND3X1 NAND3X1_35 ( .A(_380_), .B(_382_), .C(_381_), .Y(_383_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_377_) );
AND2X2 AND2X2_21 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_378_) );
OAI21X1 OAI21X1_26 ( .A(_377_), .B(_378_), .C(w_C_7_), .Y(_379_) );
NAND2X1 NAND2X1_31 ( .A(_379_), .B(_383_), .Y(_355__7_) );
INVX1 INVX1_75 ( .A(w_C_8_), .Y(_387_) );
OR2X2 OR2X2_13 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_388_) );
NAND2X1 NAND2X1_32 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_389_) );
NAND3X1 NAND3X1_36 ( .A(_387_), .B(_389_), .C(_388_), .Y(_390_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_384_) );
AND2X2 AND2X2_22 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_385_) );
OAI21X1 OAI21X1_27 ( .A(_384_), .B(_385_), .C(w_C_8_), .Y(_386_) );
NAND2X1 NAND2X1_33 ( .A(_386_), .B(_390_), .Y(_355__8_) );
INVX1 INVX1_76 ( .A(w_C_9_), .Y(_394_) );
OR2X2 OR2X2_14 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_395_) );
NAND2X1 NAND2X1_34 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_396_) );
NAND3X1 NAND3X1_37 ( .A(_394_), .B(_396_), .C(_395_), .Y(_397_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_391_) );
AND2X2 AND2X2_23 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_392_) );
OAI21X1 OAI21X1_28 ( .A(_391_), .B(_392_), .C(w_C_9_), .Y(_393_) );
NAND2X1 NAND2X1_35 ( .A(_393_), .B(_397_), .Y(_355__9_) );
INVX1 INVX1_77 ( .A(w_C_10_), .Y(_401_) );
OR2X2 OR2X2_15 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_402_) );
NAND2X1 NAND2X1_36 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_403_) );
NAND3X1 NAND3X1_38 ( .A(_401_), .B(_403_), .C(_402_), .Y(_404_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_398_) );
AND2X2 AND2X2_24 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_399_) );
OAI21X1 OAI21X1_29 ( .A(_398_), .B(_399_), .C(w_C_10_), .Y(_400_) );
NAND2X1 NAND2X1_37 ( .A(_400_), .B(_404_), .Y(_355__10_) );
INVX1 INVX1_78 ( .A(w_C_11_), .Y(_408_) );
OR2X2 OR2X2_16 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_409_) );
NAND2X1 NAND2X1_38 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_410_) );
NAND3X1 NAND3X1_39 ( .A(_408_), .B(_410_), .C(_409_), .Y(_411_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_405_) );
AND2X2 AND2X2_25 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_406_) );
OAI21X1 OAI21X1_30 ( .A(_405_), .B(_406_), .C(w_C_11_), .Y(_407_) );
NAND2X1 NAND2X1_39 ( .A(_407_), .B(_411_), .Y(_355__11_) );
INVX1 INVX1_79 ( .A(w_C_12_), .Y(_415_) );
OR2X2 OR2X2_17 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_416_) );
NAND2X1 NAND2X1_40 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_417_) );
NAND3X1 NAND3X1_40 ( .A(_415_), .B(_417_), .C(_416_), .Y(_418_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_412_) );
AND2X2 AND2X2_26 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_413_) );
OAI21X1 OAI21X1_31 ( .A(_412_), .B(_413_), .C(w_C_12_), .Y(_414_) );
NAND2X1 NAND2X1_41 ( .A(_414_), .B(_418_), .Y(_355__12_) );
INVX1 INVX1_80 ( .A(w_C_13_), .Y(_422_) );
OR2X2 OR2X2_18 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_423_) );
NAND2X1 NAND2X1_42 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_424_) );
NAND3X1 NAND3X1_41 ( .A(_422_), .B(_424_), .C(_423_), .Y(_425_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_419_) );
AND2X2 AND2X2_27 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_420_) );
OAI21X1 OAI21X1_32 ( .A(_419_), .B(_420_), .C(w_C_13_), .Y(_421_) );
NAND2X1 NAND2X1_43 ( .A(_421_), .B(_425_), .Y(_355__13_) );
INVX1 INVX1_81 ( .A(w_C_14_), .Y(_429_) );
OR2X2 OR2X2_19 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_430_) );
NAND2X1 NAND2X1_44 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_431_) );
NAND3X1 NAND3X1_42 ( .A(_429_), .B(_431_), .C(_430_), .Y(_432_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_426_) );
AND2X2 AND2X2_28 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_427_) );
OAI21X1 OAI21X1_33 ( .A(_426_), .B(_427_), .C(w_C_14_), .Y(_428_) );
NAND2X1 NAND2X1_45 ( .A(_428_), .B(_432_), .Y(_355__14_) );
INVX1 INVX1_82 ( .A(w_C_15_), .Y(_436_) );
OR2X2 OR2X2_20 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_437_) );
NAND2X1 NAND2X1_46 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_438_) );
NAND3X1 NAND3X1_43 ( .A(_436_), .B(_438_), .C(_437_), .Y(_439_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_433_) );
AND2X2 AND2X2_29 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_434_) );
OAI21X1 OAI21X1_34 ( .A(_433_), .B(_434_), .C(w_C_15_), .Y(_435_) );
NAND2X1 NAND2X1_47 ( .A(_435_), .B(_439_), .Y(_355__15_) );
INVX1 INVX1_83 ( .A(w_C_16_), .Y(_443_) );
OR2X2 OR2X2_21 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_444_) );
NAND2X1 NAND2X1_48 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_445_) );
NAND3X1 NAND3X1_44 ( .A(_443_), .B(_445_), .C(_444_), .Y(_446_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_440_) );
AND2X2 AND2X2_30 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_441_) );
OAI21X1 OAI21X1_35 ( .A(_440_), .B(_441_), .C(w_C_16_), .Y(_442_) );
NAND2X1 NAND2X1_49 ( .A(_442_), .B(_446_), .Y(_355__16_) );
INVX1 INVX1_84 ( .A(w_C_17_), .Y(_450_) );
OR2X2 OR2X2_22 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_451_) );
NAND2X1 NAND2X1_50 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_452_) );
NAND3X1 NAND3X1_45 ( .A(_450_), .B(_452_), .C(_451_), .Y(_453_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_447_) );
AND2X2 AND2X2_31 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_448_) );
OAI21X1 OAI21X1_36 ( .A(_447_), .B(_448_), .C(w_C_17_), .Y(_449_) );
NAND2X1 NAND2X1_51 ( .A(_449_), .B(_453_), .Y(_355__17_) );
INVX1 INVX1_85 ( .A(w_C_18_), .Y(_457_) );
OR2X2 OR2X2_23 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_458_) );
NAND2X1 NAND2X1_52 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_459_) );
NAND3X1 NAND3X1_46 ( .A(_457_), .B(_459_), .C(_458_), .Y(_460_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_454_) );
AND2X2 AND2X2_32 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_455_) );
OAI21X1 OAI21X1_37 ( .A(_454_), .B(_455_), .C(w_C_18_), .Y(_456_) );
NAND2X1 NAND2X1_53 ( .A(_456_), .B(_460_), .Y(_355__18_) );
INVX1 INVX1_86 ( .A(w_C_19_), .Y(_464_) );
OR2X2 OR2X2_24 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_465_) );
NAND2X1 NAND2X1_54 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_466_) );
NAND3X1 NAND3X1_47 ( .A(_464_), .B(_466_), .C(_465_), .Y(_467_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_461_) );
AND2X2 AND2X2_33 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_462_) );
OAI21X1 OAI21X1_38 ( .A(_461_), .B(_462_), .C(w_C_19_), .Y(_463_) );
NAND2X1 NAND2X1_55 ( .A(_463_), .B(_467_), .Y(_355__19_) );
INVX1 INVX1_87 ( .A(w_C_20_), .Y(_471_) );
OR2X2 OR2X2_25 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_472_) );
NAND2X1 NAND2X1_56 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_473_) );
NAND3X1 NAND3X1_48 ( .A(_471_), .B(_473_), .C(_472_), .Y(_474_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_468_) );
AND2X2 AND2X2_34 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_469_) );
OAI21X1 OAI21X1_39 ( .A(_468_), .B(_469_), .C(w_C_20_), .Y(_470_) );
NAND2X1 NAND2X1_57 ( .A(_470_), .B(_474_), .Y(_355__20_) );
INVX1 INVX1_88 ( .A(w_C_21_), .Y(_478_) );
OR2X2 OR2X2_26 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_479_) );
NAND2X1 NAND2X1_58 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_480_) );
NAND3X1 NAND3X1_49 ( .A(_478_), .B(_480_), .C(_479_), .Y(_481_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_475_) );
AND2X2 AND2X2_35 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_476_) );
OAI21X1 OAI21X1_40 ( .A(_475_), .B(_476_), .C(w_C_21_), .Y(_477_) );
NAND2X1 NAND2X1_59 ( .A(_477_), .B(_481_), .Y(_355__21_) );
INVX1 INVX1_89 ( .A(w_C_22_), .Y(_485_) );
OR2X2 OR2X2_27 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_486_) );
NAND2X1 NAND2X1_60 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_487_) );
NAND3X1 NAND3X1_50 ( .A(_485_), .B(_487_), .C(_486_), .Y(_488_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_482_) );
AND2X2 AND2X2_36 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_483_) );
OAI21X1 OAI21X1_41 ( .A(_482_), .B(_483_), .C(w_C_22_), .Y(_484_) );
NAND2X1 NAND2X1_61 ( .A(_484_), .B(_488_), .Y(_355__22_) );
INVX1 INVX1_90 ( .A(w_C_23_), .Y(_492_) );
OR2X2 OR2X2_28 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_493_) );
NAND2X1 NAND2X1_62 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_494_) );
NAND3X1 NAND3X1_51 ( .A(_492_), .B(_494_), .C(_493_), .Y(_495_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_489_) );
AND2X2 AND2X2_37 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_490_) );
OAI21X1 OAI21X1_42 ( .A(_489_), .B(_490_), .C(w_C_23_), .Y(_491_) );
NAND2X1 NAND2X1_63 ( .A(_491_), .B(_495_), .Y(_355__23_) );
INVX1 INVX1_91 ( .A(w_C_24_), .Y(_499_) );
OR2X2 OR2X2_29 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_500_) );
NAND2X1 NAND2X1_64 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_501_) );
NAND3X1 NAND3X1_52 ( .A(_499_), .B(_501_), .C(_500_), .Y(_502_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_496_) );
AND2X2 AND2X2_38 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_497_) );
OAI21X1 OAI21X1_43 ( .A(_496_), .B(_497_), .C(w_C_24_), .Y(_498_) );
NAND2X1 NAND2X1_65 ( .A(_498_), .B(_502_), .Y(_355__24_) );
INVX1 INVX1_92 ( .A(w_C_25_), .Y(_506_) );
OR2X2 OR2X2_30 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_507_) );
NAND2X1 NAND2X1_66 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_508_) );
NAND3X1 NAND3X1_53 ( .A(_506_), .B(_508_), .C(_507_), .Y(_509_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_503_) );
AND2X2 AND2X2_39 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_504_) );
OAI21X1 OAI21X1_44 ( .A(_503_), .B(_504_), .C(w_C_25_), .Y(_505_) );
NAND2X1 NAND2X1_67 ( .A(_505_), .B(_509_), .Y(_355__25_) );
INVX1 INVX1_93 ( .A(w_C_26_), .Y(_513_) );
OR2X2 OR2X2_31 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_514_) );
NAND2X1 NAND2X1_68 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_515_) );
NAND3X1 NAND3X1_54 ( .A(_513_), .B(_515_), .C(_514_), .Y(_516_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_510_) );
AND2X2 AND2X2_40 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_511_) );
OAI21X1 OAI21X1_45 ( .A(_510_), .B(_511_), .C(w_C_26_), .Y(_512_) );
NAND2X1 NAND2X1_69 ( .A(_512_), .B(_516_), .Y(_355__26_) );
INVX1 INVX1_94 ( .A(w_C_27_), .Y(_520_) );
OR2X2 OR2X2_32 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_521_) );
NAND2X1 NAND2X1_70 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_522_) );
NAND3X1 NAND3X1_55 ( .A(_520_), .B(_522_), .C(_521_), .Y(_523_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_517_) );
AND2X2 AND2X2_41 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_518_) );
OAI21X1 OAI21X1_46 ( .A(_517_), .B(_518_), .C(w_C_27_), .Y(_519_) );
NAND2X1 NAND2X1_71 ( .A(_519_), .B(_523_), .Y(_355__27_) );
INVX1 INVX1_95 ( .A(w_C_28_), .Y(_527_) );
OR2X2 OR2X2_33 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_528_) );
NAND2X1 NAND2X1_72 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_529_) );
NAND3X1 NAND3X1_56 ( .A(_527_), .B(_529_), .C(_528_), .Y(_530_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_524_) );
AND2X2 AND2X2_42 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_525_) );
OAI21X1 OAI21X1_47 ( .A(_524_), .B(_525_), .C(w_C_28_), .Y(_526_) );
NAND2X1 NAND2X1_73 ( .A(_526_), .B(_530_), .Y(_355__28_) );
INVX1 INVX1_96 ( .A(w_C_29_), .Y(_534_) );
OR2X2 OR2X2_34 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_535_) );
NAND2X1 NAND2X1_74 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_536_) );
NAND3X1 NAND3X1_57 ( .A(_534_), .B(_536_), .C(_535_), .Y(_537_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_531_) );
AND2X2 AND2X2_43 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_532_) );
OAI21X1 OAI21X1_48 ( .A(_531_), .B(_532_), .C(w_C_29_), .Y(_533_) );
NAND2X1 NAND2X1_75 ( .A(_533_), .B(_537_), .Y(_355__29_) );
INVX1 INVX1_97 ( .A(w_C_30_), .Y(_541_) );
OR2X2 OR2X2_35 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_542_) );
NAND2X1 NAND2X1_76 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_543_) );
NAND3X1 NAND3X1_58 ( .A(_541_), .B(_543_), .C(_542_), .Y(_544_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_538_) );
AND2X2 AND2X2_44 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_539_) );
OAI21X1 OAI21X1_49 ( .A(_538_), .B(_539_), .C(w_C_30_), .Y(_540_) );
NAND2X1 NAND2X1_77 ( .A(_540_), .B(_544_), .Y(_355__30_) );
INVX1 INVX1_98 ( .A(w_C_31_), .Y(_548_) );
OR2X2 OR2X2_36 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_549_) );
NAND2X1 NAND2X1_78 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_550_) );
NAND3X1 NAND3X1_59 ( .A(_548_), .B(_550_), .C(_549_), .Y(_551_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_545_) );
AND2X2 AND2X2_45 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_546_) );
OAI21X1 OAI21X1_50 ( .A(_545_), .B(_546_), .C(w_C_31_), .Y(_547_) );
NAND2X1 NAND2X1_79 ( .A(_547_), .B(_551_), .Y(_355__31_) );
INVX1 INVX1_99 ( .A(w_C_32_), .Y(_555_) );
OR2X2 OR2X2_37 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_556_) );
NAND2X1 NAND2X1_80 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_557_) );
NAND3X1 NAND3X1_60 ( .A(_555_), .B(_557_), .C(_556_), .Y(_558_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_552_) );
AND2X2 AND2X2_46 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_553_) );
OAI21X1 OAI21X1_51 ( .A(_552_), .B(_553_), .C(w_C_32_), .Y(_554_) );
NAND2X1 NAND2X1_81 ( .A(_554_), .B(_558_), .Y(_355__32_) );
INVX1 INVX1_100 ( .A(w_C_33_), .Y(_562_) );
OR2X2 OR2X2_38 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_563_) );
NAND2X1 NAND2X1_82 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_564_) );
NAND3X1 NAND3X1_61 ( .A(_562_), .B(_564_), .C(_563_), .Y(_565_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_559_) );
AND2X2 AND2X2_47 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_560_) );
OAI21X1 OAI21X1_52 ( .A(_559_), .B(_560_), .C(w_C_33_), .Y(_561_) );
NAND2X1 NAND2X1_83 ( .A(_561_), .B(_565_), .Y(_355__33_) );
INVX1 INVX1_101 ( .A(w_C_34_), .Y(_569_) );
OR2X2 OR2X2_39 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_570_) );
NAND2X1 NAND2X1_84 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_571_) );
NAND3X1 NAND3X1_62 ( .A(_569_), .B(_571_), .C(_570_), .Y(_572_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_566_) );
AND2X2 AND2X2_48 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_567_) );
OAI21X1 OAI21X1_53 ( .A(_566_), .B(_567_), .C(w_C_34_), .Y(_568_) );
NAND2X1 NAND2X1_85 ( .A(_568_), .B(_572_), .Y(_355__34_) );
INVX1 INVX1_102 ( .A(w_C_35_), .Y(_576_) );
OR2X2 OR2X2_40 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_577_) );
NAND2X1 NAND2X1_86 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_578_) );
NAND3X1 NAND3X1_63 ( .A(_576_), .B(_578_), .C(_577_), .Y(_579_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_573_) );
AND2X2 AND2X2_49 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_574_) );
OAI21X1 OAI21X1_54 ( .A(_573_), .B(_574_), .C(w_C_35_), .Y(_575_) );
NAND2X1 NAND2X1_87 ( .A(_575_), .B(_579_), .Y(_355__35_) );
INVX1 INVX1_103 ( .A(w_C_36_), .Y(_583_) );
OR2X2 OR2X2_41 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_584_) );
NAND2X1 NAND2X1_88 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_585_) );
NAND3X1 NAND3X1_64 ( .A(_583_), .B(_585_), .C(_584_), .Y(_586_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_580_) );
AND2X2 AND2X2_50 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_581_) );
OAI21X1 OAI21X1_55 ( .A(_580_), .B(_581_), .C(w_C_36_), .Y(_582_) );
NAND2X1 NAND2X1_89 ( .A(_582_), .B(_586_), .Y(_355__36_) );
INVX1 INVX1_104 ( .A(w_C_37_), .Y(_590_) );
OR2X2 OR2X2_42 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_591_) );
NAND2X1 NAND2X1_90 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_592_) );
NAND3X1 NAND3X1_65 ( .A(_590_), .B(_592_), .C(_591_), .Y(_593_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_587_) );
AND2X2 AND2X2_51 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_588_) );
OAI21X1 OAI21X1_56 ( .A(_587_), .B(_588_), .C(w_C_37_), .Y(_589_) );
NAND2X1 NAND2X1_91 ( .A(_589_), .B(_593_), .Y(_355__37_) );
INVX1 INVX1_105 ( .A(w_C_38_), .Y(_597_) );
OR2X2 OR2X2_43 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_598_) );
NAND2X1 NAND2X1_92 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_599_) );
NAND3X1 NAND3X1_66 ( .A(_597_), .B(_599_), .C(_598_), .Y(_600_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_594_) );
AND2X2 AND2X2_52 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_595_) );
OAI21X1 OAI21X1_57 ( .A(_594_), .B(_595_), .C(w_C_38_), .Y(_596_) );
NAND2X1 NAND2X1_93 ( .A(_596_), .B(_600_), .Y(_355__38_) );
INVX1 INVX1_106 ( .A(w_C_39_), .Y(_604_) );
OR2X2 OR2X2_44 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_605_) );
NAND2X1 NAND2X1_94 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_606_) );
NAND3X1 NAND3X1_67 ( .A(_604_), .B(_606_), .C(_605_), .Y(_607_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_601_) );
AND2X2 AND2X2_53 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_602_) );
OAI21X1 OAI21X1_58 ( .A(_601_), .B(_602_), .C(w_C_39_), .Y(_603_) );
NAND2X1 NAND2X1_95 ( .A(_603_), .B(_607_), .Y(_355__39_) );
INVX1 INVX1_107 ( .A(w_C_40_), .Y(_611_) );
OR2X2 OR2X2_45 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_612_) );
NAND2X1 NAND2X1_96 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_613_) );
NAND3X1 NAND3X1_68 ( .A(_611_), .B(_613_), .C(_612_), .Y(_614_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_608_) );
AND2X2 AND2X2_54 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_609_) );
OAI21X1 OAI21X1_59 ( .A(_608_), .B(_609_), .C(w_C_40_), .Y(_610_) );
NAND2X1 NAND2X1_97 ( .A(_610_), .B(_614_), .Y(_355__40_) );
INVX1 INVX1_108 ( .A(w_C_41_), .Y(_618_) );
OR2X2 OR2X2_46 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_619_) );
NAND2X1 NAND2X1_98 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_620_) );
NAND3X1 NAND3X1_69 ( .A(_618_), .B(_620_), .C(_619_), .Y(_621_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_615_) );
AND2X2 AND2X2_55 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_616_) );
OAI21X1 OAI21X1_60 ( .A(_615_), .B(_616_), .C(w_C_41_), .Y(_617_) );
NAND2X1 NAND2X1_99 ( .A(_617_), .B(_621_), .Y(_355__41_) );
INVX1 INVX1_109 ( .A(w_C_42_), .Y(_625_) );
OR2X2 OR2X2_47 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_626_) );
NAND2X1 NAND2X1_100 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_627_) );
NAND3X1 NAND3X1_70 ( .A(_625_), .B(_627_), .C(_626_), .Y(_628_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_622_) );
AND2X2 AND2X2_56 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_623_) );
OAI21X1 OAI21X1_61 ( .A(_622_), .B(_623_), .C(w_C_42_), .Y(_624_) );
NAND2X1 NAND2X1_101 ( .A(_624_), .B(_628_), .Y(_355__42_) );
INVX1 INVX1_110 ( .A(w_C_43_), .Y(_632_) );
OR2X2 OR2X2_48 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_633_) );
NAND2X1 NAND2X1_102 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_634_) );
NAND3X1 NAND3X1_71 ( .A(_632_), .B(_634_), .C(_633_), .Y(_635_) );
NOR2X1 NOR2X1_68 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_629_) );
AND2X2 AND2X2_57 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_630_) );
OAI21X1 OAI21X1_62 ( .A(_629_), .B(_630_), .C(w_C_43_), .Y(_631_) );
NAND2X1 NAND2X1_103 ( .A(_631_), .B(_635_), .Y(_355__43_) );
INVX1 INVX1_111 ( .A(w_C_44_), .Y(_639_) );
OR2X2 OR2X2_49 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_640_) );
NAND2X1 NAND2X1_104 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_641_) );
NAND3X1 NAND3X1_72 ( .A(_639_), .B(_641_), .C(_640_), .Y(_642_) );
NOR2X1 NOR2X1_69 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_636_) );
AND2X2 AND2X2_58 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_637_) );
OAI21X1 OAI21X1_63 ( .A(_636_), .B(_637_), .C(w_C_44_), .Y(_638_) );
NAND2X1 NAND2X1_105 ( .A(_638_), .B(_642_), .Y(_355__44_) );
INVX1 INVX1_112 ( .A(w_C_45_), .Y(_646_) );
OR2X2 OR2X2_50 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_647_) );
NAND2X1 NAND2X1_106 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_648_) );
NAND3X1 NAND3X1_73 ( .A(_646_), .B(_648_), .C(_647_), .Y(_649_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_643_) );
AND2X2 AND2X2_59 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_644_) );
OAI21X1 OAI21X1_64 ( .A(_643_), .B(_644_), .C(w_C_45_), .Y(_645_) );
NAND2X1 NAND2X1_107 ( .A(_645_), .B(_649_), .Y(_355__45_) );
INVX1 INVX1_113 ( .A(w_C_46_), .Y(_653_) );
OR2X2 OR2X2_51 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_654_) );
NAND2X1 NAND2X1_108 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_655_) );
NAND3X1 NAND3X1_74 ( .A(_653_), .B(_655_), .C(_654_), .Y(_656_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_650_) );
AND2X2 AND2X2_60 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_651_) );
OAI21X1 OAI21X1_65 ( .A(_650_), .B(_651_), .C(w_C_46_), .Y(_652_) );
NAND2X1 NAND2X1_109 ( .A(_652_), .B(_656_), .Y(_355__46_) );
INVX1 INVX1_114 ( .A(w_C_47_), .Y(_660_) );
OR2X2 OR2X2_52 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_661_) );
NAND2X1 NAND2X1_110 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_662_) );
NAND3X1 NAND3X1_75 ( .A(_660_), .B(_662_), .C(_661_), .Y(_663_) );
NOR2X1 NOR2X1_72 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_657_) );
AND2X2 AND2X2_61 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_658_) );
OAI21X1 OAI21X1_66 ( .A(_657_), .B(_658_), .C(w_C_47_), .Y(_659_) );
NAND2X1 NAND2X1_111 ( .A(_659_), .B(_663_), .Y(_355__47_) );
INVX1 INVX1_115 ( .A(w_C_48_), .Y(_667_) );
OR2X2 OR2X2_53 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_668_) );
NAND2X1 NAND2X1_112 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_669_) );
NAND3X1 NAND3X1_76 ( .A(_667_), .B(_669_), .C(_668_), .Y(_670_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_664_) );
AND2X2 AND2X2_62 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_665_) );
OAI21X1 OAI21X1_67 ( .A(_664_), .B(_665_), .C(w_C_48_), .Y(_666_) );
NAND2X1 NAND2X1_113 ( .A(_666_), .B(_670_), .Y(_355__48_) );
INVX1 INVX1_116 ( .A(w_C_49_), .Y(_674_) );
OR2X2 OR2X2_54 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_675_) );
NAND2X1 NAND2X1_114 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_676_) );
NAND3X1 NAND3X1_77 ( .A(_674_), .B(_676_), .C(_675_), .Y(_677_) );
NOR2X1 NOR2X1_74 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_671_) );
AND2X2 AND2X2_63 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_672_) );
OAI21X1 OAI21X1_68 ( .A(_671_), .B(_672_), .C(w_C_49_), .Y(_673_) );
NAND2X1 NAND2X1_115 ( .A(_673_), .B(_677_), .Y(_355__49_) );
INVX1 INVX1_117 ( .A(w_C_50_), .Y(_681_) );
OR2X2 OR2X2_55 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_682_) );
NAND2X1 NAND2X1_116 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_683_) );
NAND3X1 NAND3X1_78 ( .A(_681_), .B(_683_), .C(_682_), .Y(_684_) );
NOR2X1 NOR2X1_75 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_678_) );
AND2X2 AND2X2_64 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_679_) );
OAI21X1 OAI21X1_69 ( .A(_678_), .B(_679_), .C(w_C_50_), .Y(_680_) );
NAND2X1 NAND2X1_117 ( .A(_680_), .B(_684_), .Y(_355__50_) );
INVX1 INVX1_118 ( .A(w_C_51_), .Y(_688_) );
OR2X2 OR2X2_56 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_689_) );
NAND2X1 NAND2X1_118 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_690_) );
NAND3X1 NAND3X1_79 ( .A(_688_), .B(_690_), .C(_689_), .Y(_691_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_685_) );
AND2X2 AND2X2_65 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_686_) );
OAI21X1 OAI21X1_70 ( .A(_685_), .B(_686_), .C(w_C_51_), .Y(_687_) );
NAND2X1 NAND2X1_119 ( .A(_687_), .B(_691_), .Y(_355__51_) );
INVX1 INVX1_119 ( .A(w_C_52_), .Y(_695_) );
OR2X2 OR2X2_57 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_696_) );
NAND2X1 NAND2X1_120 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_697_) );
NAND3X1 NAND3X1_80 ( .A(_695_), .B(_697_), .C(_696_), .Y(_698_) );
NOR2X1 NOR2X1_77 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_692_) );
AND2X2 AND2X2_66 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_693_) );
OAI21X1 OAI21X1_71 ( .A(_692_), .B(_693_), .C(w_C_52_), .Y(_694_) );
NAND2X1 NAND2X1_121 ( .A(_694_), .B(_698_), .Y(_355__52_) );
INVX1 INVX1_120 ( .A(w_C_53_), .Y(_702_) );
OR2X2 OR2X2_58 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_703_) );
NAND2X1 NAND2X1_122 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_704_) );
NAND3X1 NAND3X1_81 ( .A(_702_), .B(_704_), .C(_703_), .Y(_705_) );
NOR2X1 NOR2X1_78 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_699_) );
AND2X2 AND2X2_67 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_700_) );
OAI21X1 OAI21X1_72 ( .A(_699_), .B(_700_), .C(w_C_53_), .Y(_701_) );
NAND2X1 NAND2X1_123 ( .A(_701_), .B(_705_), .Y(_355__53_) );
INVX1 INVX1_121 ( .A(w_C_54_), .Y(_709_) );
OR2X2 OR2X2_59 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_710_) );
NAND2X1 NAND2X1_124 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_711_) );
NAND3X1 NAND3X1_82 ( .A(_709_), .B(_711_), .C(_710_), .Y(_712_) );
NOR2X1 NOR2X1_79 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_706_) );
AND2X2 AND2X2_68 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_707_) );
OAI21X1 OAI21X1_73 ( .A(_706_), .B(_707_), .C(w_C_54_), .Y(_708_) );
NAND2X1 NAND2X1_125 ( .A(_708_), .B(_712_), .Y(_355__54_) );
INVX1 INVX1_122 ( .A(w_C_55_), .Y(_716_) );
OR2X2 OR2X2_60 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_717_) );
NAND2X1 NAND2X1_126 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_718_) );
NAND3X1 NAND3X1_83 ( .A(_716_), .B(_718_), .C(_717_), .Y(_719_) );
NOR2X1 NOR2X1_80 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_713_) );
AND2X2 AND2X2_69 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_714_) );
OAI21X1 OAI21X1_74 ( .A(_713_), .B(_714_), .C(w_C_55_), .Y(_715_) );
NAND2X1 NAND2X1_127 ( .A(_715_), .B(_719_), .Y(_355__55_) );
INVX1 INVX1_123 ( .A(w_C_56_), .Y(_723_) );
OR2X2 OR2X2_61 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_724_) );
NAND2X1 NAND2X1_128 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_725_) );
NAND3X1 NAND3X1_84 ( .A(_723_), .B(_725_), .C(_724_), .Y(_726_) );
NOR2X1 NOR2X1_81 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_720_) );
AND2X2 AND2X2_70 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_721_) );
OAI21X1 OAI21X1_75 ( .A(_720_), .B(_721_), .C(w_C_56_), .Y(_722_) );
NAND2X1 NAND2X1_129 ( .A(_722_), .B(_726_), .Y(_355__56_) );
INVX1 INVX1_124 ( .A(w_C_57_), .Y(_730_) );
OR2X2 OR2X2_62 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_731_) );
NAND2X1 NAND2X1_130 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_732_) );
NAND3X1 NAND3X1_85 ( .A(_730_), .B(_732_), .C(_731_), .Y(_733_) );
NOR2X1 NOR2X1_82 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_727_) );
AND2X2 AND2X2_71 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_728_) );
OAI21X1 OAI21X1_76 ( .A(_727_), .B(_728_), .C(w_C_57_), .Y(_729_) );
NAND2X1 NAND2X1_131 ( .A(_729_), .B(_733_), .Y(_355__57_) );
INVX1 INVX1_125 ( .A(w_C_58_), .Y(_737_) );
OR2X2 OR2X2_63 ( .A(i_add2[58]), .B(i_add1[58]), .Y(_738_) );
NAND2X1 NAND2X1_132 ( .A(i_add2[58]), .B(i_add1[58]), .Y(_739_) );
NAND3X1 NAND3X1_86 ( .A(_737_), .B(_739_), .C(_738_), .Y(_740_) );
NOR2X1 NOR2X1_83 ( .A(i_add2[58]), .B(i_add1[58]), .Y(_734_) );
AND2X2 AND2X2_72 ( .A(i_add2[58]), .B(i_add1[58]), .Y(_735_) );
OAI21X1 OAI21X1_77 ( .A(_734_), .B(_735_), .C(w_C_58_), .Y(_736_) );
NAND2X1 NAND2X1_133 ( .A(_736_), .B(_740_), .Y(_355__58_) );
INVX1 INVX1_126 ( .A(w_C_59_), .Y(_744_) );
OR2X2 OR2X2_64 ( .A(i_add2[59]), .B(i_add1[59]), .Y(_745_) );
NAND2X1 NAND2X1_134 ( .A(i_add2[59]), .B(i_add1[59]), .Y(_746_) );
NAND3X1 NAND3X1_87 ( .A(_744_), .B(_746_), .C(_745_), .Y(_747_) );
NOR2X1 NOR2X1_84 ( .A(i_add2[59]), .B(i_add1[59]), .Y(_741_) );
AND2X2 AND2X2_73 ( .A(i_add2[59]), .B(i_add1[59]), .Y(_742_) );
OAI21X1 OAI21X1_78 ( .A(_741_), .B(_742_), .C(w_C_59_), .Y(_743_) );
NAND2X1 NAND2X1_135 ( .A(_743_), .B(_747_), .Y(_355__59_) );
INVX1 INVX1_127 ( .A(w_C_60_), .Y(_751_) );
OR2X2 OR2X2_65 ( .A(i_add2[60]), .B(i_add1[60]), .Y(_752_) );
NAND2X1 NAND2X1_136 ( .A(i_add2[60]), .B(i_add1[60]), .Y(_753_) );
NAND3X1 NAND3X1_88 ( .A(_751_), .B(_753_), .C(_752_), .Y(_754_) );
NOR2X1 NOR2X1_85 ( .A(i_add2[60]), .B(i_add1[60]), .Y(_748_) );
AND2X2 AND2X2_74 ( .A(i_add2[60]), .B(i_add1[60]), .Y(_749_) );
OAI21X1 OAI21X1_79 ( .A(_748_), .B(_749_), .C(w_C_60_), .Y(_750_) );
NAND2X1 NAND2X1_137 ( .A(_750_), .B(_754_), .Y(_355__60_) );
INVX1 INVX1_128 ( .A(gnd), .Y(_758_) );
OR2X2 OR2X2_66 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_759_) );
NAND2X1 NAND2X1_138 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_760_) );
NAND3X1 NAND3X1_89 ( .A(_758_), .B(_760_), .C(_759_), .Y(_761_) );
NOR2X1 NOR2X1_86 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_755_) );
AND2X2 AND2X2_75 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_756_) );
OAI21X1 OAI21X1_80 ( .A(_755_), .B(_756_), .C(gnd), .Y(_757_) );
NAND2X1 NAND2X1_139 ( .A(_757_), .B(_761_), .Y(_355__0_) );
INVX1 INVX1_129 ( .A(w_C_1_), .Y(_765_) );
OR2X2 OR2X2_67 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_766_) );
NAND2X1 NAND2X1_140 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_767_) );
NAND3X1 NAND3X1_90 ( .A(_765_), .B(_767_), .C(_766_), .Y(_768_) );
NOR2X1 NOR2X1_87 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_762_) );
AND2X2 AND2X2_76 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_763_) );
OAI21X1 OAI21X1_81 ( .A(_762_), .B(_763_), .C(w_C_1_), .Y(_764_) );
NAND2X1 NAND2X1_141 ( .A(_764_), .B(_768_), .Y(_355__1_) );
INVX1 INVX1_130 ( .A(w_C_2_), .Y(_772_) );
OR2X2 OR2X2_68 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_773_) );
NAND2X1 NAND2X1_142 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_774_) );
NAND3X1 NAND3X1_91 ( .A(_772_), .B(_774_), .C(_773_), .Y(_775_) );
NOR2X1 NOR2X1_88 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_769_) );
AND2X2 AND2X2_77 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_770_) );
OAI21X1 OAI21X1_82 ( .A(_769_), .B(_770_), .C(w_C_2_), .Y(_771_) );
NAND2X1 NAND2X1_143 ( .A(_771_), .B(_775_), .Y(_355__2_) );
INVX1 INVX1_131 ( .A(w_C_3_), .Y(_779_) );
OR2X2 OR2X2_69 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_780_) );
NAND2X1 NAND2X1_144 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_781_) );
NAND3X1 NAND3X1_92 ( .A(_779_), .B(_781_), .C(_780_), .Y(_782_) );
NOR2X1 NOR2X1_89 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_776_) );
AND2X2 AND2X2_78 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_777_) );
OAI21X1 OAI21X1_83 ( .A(_776_), .B(_777_), .C(w_C_3_), .Y(_778_) );
NAND2X1 NAND2X1_145 ( .A(_778_), .B(_782_), .Y(_355__3_) );
INVX1 INVX1_132 ( .A(i_add1[12]), .Y(_52_) );
NOR2X1 NOR2X1_90 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_53_) );
INVX1 INVX1_133 ( .A(_53_), .Y(_54_) );
NOR2X1 NOR2X1_91 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_55_) );
INVX1 INVX1_134 ( .A(_55_), .Y(_56_) );
NAND3X1 NAND3X1_93 ( .A(_54_), .B(_56_), .C(_49_), .Y(_57_) );
OAI21X1 OAI21X1_84 ( .A(_51_), .B(_52_), .C(_57_), .Y(w_C_13_) );
NOR2X1 NOR2X1_92 ( .A(_51_), .B(_52_), .Y(_58_) );
INVX1 INVX1_135 ( .A(_58_), .Y(_59_) );
AND2X2 AND2X2_79 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_60_) );
INVX1 INVX1_136 ( .A(_60_), .Y(_61_) );
NAND3X1 NAND3X1_94 ( .A(_59_), .B(_61_), .C(_57_), .Y(_62_) );
OAI21X1 OAI21X1_85 ( .A(i_add2[13]), .B(i_add1[13]), .C(_62_), .Y(_63_) );
INVX1 INVX1_137 ( .A(_63_), .Y(w_C_14_) );
INVX1 INVX1_138 ( .A(i_add2[14]), .Y(_64_) );
INVX1 INVX1_139 ( .A(i_add1[14]), .Y(_65_) );
NOR2X1 NOR2X1_93 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_66_) );
INVX1 INVX1_140 ( .A(_66_), .Y(_67_) );
NOR2X1 NOR2X1_94 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_68_) );
INVX1 INVX1_141 ( .A(_68_), .Y(_69_) );
NAND3X1 NAND3X1_95 ( .A(_67_), .B(_69_), .C(_62_), .Y(_70_) );
OAI21X1 OAI21X1_86 ( .A(_64_), .B(_65_), .C(_70_), .Y(w_C_15_) );
NOR2X1 NOR2X1_95 ( .A(_64_), .B(_65_), .Y(_71_) );
INVX1 INVX1_142 ( .A(_71_), .Y(_72_) );
AND2X2 AND2X2_80 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_73_) );
INVX1 INVX1_143 ( .A(_73_), .Y(_74_) );
NAND3X1 NAND3X1_96 ( .A(_72_), .B(_74_), .C(_70_), .Y(_75_) );
OAI21X1 OAI21X1_87 ( .A(i_add2[15]), .B(i_add1[15]), .C(_75_), .Y(_76_) );
INVX1 INVX1_144 ( .A(_76_), .Y(w_C_16_) );
INVX1 INVX1_145 ( .A(i_add2[16]), .Y(_77_) );
INVX1 INVX1_146 ( .A(i_add1[16]), .Y(_78_) );
NOR2X1 NOR2X1_96 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_79_) );
INVX1 INVX1_147 ( .A(_79_), .Y(_80_) );
NOR2X1 NOR2X1_97 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_81_) );
INVX1 INVX1_148 ( .A(_81_), .Y(_82_) );
NAND3X1 NAND3X1_97 ( .A(_80_), .B(_82_), .C(_75_), .Y(_83_) );
OAI21X1 OAI21X1_88 ( .A(_77_), .B(_78_), .C(_83_), .Y(w_C_17_) );
NOR2X1 NOR2X1_98 ( .A(_77_), .B(_78_), .Y(_84_) );
INVX1 INVX1_149 ( .A(_84_), .Y(_85_) );
AND2X2 AND2X2_81 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_86_) );
INVX1 INVX1_150 ( .A(_86_), .Y(_87_) );
NAND3X1 NAND3X1_98 ( .A(_85_), .B(_87_), .C(_83_), .Y(_88_) );
OAI21X1 OAI21X1_89 ( .A(i_add2[17]), .B(i_add1[17]), .C(_88_), .Y(_89_) );
INVX1 INVX1_151 ( .A(_89_), .Y(w_C_18_) );
INVX1 INVX1_152 ( .A(i_add2[18]), .Y(_90_) );
INVX1 INVX1_153 ( .A(i_add1[18]), .Y(_91_) );
NOR2X1 NOR2X1_99 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_92_) );
INVX1 INVX1_154 ( .A(_92_), .Y(_93_) );
NOR2X1 NOR2X1_100 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_94_) );
INVX1 INVX1_155 ( .A(_94_), .Y(_95_) );
NAND3X1 NAND3X1_99 ( .A(_93_), .B(_95_), .C(_88_), .Y(_96_) );
OAI21X1 OAI21X1_90 ( .A(_90_), .B(_91_), .C(_96_), .Y(w_C_19_) );
NOR2X1 NOR2X1_101 ( .A(_90_), .B(_91_), .Y(_97_) );
INVX1 INVX1_156 ( .A(_97_), .Y(_98_) );
AND2X2 AND2X2_82 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_99_) );
INVX1 INVX1_157 ( .A(_99_), .Y(_100_) );
NAND3X1 NAND3X1_100 ( .A(_98_), .B(_100_), .C(_96_), .Y(_101_) );
OAI21X1 OAI21X1_91 ( .A(i_add2[19]), .B(i_add1[19]), .C(_101_), .Y(_102_) );
INVX1 INVX1_158 ( .A(_102_), .Y(w_C_20_) );
INVX1 INVX1_159 ( .A(i_add2[20]), .Y(_103_) );
INVX1 INVX1_160 ( .A(i_add1[20]), .Y(_104_) );
NOR2X1 NOR2X1_102 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_105_) );
INVX1 INVX1_161 ( .A(_105_), .Y(_106_) );
NOR2X1 NOR2X1_103 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_107_) );
INVX1 INVX1_162 ( .A(_107_), .Y(_108_) );
NAND3X1 NAND3X1_101 ( .A(_106_), .B(_108_), .C(_101_), .Y(_109_) );
OAI21X1 OAI21X1_92 ( .A(_103_), .B(_104_), .C(_109_), .Y(w_C_21_) );
NOR2X1 NOR2X1_104 ( .A(_103_), .B(_104_), .Y(_110_) );
INVX1 INVX1_163 ( .A(_110_), .Y(_111_) );
AND2X2 AND2X2_83 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_112_) );
INVX1 INVX1_164 ( .A(_112_), .Y(_113_) );
NAND3X1 NAND3X1_102 ( .A(_111_), .B(_113_), .C(_109_), .Y(_114_) );
OAI21X1 OAI21X1_93 ( .A(i_add2[21]), .B(i_add1[21]), .C(_114_), .Y(_115_) );
INVX1 INVX1_165 ( .A(_115_), .Y(w_C_22_) );
INVX1 INVX1_166 ( .A(i_add2[22]), .Y(_116_) );
INVX1 INVX1_167 ( .A(i_add1[22]), .Y(_117_) );
NOR2X1 NOR2X1_105 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_118_) );
INVX1 INVX1_168 ( .A(_118_), .Y(_119_) );
NOR2X1 NOR2X1_106 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_120_) );
INVX1 INVX1_169 ( .A(_120_), .Y(_121_) );
NAND3X1 NAND3X1_103 ( .A(_119_), .B(_121_), .C(_114_), .Y(_122_) );
OAI21X1 OAI21X1_94 ( .A(_116_), .B(_117_), .C(_122_), .Y(w_C_23_) );
NOR2X1 NOR2X1_107 ( .A(_116_), .B(_117_), .Y(_123_) );
INVX1 INVX1_170 ( .A(_123_), .Y(_124_) );
AND2X2 AND2X2_84 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_125_) );
INVX1 INVX1_171 ( .A(_125_), .Y(_126_) );
NAND3X1 NAND3X1_104 ( .A(_124_), .B(_126_), .C(_122_), .Y(_127_) );
OAI21X1 OAI21X1_95 ( .A(i_add2[23]), .B(i_add1[23]), .C(_127_), .Y(_128_) );
INVX1 INVX1_172 ( .A(_128_), .Y(w_C_24_) );
INVX1 INVX1_173 ( .A(i_add2[24]), .Y(_129_) );
INVX1 INVX1_174 ( .A(i_add1[24]), .Y(_130_) );
NOR2X1 NOR2X1_108 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_131_) );
INVX1 INVX1_175 ( .A(_131_), .Y(_132_) );
NOR2X1 NOR2X1_109 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_133_) );
INVX1 INVX1_176 ( .A(_133_), .Y(_134_) );
NAND3X1 NAND3X1_105 ( .A(_132_), .B(_134_), .C(_127_), .Y(_135_) );
OAI21X1 OAI21X1_96 ( .A(_129_), .B(_130_), .C(_135_), .Y(w_C_25_) );
NOR2X1 NOR2X1_110 ( .A(_129_), .B(_130_), .Y(_136_) );
INVX1 INVX1_177 ( .A(_136_), .Y(_137_) );
AND2X2 AND2X2_85 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_138_) );
INVX1 INVX1_178 ( .A(_138_), .Y(_139_) );
NAND3X1 NAND3X1_106 ( .A(_137_), .B(_139_), .C(_135_), .Y(_140_) );
OAI21X1 OAI21X1_97 ( .A(i_add2[25]), .B(i_add1[25]), .C(_140_), .Y(_141_) );
INVX1 INVX1_179 ( .A(_141_), .Y(w_C_26_) );
INVX1 INVX1_180 ( .A(i_add2[26]), .Y(_142_) );
INVX1 INVX1_181 ( .A(i_add1[26]), .Y(_143_) );
NOR2X1 NOR2X1_111 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_144_) );
INVX1 INVX1_182 ( .A(_144_), .Y(_145_) );
NOR2X1 NOR2X1_112 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_146_) );
INVX1 INVX1_183 ( .A(_146_), .Y(_147_) );
NAND3X1 NAND3X1_107 ( .A(_145_), .B(_147_), .C(_140_), .Y(_148_) );
OAI21X1 OAI21X1_98 ( .A(_142_), .B(_143_), .C(_148_), .Y(w_C_27_) );
NOR2X1 NOR2X1_113 ( .A(_142_), .B(_143_), .Y(_149_) );
INVX1 INVX1_184 ( .A(_149_), .Y(_150_) );
AND2X2 AND2X2_86 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_151_) );
INVX1 INVX1_185 ( .A(_151_), .Y(_152_) );
NAND3X1 NAND3X1_108 ( .A(_150_), .B(_152_), .C(_148_), .Y(_153_) );
OAI21X1 OAI21X1_99 ( .A(i_add2[27]), .B(i_add1[27]), .C(_153_), .Y(_154_) );
INVX1 INVX1_186 ( .A(_154_), .Y(w_C_28_) );
INVX1 INVX1_187 ( .A(i_add2[28]), .Y(_155_) );
INVX1 INVX1_188 ( .A(i_add1[28]), .Y(_156_) );
NOR2X1 NOR2X1_114 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_157_) );
INVX1 INVX1_189 ( .A(_157_), .Y(_158_) );
NOR2X1 NOR2X1_115 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_159_) );
INVX1 INVX1_190 ( .A(_159_), .Y(_160_) );
NAND3X1 NAND3X1_109 ( .A(_158_), .B(_160_), .C(_153_), .Y(_161_) );
OAI21X1 OAI21X1_100 ( .A(_155_), .B(_156_), .C(_161_), .Y(w_C_29_) );
NOR2X1 NOR2X1_116 ( .A(_155_), .B(_156_), .Y(_162_) );
INVX1 INVX1_191 ( .A(_162_), .Y(_163_) );
AND2X2 AND2X2_87 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_164_) );
INVX1 INVX1_192 ( .A(_164_), .Y(_165_) );
NAND3X1 NAND3X1_110 ( .A(_163_), .B(_165_), .C(_161_), .Y(_166_) );
OAI21X1 OAI21X1_101 ( .A(i_add2[29]), .B(i_add1[29]), .C(_166_), .Y(_167_) );
INVX1 INVX1_193 ( .A(_167_), .Y(w_C_30_) );
INVX1 INVX1_194 ( .A(i_add2[30]), .Y(_168_) );
INVX1 INVX1_195 ( .A(i_add1[30]), .Y(_169_) );
NOR2X1 NOR2X1_117 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_170_) );
INVX1 INVX1_196 ( .A(_170_), .Y(_171_) );
NOR2X1 NOR2X1_118 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_172_) );
INVX1 INVX1_197 ( .A(_172_), .Y(_173_) );
NAND3X1 NAND3X1_111 ( .A(_171_), .B(_173_), .C(_166_), .Y(_174_) );
OAI21X1 OAI21X1_102 ( .A(_168_), .B(_169_), .C(_174_), .Y(w_C_31_) );
NOR2X1 NOR2X1_119 ( .A(_168_), .B(_169_), .Y(_175_) );
INVX1 INVX1_198 ( .A(_175_), .Y(_176_) );
AND2X2 AND2X2_88 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_177_) );
INVX1 INVX1_199 ( .A(_177_), .Y(_178_) );
NAND3X1 NAND3X1_112 ( .A(_176_), .B(_178_), .C(_174_), .Y(_179_) );
OAI21X1 OAI21X1_103 ( .A(i_add2[31]), .B(i_add1[31]), .C(_179_), .Y(_180_) );
INVX1 INVX1_200 ( .A(_180_), .Y(w_C_32_) );
INVX1 INVX1_201 ( .A(i_add2[32]), .Y(_181_) );
INVX1 INVX1_202 ( .A(i_add1[32]), .Y(_182_) );
NOR2X1 NOR2X1_120 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_183_) );
INVX1 INVX1_203 ( .A(_183_), .Y(_184_) );
NOR2X1 NOR2X1_121 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_185_) );
INVX1 INVX1_204 ( .A(_185_), .Y(_186_) );
NAND3X1 NAND3X1_113 ( .A(_184_), .B(_186_), .C(_179_), .Y(_187_) );
OAI21X1 OAI21X1_104 ( .A(_181_), .B(_182_), .C(_187_), .Y(w_C_33_) );
NOR2X1 NOR2X1_122 ( .A(_181_), .B(_182_), .Y(_188_) );
INVX1 INVX1_205 ( .A(_188_), .Y(_189_) );
AND2X2 AND2X2_89 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_190_) );
INVX1 INVX1_206 ( .A(_190_), .Y(_191_) );
NAND3X1 NAND3X1_114 ( .A(_189_), .B(_191_), .C(_187_), .Y(_192_) );
OAI21X1 OAI21X1_105 ( .A(i_add2[33]), .B(i_add1[33]), .C(_192_), .Y(_193_) );
INVX1 INVX1_207 ( .A(_193_), .Y(w_C_34_) );
INVX1 INVX1_208 ( .A(i_add2[34]), .Y(_194_) );
INVX1 INVX1_209 ( .A(i_add1[34]), .Y(_195_) );
NOR2X1 NOR2X1_123 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_196_) );
INVX1 INVX1_210 ( .A(_196_), .Y(_197_) );
NOR2X1 NOR2X1_124 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_198_) );
INVX1 INVX1_211 ( .A(_198_), .Y(_199_) );
NAND3X1 NAND3X1_115 ( .A(_197_), .B(_199_), .C(_192_), .Y(_200_) );
OAI21X1 OAI21X1_106 ( .A(_194_), .B(_195_), .C(_200_), .Y(w_C_35_) );
NOR2X1 NOR2X1_125 ( .A(_194_), .B(_195_), .Y(_201_) );
INVX1 INVX1_212 ( .A(_201_), .Y(_202_) );
AND2X2 AND2X2_90 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_203_) );
INVX1 INVX1_213 ( .A(_203_), .Y(_204_) );
NAND3X1 NAND3X1_116 ( .A(_202_), .B(_204_), .C(_200_), .Y(_205_) );
OAI21X1 OAI21X1_107 ( .A(i_add2[35]), .B(i_add1[35]), .C(_205_), .Y(_206_) );
INVX1 INVX1_214 ( .A(_206_), .Y(w_C_36_) );
INVX1 INVX1_215 ( .A(i_add2[36]), .Y(_207_) );
INVX1 INVX1_216 ( .A(i_add1[36]), .Y(_208_) );
NOR2X1 NOR2X1_126 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_209_) );
INVX1 INVX1_217 ( .A(_209_), .Y(_210_) );
NOR2X1 NOR2X1_127 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_211_) );
INVX1 INVX1_218 ( .A(_211_), .Y(_212_) );
NAND3X1 NAND3X1_117 ( .A(_210_), .B(_212_), .C(_205_), .Y(_213_) );
OAI21X1 OAI21X1_108 ( .A(_207_), .B(_208_), .C(_213_), .Y(w_C_37_) );
NOR2X1 NOR2X1_128 ( .A(_207_), .B(_208_), .Y(_214_) );
INVX1 INVX1_219 ( .A(_214_), .Y(_215_) );
AND2X2 AND2X2_91 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_216_) );
INVX1 INVX1_220 ( .A(_216_), .Y(_217_) );
NAND3X1 NAND3X1_118 ( .A(_215_), .B(_217_), .C(_213_), .Y(_218_) );
OAI21X1 OAI21X1_109 ( .A(i_add2[37]), .B(i_add1[37]), .C(_218_), .Y(_219_) );
INVX1 INVX1_221 ( .A(_219_), .Y(w_C_38_) );
INVX1 INVX1_222 ( .A(i_add2[38]), .Y(_220_) );
INVX1 INVX1_223 ( .A(i_add1[38]), .Y(_221_) );
NOR2X1 NOR2X1_129 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_222_) );
INVX1 INVX1_224 ( .A(_222_), .Y(_223_) );
NOR2X1 NOR2X1_130 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_224_) );
INVX1 INVX1_225 ( .A(_224_), .Y(_225_) );
NAND3X1 NAND3X1_119 ( .A(_223_), .B(_225_), .C(_218_), .Y(_226_) );
OAI21X1 OAI21X1_110 ( .A(_220_), .B(_221_), .C(_226_), .Y(w_C_39_) );
NOR2X1 NOR2X1_131 ( .A(_220_), .B(_221_), .Y(_227_) );
INVX1 INVX1_226 ( .A(_227_), .Y(_228_) );
AND2X2 AND2X2_92 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_229_) );
INVX1 INVX1_227 ( .A(_229_), .Y(_230_) );
NAND3X1 NAND3X1_120 ( .A(_228_), .B(_230_), .C(_226_), .Y(_231_) );
OAI21X1 OAI21X1_111 ( .A(i_add2[39]), .B(i_add1[39]), .C(_231_), .Y(_232_) );
INVX1 INVX1_228 ( .A(_232_), .Y(w_C_40_) );
INVX1 INVX1_229 ( .A(i_add2[40]), .Y(_233_) );
INVX1 INVX1_230 ( .A(i_add1[40]), .Y(_234_) );
NOR2X1 NOR2X1_132 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_235_) );
INVX1 INVX1_231 ( .A(_235_), .Y(_236_) );
NOR2X1 NOR2X1_133 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_237_) );
INVX1 INVX1_232 ( .A(_237_), .Y(_238_) );
NAND3X1 NAND3X1_121 ( .A(_236_), .B(_238_), .C(_231_), .Y(_239_) );
OAI21X1 OAI21X1_112 ( .A(_233_), .B(_234_), .C(_239_), .Y(w_C_41_) );
BUFX2 BUFX2_63 ( .A(w_C_61_), .Y(_355__61_) );
BUFX2 BUFX2_64 ( .A(gnd), .Y(w_C_0_) );
endmodule
