module CSkipA_43bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [42:0] i_add_term1;
input [42:0] i_add_term2;
output [42:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

OAI21X1 OAI21X1_1 ( .A(_403_), .B(_399_), .C(_26__1_), .Y(_400_) );
NAND2X1 NAND2X1_1 ( .A(_400_), .B(_398_), .Y(_0__33_) );
INVX1 INVX1_1 ( .A(_26__2_), .Y(_408_) );
NAND2X1 NAND2X1_2 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_409_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_410_) );
OAI21X1 OAI21X1_2 ( .A(_408_), .B(_410_), .C(_409_), .Y(_26__3_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_404_) );
NAND3X1 NAND3X1_1 ( .A(_408_), .B(_409_), .C(_404_), .Y(_405_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_406_) );
OAI21X1 OAI21X1_3 ( .A(_410_), .B(_406_), .C(_26__2_), .Y(_407_) );
NAND2X1 NAND2X1_3 ( .A(_407_), .B(_405_), .Y(_0__34_) );
INVX1 INVX1_2 ( .A(i_add_term1[32]), .Y(_411_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[32]), .B(_411_), .Y(_412_) );
INVX1 INVX1_3 ( .A(i_add_term2[32]), .Y(_413_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term1[32]), .B(_413_), .Y(_414_) );
INVX1 INVX1_4 ( .A(i_add_term1[33]), .Y(_415_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[33]), .B(_415_), .Y(_416_) );
INVX1 INVX1_5 ( .A(i_add_term2[33]), .Y(_417_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term1[33]), .B(_417_), .Y(_418_) );
OAI22X1 OAI22X1_1 ( .A(_412_), .B(_414_), .C(_416_), .D(_418_), .Y(_419_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_420_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_421_) );
NOR2X1 NOR2X1_7 ( .A(_420_), .B(_421_), .Y(_422_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_423_) );
NAND2X1 NAND2X1_4 ( .A(_422_), .B(_423_), .Y(_424_) );
NOR2X1 NOR2X1_8 ( .A(_419_), .B(_424_), .Y(_27_) );
INVX1 INVX1_6 ( .A(_25_), .Y(_425_) );
NAND2X1 NAND2X1_5 ( .A(gnd), .B(_27_), .Y(_426_) );
OAI21X1 OAI21X1_4 ( .A(_27_), .B(_425_), .C(_426_), .Y(w_cout_9_) );
INVX1 INVX1_7 ( .A(w_cout_9_), .Y(_431_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_432_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_433_) );
OAI21X1 OAI21X1_5 ( .A(_431_), .B(_433_), .C(_432_), .Y(_29__1_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_427_) );
NAND3X1 NAND3X1_2 ( .A(_431_), .B(_432_), .C(_427_), .Y(_428_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_429_) );
OAI21X1 OAI21X1_6 ( .A(_433_), .B(_429_), .C(w_cout_9_), .Y(_430_) );
NAND2X1 NAND2X1_7 ( .A(_430_), .B(_428_), .Y(_0__36_) );
INVX1 INVX1_8 ( .A(_29__3_), .Y(_438_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_439_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_440_) );
OAI21X1 OAI21X1_7 ( .A(_438_), .B(_440_), .C(_439_), .Y(_28_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_434_) );
NAND3X1 NAND3X1_3 ( .A(_438_), .B(_439_), .C(_434_), .Y(_435_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_436_) );
OAI21X1 OAI21X1_8 ( .A(_440_), .B(_436_), .C(_29__3_), .Y(_437_) );
NAND2X1 NAND2X1_9 ( .A(_437_), .B(_435_), .Y(_0__39_) );
INVX1 INVX1_9 ( .A(_29__1_), .Y(_445_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_446_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_447_) );
OAI21X1 OAI21X1_9 ( .A(_445_), .B(_447_), .C(_446_), .Y(_29__2_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_441_) );
NAND3X1 NAND3X1_4 ( .A(_445_), .B(_446_), .C(_441_), .Y(_442_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_443_) );
OAI21X1 OAI21X1_10 ( .A(_447_), .B(_443_), .C(_29__1_), .Y(_444_) );
NAND2X1 NAND2X1_11 ( .A(_444_), .B(_442_), .Y(_0__37_) );
INVX1 INVX1_10 ( .A(_29__2_), .Y(_452_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_453_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_454_) );
OAI21X1 OAI21X1_11 ( .A(_452_), .B(_454_), .C(_453_), .Y(_29__3_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_448_) );
NAND3X1 NAND3X1_5 ( .A(_452_), .B(_453_), .C(_448_), .Y(_449_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_450_) );
OAI21X1 OAI21X1_12 ( .A(_454_), .B(_450_), .C(_29__2_), .Y(_451_) );
NAND2X1 NAND2X1_13 ( .A(_451_), .B(_449_), .Y(_0__38_) );
INVX1 INVX1_11 ( .A(i_add_term1[36]), .Y(_455_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[36]), .B(_455_), .Y(_456_) );
INVX1 INVX1_12 ( .A(i_add_term2[36]), .Y(_457_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term1[36]), .B(_457_), .Y(_458_) );
INVX1 INVX1_13 ( .A(i_add_term1[37]), .Y(_459_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[37]), .B(_459_), .Y(_460_) );
INVX1 INVX1_14 ( .A(i_add_term2[37]), .Y(_461_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term1[37]), .B(_461_), .Y(_462_) );
OAI22X1 OAI22X1_2 ( .A(_456_), .B(_458_), .C(_460_), .D(_462_), .Y(_463_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_464_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_465_) );
NOR2X1 NOR2X1_18 ( .A(_464_), .B(_465_), .Y(_466_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_467_) );
NAND2X1 NAND2X1_14 ( .A(_466_), .B(_467_), .Y(_468_) );
NOR2X1 NOR2X1_19 ( .A(_463_), .B(_468_), .Y(_30_) );
INVX1 INVX1_15 ( .A(_28_), .Y(_469_) );
NAND2X1 NAND2X1_15 ( .A(gnd), .B(_30_), .Y(_470_) );
OAI21X1 OAI21X1_13 ( .A(_30_), .B(_469_), .C(_470_), .Y(cskip3_inst_cin) );
INVX1 INVX1_16 ( .A(cskip3_inst_cin), .Y(_475_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_476_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_477_) );
OAI21X1 OAI21X1_14 ( .A(_475_), .B(_477_), .C(_476_), .Y(cskip3_inst_rca0_fa0_o_carry) );
OR2X2 OR2X2_6 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_471_) );
NAND3X1 NAND3X1_6 ( .A(_475_), .B(_476_), .C(_471_), .Y(_472_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_473_) );
OAI21X1 OAI21X1_15 ( .A(_477_), .B(_473_), .C(cskip3_inst_cin), .Y(_474_) );
NAND2X1 NAND2X1_17 ( .A(_474_), .B(_472_), .Y(cskip3_inst_rca0_fa0_o_sum) );
INVX1 INVX1_17 ( .A(cskip3_inst_rca0_fa0_o_carry), .Y(_482_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_483_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_484_) );
OAI21X1 OAI21X1_16 ( .A(_482_), .B(_484_), .C(_483_), .Y(cskip3_inst_rca0_fa1_o_carry) );
OR2X2 OR2X2_7 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_478_) );
NAND3X1 NAND3X1_7 ( .A(_482_), .B(_483_), .C(_478_), .Y(_479_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_480_) );
OAI21X1 OAI21X1_17 ( .A(_484_), .B(_480_), .C(cskip3_inst_rca0_fa0_o_carry), .Y(_481_) );
NAND2X1 NAND2X1_19 ( .A(_481_), .B(_479_), .Y(cskip3_inst_rca0_fa1_o_sum) );
INVX1 INVX1_18 ( .A(cskip3_inst_rca0_fa1_o_carry), .Y(_489_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_490_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_491_) );
OAI21X1 OAI21X1_18 ( .A(_489_), .B(_491_), .C(_490_), .Y(cskip3_inst_cout0) );
OR2X2 OR2X2_8 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_485_) );
NAND3X1 NAND3X1_8 ( .A(_489_), .B(_490_), .C(_485_), .Y(_486_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_487_) );
OAI21X1 OAI21X1_19 ( .A(_491_), .B(_487_), .C(cskip3_inst_rca0_fa1_o_carry), .Y(_488_) );
NAND2X1 NAND2X1_21 ( .A(_488_), .B(_486_), .Y(cskip3_inst_rca0_fa2_o_sum) );
OR2X2 OR2X2_9 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_495_) );
NAND2X1 NAND2X1_22 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_496_) );
NAND2X1 NAND2X1_23 ( .A(_496_), .B(_495_), .Y(_492_) );
XNOR2X1 XNOR2X1_1 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_493_) );
XNOR2X1 XNOR2X1_2 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_494_) );
NOR3X1 NOR3X1_1 ( .A(_492_), .B(_493_), .C(_494_), .Y(cskip3_inst_skip0_P) );
INVX1 INVX1_19 ( .A(cskip3_inst_cout0), .Y(_497_) );
NAND2X1 NAND2X1_24 ( .A(gnd), .B(cskip3_inst_skip0_P), .Y(_498_) );
OAI21X1 OAI21X1_20 ( .A(cskip3_inst_skip0_P), .B(_497_), .C(_498_), .Y(w_cout_11_) );
BUFX2 BUFX2_1 ( .A(w_cout_11_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(cskip3_inst_rca0_fa0_o_sum), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(cskip3_inst_rca0_fa1_o_sum), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(cskip3_inst_rca0_fa2_o_sum), .Y(sum[42]) );
INVX1 INVX1_20 ( .A(gnd), .Y(_35_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_36_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_37_) );
OAI21X1 OAI21X1_21 ( .A(_35_), .B(_37_), .C(_36_), .Y(_2__1_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_31_) );
NAND3X1 NAND3X1_9 ( .A(_35_), .B(_36_), .C(_31_), .Y(_32_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_33_) );
OAI21X1 OAI21X1_22 ( .A(_37_), .B(_33_), .C(gnd), .Y(_34_) );
NAND2X1 NAND2X1_26 ( .A(_34_), .B(_32_), .Y(_0__0_) );
INVX1 INVX1_21 ( .A(_2__3_), .Y(_42_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_43_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_44_) );
OAI21X1 OAI21X1_23 ( .A(_42_), .B(_44_), .C(_43_), .Y(_1_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_38_) );
NAND3X1 NAND3X1_10 ( .A(_42_), .B(_43_), .C(_38_), .Y(_39_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_40_) );
OAI21X1 OAI21X1_24 ( .A(_44_), .B(_40_), .C(_2__3_), .Y(_41_) );
NAND2X1 NAND2X1_28 ( .A(_41_), .B(_39_), .Y(_0__3_) );
INVX1 INVX1_22 ( .A(_2__1_), .Y(_49_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_50_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_51_) );
OAI21X1 OAI21X1_25 ( .A(_49_), .B(_51_), .C(_50_), .Y(_2__2_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_45_) );
NAND3X1 NAND3X1_11 ( .A(_49_), .B(_50_), .C(_45_), .Y(_46_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_47_) );
OAI21X1 OAI21X1_26 ( .A(_51_), .B(_47_), .C(_2__1_), .Y(_48_) );
NAND2X1 NAND2X1_30 ( .A(_48_), .B(_46_), .Y(_0__1_) );
INVX1 INVX1_23 ( .A(_2__2_), .Y(_56_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_57_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_58_) );
OAI21X1 OAI21X1_27 ( .A(_56_), .B(_58_), .C(_57_), .Y(_2__3_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_52_) );
NAND3X1 NAND3X1_12 ( .A(_56_), .B(_57_), .C(_52_), .Y(_53_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_54_) );
OAI21X1 OAI21X1_28 ( .A(_58_), .B(_54_), .C(_2__2_), .Y(_55_) );
NAND2X1 NAND2X1_32 ( .A(_55_), .B(_53_), .Y(_0__2_) );
INVX1 INVX1_24 ( .A(i_add_term1[0]), .Y(_59_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[0]), .B(_59_), .Y(_60_) );
INVX1 INVX1_25 ( .A(i_add_term2[0]), .Y(_61_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term1[0]), .B(_61_), .Y(_62_) );
INVX1 INVX1_26 ( .A(i_add_term1[1]), .Y(_63_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[1]), .B(_63_), .Y(_64_) );
INVX1 INVX1_27 ( .A(i_add_term2[1]), .Y(_65_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term1[1]), .B(_65_), .Y(_66_) );
OAI22X1 OAI22X1_3 ( .A(_60_), .B(_62_), .C(_64_), .D(_66_), .Y(_67_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_68_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_69_) );
NOR2X1 NOR2X1_32 ( .A(_68_), .B(_69_), .Y(_70_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_71_) );
NAND2X1 NAND2X1_33 ( .A(_70_), .B(_71_), .Y(_72_) );
NOR2X1 NOR2X1_33 ( .A(_67_), .B(_72_), .Y(_3_) );
INVX1 INVX1_28 ( .A(_1_), .Y(_73_) );
NAND2X1 NAND2X1_34 ( .A(gnd), .B(_3_), .Y(_74_) );
OAI21X1 OAI21X1_29 ( .A(_3_), .B(_73_), .C(_74_), .Y(w_cout_1_) );
INVX1 INVX1_29 ( .A(w_cout_1_), .Y(_79_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_80_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_81_) );
OAI21X1 OAI21X1_30 ( .A(_79_), .B(_81_), .C(_80_), .Y(_5__1_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_75_) );
NAND3X1 NAND3X1_13 ( .A(_79_), .B(_80_), .C(_75_), .Y(_76_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_77_) );
OAI21X1 OAI21X1_31 ( .A(_81_), .B(_77_), .C(w_cout_1_), .Y(_78_) );
NAND2X1 NAND2X1_36 ( .A(_78_), .B(_76_), .Y(_0__4_) );
INVX1 INVX1_30 ( .A(_5__3_), .Y(_86_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_87_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_88_) );
OAI21X1 OAI21X1_32 ( .A(_86_), .B(_88_), .C(_87_), .Y(_4_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_82_) );
NAND3X1 NAND3X1_14 ( .A(_86_), .B(_87_), .C(_82_), .Y(_83_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_84_) );
OAI21X1 OAI21X1_33 ( .A(_88_), .B(_84_), .C(_5__3_), .Y(_85_) );
NAND2X1 NAND2X1_38 ( .A(_85_), .B(_83_), .Y(_0__7_) );
INVX1 INVX1_31 ( .A(_5__1_), .Y(_93_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_94_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_95_) );
OAI21X1 OAI21X1_34 ( .A(_93_), .B(_95_), .C(_94_), .Y(_5__2_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_89_) );
NAND3X1 NAND3X1_15 ( .A(_93_), .B(_94_), .C(_89_), .Y(_90_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_91_) );
OAI21X1 OAI21X1_35 ( .A(_95_), .B(_91_), .C(_5__1_), .Y(_92_) );
NAND2X1 NAND2X1_40 ( .A(_92_), .B(_90_), .Y(_0__5_) );
INVX1 INVX1_32 ( .A(_5__2_), .Y(_100_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_101_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_102_) );
OAI21X1 OAI21X1_36 ( .A(_100_), .B(_102_), .C(_101_), .Y(_5__3_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_96_) );
NAND3X1 NAND3X1_16 ( .A(_100_), .B(_101_), .C(_96_), .Y(_97_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_98_) );
OAI21X1 OAI21X1_37 ( .A(_102_), .B(_98_), .C(_5__2_), .Y(_99_) );
NAND2X1 NAND2X1_42 ( .A(_99_), .B(_97_), .Y(_0__6_) );
INVX1 INVX1_33 ( .A(i_add_term1[4]), .Y(_103_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[4]), .B(_103_), .Y(_104_) );
INVX1 INVX1_34 ( .A(i_add_term2[4]), .Y(_105_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term1[4]), .B(_105_), .Y(_106_) );
INVX1 INVX1_35 ( .A(i_add_term1[5]), .Y(_107_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[5]), .B(_107_), .Y(_108_) );
INVX1 INVX1_36 ( .A(i_add_term2[5]), .Y(_109_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term1[5]), .B(_109_), .Y(_110_) );
OAI22X1 OAI22X1_4 ( .A(_104_), .B(_106_), .C(_108_), .D(_110_), .Y(_111_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_112_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_113_) );
NOR2X1 NOR2X1_43 ( .A(_112_), .B(_113_), .Y(_114_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_115_) );
NAND2X1 NAND2X1_43 ( .A(_114_), .B(_115_), .Y(_116_) );
NOR2X1 NOR2X1_44 ( .A(_111_), .B(_116_), .Y(_6_) );
INVX1 INVX1_37 ( .A(_4_), .Y(_117_) );
NAND2X1 NAND2X1_44 ( .A(gnd), .B(_6_), .Y(_118_) );
OAI21X1 OAI21X1_38 ( .A(_6_), .B(_117_), .C(_118_), .Y(w_cout_2_) );
INVX1 INVX1_38 ( .A(w_cout_2_), .Y(_123_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_124_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_125_) );
OAI21X1 OAI21X1_39 ( .A(_123_), .B(_125_), .C(_124_), .Y(_8__1_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_119_) );
NAND3X1 NAND3X1_17 ( .A(_123_), .B(_124_), .C(_119_), .Y(_120_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_121_) );
OAI21X1 OAI21X1_40 ( .A(_125_), .B(_121_), .C(w_cout_2_), .Y(_122_) );
NAND2X1 NAND2X1_46 ( .A(_122_), .B(_120_), .Y(_0__8_) );
INVX1 INVX1_39 ( .A(_8__3_), .Y(_130_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_131_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_132_) );
OAI21X1 OAI21X1_41 ( .A(_130_), .B(_132_), .C(_131_), .Y(_7_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_126_) );
NAND3X1 NAND3X1_18 ( .A(_130_), .B(_131_), .C(_126_), .Y(_127_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_128_) );
OAI21X1 OAI21X1_42 ( .A(_132_), .B(_128_), .C(_8__3_), .Y(_129_) );
NAND2X1 NAND2X1_48 ( .A(_129_), .B(_127_), .Y(_0__11_) );
INVX1 INVX1_40 ( .A(_8__1_), .Y(_137_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_138_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_139_) );
OAI21X1 OAI21X1_43 ( .A(_137_), .B(_139_), .C(_138_), .Y(_8__2_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_133_) );
NAND3X1 NAND3X1_19 ( .A(_137_), .B(_138_), .C(_133_), .Y(_134_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_135_) );
OAI21X1 OAI21X1_44 ( .A(_139_), .B(_135_), .C(_8__1_), .Y(_136_) );
NAND2X1 NAND2X1_50 ( .A(_136_), .B(_134_), .Y(_0__9_) );
INVX1 INVX1_41 ( .A(_8__2_), .Y(_144_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_145_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_146_) );
OAI21X1 OAI21X1_45 ( .A(_144_), .B(_146_), .C(_145_), .Y(_8__3_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_140_) );
NAND3X1 NAND3X1_20 ( .A(_144_), .B(_145_), .C(_140_), .Y(_141_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_142_) );
OAI21X1 OAI21X1_46 ( .A(_146_), .B(_142_), .C(_8__2_), .Y(_143_) );
NAND2X1 NAND2X1_52 ( .A(_143_), .B(_141_), .Y(_0__10_) );
INVX1 INVX1_42 ( .A(i_add_term1[8]), .Y(_147_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[8]), .B(_147_), .Y(_148_) );
INVX1 INVX1_43 ( .A(i_add_term2[8]), .Y(_149_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term1[8]), .B(_149_), .Y(_150_) );
INVX1 INVX1_44 ( .A(i_add_term1[9]), .Y(_151_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[9]), .B(_151_), .Y(_152_) );
INVX1 INVX1_45 ( .A(i_add_term2[9]), .Y(_153_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term1[9]), .B(_153_), .Y(_154_) );
OAI22X1 OAI22X1_5 ( .A(_148_), .B(_150_), .C(_152_), .D(_154_), .Y(_155_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_156_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_157_) );
NOR2X1 NOR2X1_54 ( .A(_156_), .B(_157_), .Y(_158_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_159_) );
NAND2X1 NAND2X1_53 ( .A(_158_), .B(_159_), .Y(_160_) );
NOR2X1 NOR2X1_55 ( .A(_155_), .B(_160_), .Y(_9_) );
INVX1 INVX1_46 ( .A(_7_), .Y(_161_) );
NAND2X1 NAND2X1_54 ( .A(gnd), .B(_9_), .Y(_162_) );
OAI21X1 OAI21X1_47 ( .A(_9_), .B(_161_), .C(_162_), .Y(w_cout_3_) );
INVX1 INVX1_47 ( .A(w_cout_3_), .Y(_167_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_168_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_169_) );
OAI21X1 OAI21X1_48 ( .A(_167_), .B(_169_), .C(_168_), .Y(_11__1_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_163_) );
NAND3X1 NAND3X1_21 ( .A(_167_), .B(_168_), .C(_163_), .Y(_164_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_165_) );
OAI21X1 OAI21X1_49 ( .A(_169_), .B(_165_), .C(w_cout_3_), .Y(_166_) );
NAND2X1 NAND2X1_56 ( .A(_166_), .B(_164_), .Y(_0__12_) );
INVX1 INVX1_48 ( .A(_11__3_), .Y(_174_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_175_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_176_) );
OAI21X1 OAI21X1_50 ( .A(_174_), .B(_176_), .C(_175_), .Y(_10_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_170_) );
NAND3X1 NAND3X1_22 ( .A(_174_), .B(_175_), .C(_170_), .Y(_171_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_172_) );
OAI21X1 OAI21X1_51 ( .A(_176_), .B(_172_), .C(_11__3_), .Y(_173_) );
NAND2X1 NAND2X1_58 ( .A(_173_), .B(_171_), .Y(_0__15_) );
INVX1 INVX1_49 ( .A(_11__1_), .Y(_181_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_182_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_183_) );
OAI21X1 OAI21X1_52 ( .A(_181_), .B(_183_), .C(_182_), .Y(_11__2_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_177_) );
NAND3X1 NAND3X1_23 ( .A(_181_), .B(_182_), .C(_177_), .Y(_178_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_179_) );
OAI21X1 OAI21X1_53 ( .A(_183_), .B(_179_), .C(_11__1_), .Y(_180_) );
NAND2X1 NAND2X1_60 ( .A(_180_), .B(_178_), .Y(_0__13_) );
INVX1 INVX1_50 ( .A(_11__2_), .Y(_188_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_189_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_190_) );
OAI21X1 OAI21X1_54 ( .A(_188_), .B(_190_), .C(_189_), .Y(_11__3_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_184_) );
NAND3X1 NAND3X1_24 ( .A(_188_), .B(_189_), .C(_184_), .Y(_185_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_186_) );
OAI21X1 OAI21X1_55 ( .A(_190_), .B(_186_), .C(_11__2_), .Y(_187_) );
NAND2X1 NAND2X1_62 ( .A(_187_), .B(_185_), .Y(_0__14_) );
INVX1 INVX1_51 ( .A(i_add_term1[12]), .Y(_191_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[12]), .B(_191_), .Y(_192_) );
INVX1 INVX1_52 ( .A(i_add_term2[12]), .Y(_193_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term1[12]), .B(_193_), .Y(_194_) );
INVX1 INVX1_53 ( .A(i_add_term1[13]), .Y(_195_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[13]), .B(_195_), .Y(_196_) );
INVX1 INVX1_54 ( .A(i_add_term2[13]), .Y(_197_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term1[13]), .B(_197_), .Y(_198_) );
OAI22X1 OAI22X1_6 ( .A(_192_), .B(_194_), .C(_196_), .D(_198_), .Y(_199_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_200_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_201_) );
NOR2X1 NOR2X1_65 ( .A(_200_), .B(_201_), .Y(_202_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_203_) );
NAND2X1 NAND2X1_63 ( .A(_202_), .B(_203_), .Y(_204_) );
NOR2X1 NOR2X1_66 ( .A(_199_), .B(_204_), .Y(_12_) );
INVX1 INVX1_55 ( .A(_10_), .Y(_205_) );
NAND2X1 NAND2X1_64 ( .A(gnd), .B(_12_), .Y(_206_) );
OAI21X1 OAI21X1_56 ( .A(_12_), .B(_205_), .C(_206_), .Y(w_cout_4_) );
INVX1 INVX1_56 ( .A(w_cout_4_), .Y(_211_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_212_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_213_) );
OAI21X1 OAI21X1_57 ( .A(_211_), .B(_213_), .C(_212_), .Y(_14__1_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_207_) );
NAND3X1 NAND3X1_25 ( .A(_211_), .B(_212_), .C(_207_), .Y(_208_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_209_) );
OAI21X1 OAI21X1_58 ( .A(_213_), .B(_209_), .C(w_cout_4_), .Y(_210_) );
NAND2X1 NAND2X1_66 ( .A(_210_), .B(_208_), .Y(_0__16_) );
INVX1 INVX1_57 ( .A(_14__3_), .Y(_218_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_219_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_220_) );
OAI21X1 OAI21X1_59 ( .A(_218_), .B(_220_), .C(_219_), .Y(_13_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_214_) );
NAND3X1 NAND3X1_26 ( .A(_218_), .B(_219_), .C(_214_), .Y(_215_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_216_) );
OAI21X1 OAI21X1_60 ( .A(_220_), .B(_216_), .C(_14__3_), .Y(_217_) );
NAND2X1 NAND2X1_68 ( .A(_217_), .B(_215_), .Y(_0__19_) );
INVX1 INVX1_58 ( .A(_14__1_), .Y(_225_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_226_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_227_) );
OAI21X1 OAI21X1_61 ( .A(_225_), .B(_227_), .C(_226_), .Y(_14__2_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_221_) );
NAND3X1 NAND3X1_27 ( .A(_225_), .B(_226_), .C(_221_), .Y(_222_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_223_) );
OAI21X1 OAI21X1_62 ( .A(_227_), .B(_223_), .C(_14__1_), .Y(_224_) );
NAND2X1 NAND2X1_70 ( .A(_224_), .B(_222_), .Y(_0__17_) );
INVX1 INVX1_59 ( .A(_14__2_), .Y(_232_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_233_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_234_) );
OAI21X1 OAI21X1_63 ( .A(_232_), .B(_234_), .C(_233_), .Y(_14__3_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_228_) );
NAND3X1 NAND3X1_28 ( .A(_232_), .B(_233_), .C(_228_), .Y(_229_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_230_) );
OAI21X1 OAI21X1_64 ( .A(_234_), .B(_230_), .C(_14__2_), .Y(_231_) );
NAND2X1 NAND2X1_72 ( .A(_231_), .B(_229_), .Y(_0__18_) );
INVX1 INVX1_60 ( .A(i_add_term1[16]), .Y(_235_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[16]), .B(_235_), .Y(_236_) );
INVX1 INVX1_61 ( .A(i_add_term2[16]), .Y(_237_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term1[16]), .B(_237_), .Y(_238_) );
INVX1 INVX1_62 ( .A(i_add_term1[17]), .Y(_239_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[17]), .B(_239_), .Y(_240_) );
INVX1 INVX1_63 ( .A(i_add_term2[17]), .Y(_241_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term1[17]), .B(_241_), .Y(_242_) );
OAI22X1 OAI22X1_7 ( .A(_236_), .B(_238_), .C(_240_), .D(_242_), .Y(_243_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_244_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_245_) );
NOR2X1 NOR2X1_76 ( .A(_244_), .B(_245_), .Y(_246_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_247_) );
NAND2X1 NAND2X1_73 ( .A(_246_), .B(_247_), .Y(_248_) );
NOR2X1 NOR2X1_77 ( .A(_243_), .B(_248_), .Y(_15_) );
INVX1 INVX1_64 ( .A(_13_), .Y(_249_) );
NAND2X1 NAND2X1_74 ( .A(gnd), .B(_15_), .Y(_250_) );
OAI21X1 OAI21X1_65 ( .A(_15_), .B(_249_), .C(_250_), .Y(w_cout_5_) );
INVX1 INVX1_65 ( .A(w_cout_5_), .Y(_255_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_256_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_257_) );
OAI21X1 OAI21X1_66 ( .A(_255_), .B(_257_), .C(_256_), .Y(_17__1_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_251_) );
NAND3X1 NAND3X1_29 ( .A(_255_), .B(_256_), .C(_251_), .Y(_252_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_253_) );
OAI21X1 OAI21X1_67 ( .A(_257_), .B(_253_), .C(w_cout_5_), .Y(_254_) );
NAND2X1 NAND2X1_76 ( .A(_254_), .B(_252_), .Y(_0__20_) );
INVX1 INVX1_66 ( .A(_17__3_), .Y(_262_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_263_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_264_) );
OAI21X1 OAI21X1_68 ( .A(_262_), .B(_264_), .C(_263_), .Y(_16_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_258_) );
NAND3X1 NAND3X1_30 ( .A(_262_), .B(_263_), .C(_258_), .Y(_259_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_260_) );
OAI21X1 OAI21X1_69 ( .A(_264_), .B(_260_), .C(_17__3_), .Y(_261_) );
NAND2X1 NAND2X1_78 ( .A(_261_), .B(_259_), .Y(_0__23_) );
INVX1 INVX1_67 ( .A(_17__1_), .Y(_269_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_270_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_271_) );
OAI21X1 OAI21X1_70 ( .A(_269_), .B(_271_), .C(_270_), .Y(_17__2_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_265_) );
NAND3X1 NAND3X1_31 ( .A(_269_), .B(_270_), .C(_265_), .Y(_266_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_267_) );
OAI21X1 OAI21X1_71 ( .A(_271_), .B(_267_), .C(_17__1_), .Y(_268_) );
NAND2X1 NAND2X1_80 ( .A(_268_), .B(_266_), .Y(_0__21_) );
INVX1 INVX1_68 ( .A(_17__2_), .Y(_276_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_277_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_278_) );
OAI21X1 OAI21X1_72 ( .A(_276_), .B(_278_), .C(_277_), .Y(_17__3_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_272_) );
NAND3X1 NAND3X1_32 ( .A(_276_), .B(_277_), .C(_272_), .Y(_273_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_274_) );
OAI21X1 OAI21X1_73 ( .A(_278_), .B(_274_), .C(_17__2_), .Y(_275_) );
NAND2X1 NAND2X1_82 ( .A(_275_), .B(_273_), .Y(_0__22_) );
INVX1 INVX1_69 ( .A(i_add_term1[20]), .Y(_279_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[20]), .B(_279_), .Y(_280_) );
INVX1 INVX1_70 ( .A(i_add_term2[20]), .Y(_281_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term1[20]), .B(_281_), .Y(_282_) );
INVX1 INVX1_71 ( .A(i_add_term1[21]), .Y(_283_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[21]), .B(_283_), .Y(_284_) );
INVX1 INVX1_72 ( .A(i_add_term2[21]), .Y(_285_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term1[21]), .B(_285_), .Y(_286_) );
OAI22X1 OAI22X1_8 ( .A(_280_), .B(_282_), .C(_284_), .D(_286_), .Y(_287_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_288_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_289_) );
NOR2X1 NOR2X1_87 ( .A(_288_), .B(_289_), .Y(_290_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_291_) );
NAND2X1 NAND2X1_83 ( .A(_290_), .B(_291_), .Y(_292_) );
NOR2X1 NOR2X1_88 ( .A(_287_), .B(_292_), .Y(_18_) );
INVX1 INVX1_73 ( .A(_16_), .Y(_293_) );
NAND2X1 NAND2X1_84 ( .A(gnd), .B(_18_), .Y(_294_) );
OAI21X1 OAI21X1_74 ( .A(_18_), .B(_293_), .C(_294_), .Y(w_cout_6_) );
INVX1 INVX1_74 ( .A(w_cout_6_), .Y(_299_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_300_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_301_) );
OAI21X1 OAI21X1_75 ( .A(_299_), .B(_301_), .C(_300_), .Y(_20__1_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_295_) );
NAND3X1 NAND3X1_33 ( .A(_299_), .B(_300_), .C(_295_), .Y(_296_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_297_) );
OAI21X1 OAI21X1_76 ( .A(_301_), .B(_297_), .C(w_cout_6_), .Y(_298_) );
NAND2X1 NAND2X1_86 ( .A(_298_), .B(_296_), .Y(_0__24_) );
INVX1 INVX1_75 ( .A(_20__3_), .Y(_306_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_307_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_308_) );
OAI21X1 OAI21X1_77 ( .A(_306_), .B(_308_), .C(_307_), .Y(_19_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_302_) );
NAND3X1 NAND3X1_34 ( .A(_306_), .B(_307_), .C(_302_), .Y(_303_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_304_) );
OAI21X1 OAI21X1_78 ( .A(_308_), .B(_304_), .C(_20__3_), .Y(_305_) );
NAND2X1 NAND2X1_88 ( .A(_305_), .B(_303_), .Y(_0__27_) );
INVX1 INVX1_76 ( .A(_20__1_), .Y(_313_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_314_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_315_) );
OAI21X1 OAI21X1_79 ( .A(_313_), .B(_315_), .C(_314_), .Y(_20__2_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_309_) );
NAND3X1 NAND3X1_35 ( .A(_313_), .B(_314_), .C(_309_), .Y(_310_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_311_) );
OAI21X1 OAI21X1_80 ( .A(_315_), .B(_311_), .C(_20__1_), .Y(_312_) );
NAND2X1 NAND2X1_90 ( .A(_312_), .B(_310_), .Y(_0__25_) );
INVX1 INVX1_77 ( .A(_20__2_), .Y(_320_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_321_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_322_) );
OAI21X1 OAI21X1_81 ( .A(_320_), .B(_322_), .C(_321_), .Y(_20__3_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_316_) );
NAND3X1 NAND3X1_36 ( .A(_320_), .B(_321_), .C(_316_), .Y(_317_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_318_) );
OAI21X1 OAI21X1_82 ( .A(_322_), .B(_318_), .C(_20__2_), .Y(_319_) );
NAND2X1 NAND2X1_92 ( .A(_319_), .B(_317_), .Y(_0__26_) );
INVX1 INVX1_78 ( .A(i_add_term1[24]), .Y(_323_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[24]), .B(_323_), .Y(_324_) );
INVX1 INVX1_79 ( .A(i_add_term2[24]), .Y(_325_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term1[24]), .B(_325_), .Y(_326_) );
INVX1 INVX1_80 ( .A(i_add_term1[25]), .Y(_327_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[25]), .B(_327_), .Y(_328_) );
INVX1 INVX1_81 ( .A(i_add_term2[25]), .Y(_329_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term1[25]), .B(_329_), .Y(_330_) );
OAI22X1 OAI22X1_9 ( .A(_324_), .B(_326_), .C(_328_), .D(_330_), .Y(_331_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_332_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_333_) );
NOR2X1 NOR2X1_98 ( .A(_332_), .B(_333_), .Y(_334_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_335_) );
NAND2X1 NAND2X1_93 ( .A(_334_), .B(_335_), .Y(_336_) );
NOR2X1 NOR2X1_99 ( .A(_331_), .B(_336_), .Y(_21_) );
INVX1 INVX1_82 ( .A(_19_), .Y(_337_) );
NAND2X1 NAND2X1_94 ( .A(gnd), .B(_21_), .Y(_338_) );
OAI21X1 OAI21X1_83 ( .A(_21_), .B(_337_), .C(_338_), .Y(w_cout_7_) );
INVX1 INVX1_83 ( .A(w_cout_7_), .Y(_343_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_344_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_345_) );
OAI21X1 OAI21X1_84 ( .A(_343_), .B(_345_), .C(_344_), .Y(_23__1_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_339_) );
NAND3X1 NAND3X1_37 ( .A(_343_), .B(_344_), .C(_339_), .Y(_340_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_341_) );
OAI21X1 OAI21X1_85 ( .A(_345_), .B(_341_), .C(w_cout_7_), .Y(_342_) );
NAND2X1 NAND2X1_96 ( .A(_342_), .B(_340_), .Y(_0__28_) );
INVX1 INVX1_84 ( .A(_23__3_), .Y(_350_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_351_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_352_) );
OAI21X1 OAI21X1_86 ( .A(_350_), .B(_352_), .C(_351_), .Y(_22_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_346_) );
NAND3X1 NAND3X1_38 ( .A(_350_), .B(_351_), .C(_346_), .Y(_347_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_348_) );
OAI21X1 OAI21X1_87 ( .A(_352_), .B(_348_), .C(_23__3_), .Y(_349_) );
NAND2X1 NAND2X1_98 ( .A(_349_), .B(_347_), .Y(_0__31_) );
INVX1 INVX1_85 ( .A(_23__1_), .Y(_357_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_358_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_359_) );
OAI21X1 OAI21X1_88 ( .A(_357_), .B(_359_), .C(_358_), .Y(_23__2_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_353_) );
NAND3X1 NAND3X1_39 ( .A(_357_), .B(_358_), .C(_353_), .Y(_354_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_355_) );
OAI21X1 OAI21X1_89 ( .A(_359_), .B(_355_), .C(_23__1_), .Y(_356_) );
NAND2X1 NAND2X1_100 ( .A(_356_), .B(_354_), .Y(_0__29_) );
INVX1 INVX1_86 ( .A(_23__2_), .Y(_364_) );
NAND2X1 NAND2X1_101 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_365_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_366_) );
OAI21X1 OAI21X1_90 ( .A(_364_), .B(_366_), .C(_365_), .Y(_23__3_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_360_) );
NAND3X1 NAND3X1_40 ( .A(_364_), .B(_365_), .C(_360_), .Y(_361_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_362_) );
OAI21X1 OAI21X1_91 ( .A(_366_), .B(_362_), .C(_23__2_), .Y(_363_) );
NAND2X1 NAND2X1_102 ( .A(_363_), .B(_361_), .Y(_0__30_) );
INVX1 INVX1_87 ( .A(i_add_term1[28]), .Y(_367_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term2[28]), .B(_367_), .Y(_368_) );
INVX1 INVX1_88 ( .A(i_add_term2[28]), .Y(_369_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term1[28]), .B(_369_), .Y(_370_) );
INVX1 INVX1_89 ( .A(i_add_term1[29]), .Y(_371_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term2[29]), .B(_371_), .Y(_372_) );
INVX1 INVX1_90 ( .A(i_add_term2[29]), .Y(_373_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term1[29]), .B(_373_), .Y(_374_) );
OAI22X1 OAI22X1_10 ( .A(_368_), .B(_370_), .C(_372_), .D(_374_), .Y(_375_) );
NOR2X1 NOR2X1_108 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_376_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_377_) );
NOR2X1 NOR2X1_109 ( .A(_376_), .B(_377_), .Y(_378_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_379_) );
NAND2X1 NAND2X1_103 ( .A(_378_), .B(_379_), .Y(_380_) );
NOR2X1 NOR2X1_110 ( .A(_375_), .B(_380_), .Y(_24_) );
INVX1 INVX1_91 ( .A(_22_), .Y(_381_) );
NAND2X1 NAND2X1_104 ( .A(gnd), .B(_24_), .Y(_382_) );
OAI21X1 OAI21X1_92 ( .A(_24_), .B(_381_), .C(_382_), .Y(w_cout_8_) );
INVX1 INVX1_92 ( .A(w_cout_8_), .Y(_387_) );
NAND2X1 NAND2X1_105 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_388_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_389_) );
OAI21X1 OAI21X1_93 ( .A(_387_), .B(_389_), .C(_388_), .Y(_26__1_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_383_) );
NAND3X1 NAND3X1_41 ( .A(_387_), .B(_388_), .C(_383_), .Y(_384_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_385_) );
OAI21X1 OAI21X1_94 ( .A(_389_), .B(_385_), .C(w_cout_8_), .Y(_386_) );
NAND2X1 NAND2X1_106 ( .A(_386_), .B(_384_), .Y(_0__32_) );
INVX1 INVX1_93 ( .A(_26__3_), .Y(_394_) );
NAND2X1 NAND2X1_107 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_395_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_396_) );
OAI21X1 OAI21X1_95 ( .A(_394_), .B(_396_), .C(_395_), .Y(_25_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_390_) );
NAND3X1 NAND3X1_42 ( .A(_394_), .B(_395_), .C(_390_), .Y(_391_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_392_) );
OAI21X1 OAI21X1_96 ( .A(_396_), .B(_392_), .C(_26__3_), .Y(_393_) );
NAND2X1 NAND2X1_108 ( .A(_393_), .B(_391_), .Y(_0__35_) );
INVX1 INVX1_94 ( .A(_26__1_), .Y(_401_) );
NAND2X1 NAND2X1_109 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_402_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_403_) );
OAI21X1 OAI21X1_97 ( .A(_401_), .B(_403_), .C(_402_), .Y(_26__2_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_397_) );
NAND3X1 NAND3X1_43 ( .A(_401_), .B(_402_), .C(_397_), .Y(_398_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_399_) );
BUFX2 BUFX2_45 ( .A(cskip3_inst_rca0_fa0_o_sum), .Y(_0__40_) );
BUFX2 BUFX2_46 ( .A(cskip3_inst_rca0_fa1_o_sum), .Y(_0__41_) );
BUFX2 BUFX2_47 ( .A(cskip3_inst_rca0_fa2_o_sum), .Y(_0__42_) );
BUFX2 BUFX2_48 ( .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_49 ( .A(cskip3_inst_cin), .Y(w_cout_10_) );
endmodule
