module CSkipA_50bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term1[45], i_add_term1[46], i_add_term1[47], i_add_term1[48], i_add_term1[49], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], i_add_term2[45], i_add_term2[46], i_add_term2[47], i_add_term2[48], i_add_term2[49], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], sum[45], sum[46], sum[47], sum[48], sum[49], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term1[45];
input i_add_term1[46];
input i_add_term1[47];
input i_add_term1[48];
input i_add_term1[49];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
input i_add_term2[45];
input i_add_term2[46];
input i_add_term2[47];
input i_add_term2[48];
input i_add_term2[49];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output sum[45];
output sum[46];
output sum[47];
output sum[48];
output sum[49];
output cout;

INVX1 INVX1_1 ( .A(i_add_term1[24]), .Y(_329_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[24]), .B(_329_), .Y(_330_) );
INVX1 INVX1_2 ( .A(i_add_term2[24]), .Y(_331_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term1[24]), .B(_331_), .Y(_332_) );
INVX1 INVX1_3 ( .A(i_add_term1[25]), .Y(_333_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[25]), .B(_333_), .Y(_334_) );
INVX1 INVX1_4 ( .A(i_add_term2[25]), .Y(_335_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term1[25]), .B(_335_), .Y(_336_) );
OAI22X1 OAI22X1_1 ( .A(_330_), .B(_332_), .C(_334_), .D(_336_), .Y(_337_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_338_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_339_) );
NOR2X1 NOR2X1_6 ( .A(_338_), .B(_339_), .Y(_340_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_341_) );
NAND2X1 NAND2X1_1 ( .A(_340_), .B(_341_), .Y(_342_) );
NOR2X1 NOR2X1_7 ( .A(_337_), .B(_342_), .Y(_21_) );
INVX1 INVX1_5 ( .A(_19_), .Y(_343_) );
NAND2X1 NAND2X1_2 ( .A(1'b0), .B(_21_), .Y(_344_) );
OAI21X1 OAI21X1_1 ( .A(_21_), .B(_343_), .C(_344_), .Y(w_cout_7_) );
INVX1 INVX1_6 ( .A(w_cout_7_), .Y(_349_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_350_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_351_) );
OAI21X1 OAI21X1_2 ( .A(_349_), .B(_351_), .C(_350_), .Y(_23__1_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_345_) );
NAND3X1 NAND3X1_1 ( .A(_349_), .B(_350_), .C(_345_), .Y(_346_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_347_) );
OAI21X1 OAI21X1_3 ( .A(_351_), .B(_347_), .C(w_cout_7_), .Y(_348_) );
NAND2X1 NAND2X1_4 ( .A(_348_), .B(_346_), .Y(_0__28_) );
INVX1 INVX1_7 ( .A(_23__3_), .Y(_356_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_357_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_358_) );
OAI21X1 OAI21X1_4 ( .A(_356_), .B(_358_), .C(_357_), .Y(_22_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_352_) );
NAND3X1 NAND3X1_2 ( .A(_356_), .B(_357_), .C(_352_), .Y(_353_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_354_) );
OAI21X1 OAI21X1_5 ( .A(_358_), .B(_354_), .C(_23__3_), .Y(_355_) );
NAND2X1 NAND2X1_6 ( .A(_355_), .B(_353_), .Y(_0__31_) );
INVX1 INVX1_8 ( .A(_23__1_), .Y(_363_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_364_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_365_) );
OAI21X1 OAI21X1_6 ( .A(_363_), .B(_365_), .C(_364_), .Y(_23__2_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_359_) );
NAND3X1 NAND3X1_3 ( .A(_363_), .B(_364_), .C(_359_), .Y(_360_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_361_) );
OAI21X1 OAI21X1_7 ( .A(_365_), .B(_361_), .C(_23__1_), .Y(_362_) );
NAND2X1 NAND2X1_8 ( .A(_362_), .B(_360_), .Y(_0__29_) );
INVX1 INVX1_9 ( .A(_23__2_), .Y(_370_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_371_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_372_) );
OAI21X1 OAI21X1_8 ( .A(_370_), .B(_372_), .C(_371_), .Y(_23__3_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_366_) );
NAND3X1 NAND3X1_4 ( .A(_370_), .B(_371_), .C(_366_), .Y(_367_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_368_) );
OAI21X1 OAI21X1_9 ( .A(_372_), .B(_368_), .C(_23__2_), .Y(_369_) );
NAND2X1 NAND2X1_10 ( .A(_369_), .B(_367_), .Y(_0__30_) );
INVX1 INVX1_10 ( .A(i_add_term1[28]), .Y(_373_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[28]), .B(_373_), .Y(_374_) );
INVX1 INVX1_11 ( .A(i_add_term2[28]), .Y(_375_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term1[28]), .B(_375_), .Y(_376_) );
INVX1 INVX1_12 ( .A(i_add_term1[29]), .Y(_377_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[29]), .B(_377_), .Y(_378_) );
INVX1 INVX1_13 ( .A(i_add_term2[29]), .Y(_379_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term1[29]), .B(_379_), .Y(_380_) );
OAI22X1 OAI22X1_2 ( .A(_374_), .B(_376_), .C(_378_), .D(_380_), .Y(_381_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_382_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_383_) );
NOR2X1 NOR2X1_17 ( .A(_382_), .B(_383_), .Y(_384_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_385_) );
NAND2X1 NAND2X1_11 ( .A(_384_), .B(_385_), .Y(_386_) );
NOR2X1 NOR2X1_18 ( .A(_381_), .B(_386_), .Y(_24_) );
INVX1 INVX1_14 ( .A(_22_), .Y(_387_) );
NAND2X1 NAND2X1_12 ( .A(1'b0), .B(_24_), .Y(_388_) );
OAI21X1 OAI21X1_10 ( .A(_24_), .B(_387_), .C(_388_), .Y(w_cout_8_) );
INVX1 INVX1_15 ( .A(w_cout_8_), .Y(_393_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_394_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_395_) );
OAI21X1 OAI21X1_11 ( .A(_393_), .B(_395_), .C(_394_), .Y(_26__1_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_389_) );
NAND3X1 NAND3X1_5 ( .A(_393_), .B(_394_), .C(_389_), .Y(_390_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_391_) );
OAI21X1 OAI21X1_12 ( .A(_395_), .B(_391_), .C(w_cout_8_), .Y(_392_) );
NAND2X1 NAND2X1_14 ( .A(_392_), .B(_390_), .Y(_0__32_) );
INVX1 INVX1_16 ( .A(_26__3_), .Y(_400_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_401_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_402_) );
OAI21X1 OAI21X1_13 ( .A(_400_), .B(_402_), .C(_401_), .Y(_25_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_396_) );
NAND3X1 NAND3X1_6 ( .A(_400_), .B(_401_), .C(_396_), .Y(_397_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_398_) );
OAI21X1 OAI21X1_14 ( .A(_402_), .B(_398_), .C(_26__3_), .Y(_399_) );
NAND2X1 NAND2X1_16 ( .A(_399_), .B(_397_), .Y(_0__35_) );
INVX1 INVX1_17 ( .A(_26__1_), .Y(_407_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_408_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_409_) );
OAI21X1 OAI21X1_15 ( .A(_407_), .B(_409_), .C(_408_), .Y(_26__2_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_403_) );
NAND3X1 NAND3X1_7 ( .A(_407_), .B(_408_), .C(_403_), .Y(_404_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_405_) );
OAI21X1 OAI21X1_16 ( .A(_409_), .B(_405_), .C(_26__1_), .Y(_406_) );
NAND2X1 NAND2X1_18 ( .A(_406_), .B(_404_), .Y(_0__33_) );
INVX1 INVX1_18 ( .A(_26__2_), .Y(_414_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_415_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_416_) );
OAI21X1 OAI21X1_17 ( .A(_414_), .B(_416_), .C(_415_), .Y(_26__3_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_410_) );
NAND3X1 NAND3X1_8 ( .A(_414_), .B(_415_), .C(_410_), .Y(_411_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_412_) );
OAI21X1 OAI21X1_18 ( .A(_416_), .B(_412_), .C(_26__2_), .Y(_413_) );
NAND2X1 NAND2X1_20 ( .A(_413_), .B(_411_), .Y(_0__34_) );
INVX1 INVX1_19 ( .A(i_add_term1[32]), .Y(_417_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[32]), .B(_417_), .Y(_418_) );
INVX1 INVX1_20 ( .A(i_add_term2[32]), .Y(_419_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term1[32]), .B(_419_), .Y(_420_) );
INVX1 INVX1_21 ( .A(i_add_term1[33]), .Y(_421_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[33]), .B(_421_), .Y(_422_) );
INVX1 INVX1_22 ( .A(i_add_term2[33]), .Y(_423_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term1[33]), .B(_423_), .Y(_424_) );
OAI22X1 OAI22X1_3 ( .A(_418_), .B(_420_), .C(_422_), .D(_424_), .Y(_425_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_426_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_427_) );
NOR2X1 NOR2X1_28 ( .A(_426_), .B(_427_), .Y(_428_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_429_) );
NAND2X1 NAND2X1_21 ( .A(_428_), .B(_429_), .Y(_430_) );
NOR2X1 NOR2X1_29 ( .A(_425_), .B(_430_), .Y(_27_) );
INVX1 INVX1_23 ( .A(_25_), .Y(_431_) );
NAND2X1 NAND2X1_22 ( .A(1'b0), .B(_27_), .Y(_432_) );
OAI21X1 OAI21X1_19 ( .A(_27_), .B(_431_), .C(_432_), .Y(w_cout_9_) );
INVX1 INVX1_24 ( .A(w_cout_9_), .Y(_437_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_438_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_439_) );
OAI21X1 OAI21X1_20 ( .A(_437_), .B(_439_), .C(_438_), .Y(_29__1_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_433_) );
NAND3X1 NAND3X1_9 ( .A(_437_), .B(_438_), .C(_433_), .Y(_434_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_435_) );
OAI21X1 OAI21X1_21 ( .A(_439_), .B(_435_), .C(w_cout_9_), .Y(_436_) );
NAND2X1 NAND2X1_24 ( .A(_436_), .B(_434_), .Y(_0__36_) );
INVX1 INVX1_25 ( .A(_29__3_), .Y(_444_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_445_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_446_) );
OAI21X1 OAI21X1_22 ( .A(_444_), .B(_446_), .C(_445_), .Y(_28_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_440_) );
NAND3X1 NAND3X1_10 ( .A(_444_), .B(_445_), .C(_440_), .Y(_441_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_442_) );
OAI21X1 OAI21X1_23 ( .A(_446_), .B(_442_), .C(_29__3_), .Y(_443_) );
NAND2X1 NAND2X1_26 ( .A(_443_), .B(_441_), .Y(_0__39_) );
INVX1 INVX1_26 ( .A(_29__1_), .Y(_451_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_452_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_453_) );
OAI21X1 OAI21X1_24 ( .A(_451_), .B(_453_), .C(_452_), .Y(_29__2_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_447_) );
NAND3X1 NAND3X1_11 ( .A(_451_), .B(_452_), .C(_447_), .Y(_448_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_449_) );
OAI21X1 OAI21X1_25 ( .A(_453_), .B(_449_), .C(_29__1_), .Y(_450_) );
NAND2X1 NAND2X1_28 ( .A(_450_), .B(_448_), .Y(_0__37_) );
INVX1 INVX1_27 ( .A(_29__2_), .Y(_458_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_459_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_460_) );
OAI21X1 OAI21X1_26 ( .A(_458_), .B(_460_), .C(_459_), .Y(_29__3_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_454_) );
NAND3X1 NAND3X1_12 ( .A(_458_), .B(_459_), .C(_454_), .Y(_455_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_456_) );
OAI21X1 OAI21X1_27 ( .A(_460_), .B(_456_), .C(_29__2_), .Y(_457_) );
NAND2X1 NAND2X1_30 ( .A(_457_), .B(_455_), .Y(_0__38_) );
INVX1 INVX1_28 ( .A(i_add_term1[36]), .Y(_461_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[36]), .B(_461_), .Y(_462_) );
INVX1 INVX1_29 ( .A(i_add_term2[36]), .Y(_463_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term1[36]), .B(_463_), .Y(_464_) );
INVX1 INVX1_30 ( .A(i_add_term1[37]), .Y(_465_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[37]), .B(_465_), .Y(_466_) );
INVX1 INVX1_31 ( .A(i_add_term2[37]), .Y(_467_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term1[37]), .B(_467_), .Y(_468_) );
OAI22X1 OAI22X1_4 ( .A(_462_), .B(_464_), .C(_466_), .D(_468_), .Y(_469_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_470_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_471_) );
NOR2X1 NOR2X1_39 ( .A(_470_), .B(_471_), .Y(_472_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_473_) );
NAND2X1 NAND2X1_31 ( .A(_472_), .B(_473_), .Y(_474_) );
NOR2X1 NOR2X1_40 ( .A(_469_), .B(_474_), .Y(_30_) );
INVX1 INVX1_32 ( .A(_28_), .Y(_475_) );
NAND2X1 NAND2X1_32 ( .A(1'b0), .B(_30_), .Y(_476_) );
OAI21X1 OAI21X1_28 ( .A(_30_), .B(_475_), .C(_476_), .Y(w_cout_10_) );
INVX1 INVX1_33 ( .A(w_cout_10_), .Y(_481_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_482_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_483_) );
OAI21X1 OAI21X1_29 ( .A(_481_), .B(_483_), .C(_482_), .Y(_32__1_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_477_) );
NAND3X1 NAND3X1_13 ( .A(_481_), .B(_482_), .C(_477_), .Y(_478_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_479_) );
OAI21X1 OAI21X1_30 ( .A(_483_), .B(_479_), .C(w_cout_10_), .Y(_480_) );
NAND2X1 NAND2X1_34 ( .A(_480_), .B(_478_), .Y(_0__40_) );
INVX1 INVX1_34 ( .A(_32__3_), .Y(_488_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_489_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_490_) );
OAI21X1 OAI21X1_31 ( .A(_488_), .B(_490_), .C(_489_), .Y(_31_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_484_) );
NAND3X1 NAND3X1_14 ( .A(_488_), .B(_489_), .C(_484_), .Y(_485_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_486_) );
OAI21X1 OAI21X1_32 ( .A(_490_), .B(_486_), .C(_32__3_), .Y(_487_) );
NAND2X1 NAND2X1_36 ( .A(_487_), .B(_485_), .Y(_0__43_) );
INVX1 INVX1_35 ( .A(_32__1_), .Y(_495_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_496_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_497_) );
OAI21X1 OAI21X1_33 ( .A(_495_), .B(_497_), .C(_496_), .Y(_32__2_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_491_) );
NAND3X1 NAND3X1_15 ( .A(_495_), .B(_496_), .C(_491_), .Y(_492_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_493_) );
OAI21X1 OAI21X1_34 ( .A(_497_), .B(_493_), .C(_32__1_), .Y(_494_) );
NAND2X1 NAND2X1_38 ( .A(_494_), .B(_492_), .Y(_0__41_) );
INVX1 INVX1_36 ( .A(_32__2_), .Y(_502_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_503_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_504_) );
OAI21X1 OAI21X1_35 ( .A(_502_), .B(_504_), .C(_503_), .Y(_32__3_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_498_) );
NAND3X1 NAND3X1_16 ( .A(_502_), .B(_503_), .C(_498_), .Y(_499_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_500_) );
OAI21X1 OAI21X1_36 ( .A(_504_), .B(_500_), .C(_32__2_), .Y(_501_) );
NAND2X1 NAND2X1_40 ( .A(_501_), .B(_499_), .Y(_0__42_) );
INVX1 INVX1_37 ( .A(i_add_term1[40]), .Y(_505_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[40]), .B(_505_), .Y(_506_) );
INVX1 INVX1_38 ( .A(i_add_term2[40]), .Y(_507_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term1[40]), .B(_507_), .Y(_508_) );
INVX1 INVX1_39 ( .A(i_add_term1[41]), .Y(_509_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[41]), .B(_509_), .Y(_510_) );
INVX1 INVX1_40 ( .A(i_add_term2[41]), .Y(_511_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term1[41]), .B(_511_), .Y(_512_) );
OAI22X1 OAI22X1_5 ( .A(_506_), .B(_508_), .C(_510_), .D(_512_), .Y(_513_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_514_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_515_) );
NOR2X1 NOR2X1_50 ( .A(_514_), .B(_515_), .Y(_516_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_517_) );
NAND2X1 NAND2X1_41 ( .A(_516_), .B(_517_), .Y(_518_) );
NOR2X1 NOR2X1_51 ( .A(_513_), .B(_518_), .Y(_33_) );
INVX1 INVX1_41 ( .A(_31_), .Y(_519_) );
NAND2X1 NAND2X1_42 ( .A(1'b0), .B(_33_), .Y(_520_) );
OAI21X1 OAI21X1_37 ( .A(_33_), .B(_519_), .C(_520_), .Y(w_cout_11_) );
INVX1 INVX1_42 ( .A(w_cout_11_), .Y(_525_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_526_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_527_) );
OAI21X1 OAI21X1_38 ( .A(_525_), .B(_527_), .C(_526_), .Y(_35__1_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_521_) );
NAND3X1 NAND3X1_17 ( .A(_525_), .B(_526_), .C(_521_), .Y(_522_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_523_) );
OAI21X1 OAI21X1_39 ( .A(_527_), .B(_523_), .C(w_cout_11_), .Y(_524_) );
NAND2X1 NAND2X1_44 ( .A(_524_), .B(_522_), .Y(_0__44_) );
INVX1 INVX1_43 ( .A(_35__3_), .Y(_532_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_533_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_534_) );
OAI21X1 OAI21X1_40 ( .A(_532_), .B(_534_), .C(_533_), .Y(_34_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_528_) );
NAND3X1 NAND3X1_18 ( .A(_532_), .B(_533_), .C(_528_), .Y(_529_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_530_) );
OAI21X1 OAI21X1_41 ( .A(_534_), .B(_530_), .C(_35__3_), .Y(_531_) );
NAND2X1 NAND2X1_46 ( .A(_531_), .B(_529_), .Y(_0__47_) );
INVX1 INVX1_44 ( .A(_35__1_), .Y(_539_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_540_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_541_) );
OAI21X1 OAI21X1_42 ( .A(_539_), .B(_541_), .C(_540_), .Y(_35__2_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_535_) );
NAND3X1 NAND3X1_19 ( .A(_539_), .B(_540_), .C(_535_), .Y(_536_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_537_) );
OAI21X1 OAI21X1_43 ( .A(_541_), .B(_537_), .C(_35__1_), .Y(_538_) );
NAND2X1 NAND2X1_48 ( .A(_538_), .B(_536_), .Y(_0__45_) );
INVX1 INVX1_45 ( .A(_35__2_), .Y(_546_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_547_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_548_) );
OAI21X1 OAI21X1_44 ( .A(_546_), .B(_548_), .C(_547_), .Y(_35__3_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_542_) );
NAND3X1 NAND3X1_20 ( .A(_546_), .B(_547_), .C(_542_), .Y(_543_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_544_) );
OAI21X1 OAI21X1_45 ( .A(_548_), .B(_544_), .C(_35__2_), .Y(_545_) );
NAND2X1 NAND2X1_50 ( .A(_545_), .B(_543_), .Y(_0__46_) );
INVX1 INVX1_46 ( .A(i_add_term1[44]), .Y(_549_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[44]), .B(_549_), .Y(_550_) );
INVX1 INVX1_47 ( .A(i_add_term2[44]), .Y(_551_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term1[44]), .B(_551_), .Y(_552_) );
INVX1 INVX1_48 ( .A(i_add_term1[45]), .Y(_553_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[45]), .B(_553_), .Y(_554_) );
INVX1 INVX1_49 ( .A(i_add_term2[45]), .Y(_555_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term1[45]), .B(_555_), .Y(_556_) );
OAI22X1 OAI22X1_6 ( .A(_550_), .B(_552_), .C(_554_), .D(_556_), .Y(_557_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_558_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_559_) );
NOR2X1 NOR2X1_61 ( .A(_558_), .B(_559_), .Y(_560_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_561_) );
NAND2X1 NAND2X1_51 ( .A(_560_), .B(_561_), .Y(_562_) );
NOR2X1 NOR2X1_62 ( .A(_557_), .B(_562_), .Y(_36_) );
INVX1 INVX1_50 ( .A(_34_), .Y(_563_) );
NAND2X1 NAND2X1_52 ( .A(1'b0), .B(_36_), .Y(_564_) );
OAI21X1 OAI21X1_46 ( .A(_36_), .B(_563_), .C(_564_), .Y(cskip2_inst_cin) );
INVX1 INVX1_51 ( .A(cskip2_inst_cin), .Y(_569_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_570_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_571_) );
OAI21X1 OAI21X1_47 ( .A(_569_), .B(_571_), .C(_570_), .Y(cskip2_inst_rca0_c) );
OR2X2 OR2X2_21 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_565_) );
NAND3X1 NAND3X1_21 ( .A(_569_), .B(_570_), .C(_565_), .Y(_566_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_567_) );
OAI21X1 OAI21X1_48 ( .A(_571_), .B(_567_), .C(cskip2_inst_cin), .Y(_568_) );
NAND2X1 NAND2X1_54 ( .A(_568_), .B(_566_), .Y(cskip2_inst_rca0_fa0_o_sum) );
INVX1 INVX1_52 ( .A(cskip2_inst_rca0_c), .Y(_576_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_577_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_578_) );
OAI21X1 OAI21X1_49 ( .A(_576_), .B(_578_), .C(_577_), .Y(cskip2_inst_cout0) );
OR2X2 OR2X2_22 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_572_) );
NAND3X1 NAND3X1_22 ( .A(_576_), .B(_577_), .C(_572_), .Y(_573_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_574_) );
OAI21X1 OAI21X1_50 ( .A(_578_), .B(_574_), .C(cskip2_inst_rca0_c), .Y(_575_) );
NAND2X1 NAND2X1_56 ( .A(_575_), .B(_573_), .Y(cskip2_inst_rca0_fa31_o_sum) );
INVX1 INVX1_53 ( .A(i_add_term1[49]), .Y(_583_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[49]), .B(_583_), .Y(_584_) );
INVX1 INVX1_54 ( .A(i_add_term2[49]), .Y(_585_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term1[49]), .B(_585_), .Y(_586_) );
INVX1 INVX1_55 ( .A(i_add_term1[48]), .Y(_579_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[48]), .B(_579_), .Y(_580_) );
INVX1 INVX1_56 ( .A(i_add_term2[48]), .Y(_581_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term1[48]), .B(_581_), .Y(_582_) );
AOI22X1 AOI22X1_1 ( .A(_584_), .B(_586_), .C(_580_), .D(_582_), .Y(cskip2_inst_skip0_P) );
INVX1 INVX1_57 ( .A(cskip2_inst_cout0), .Y(_587_) );
NAND2X1 NAND2X1_61 ( .A(1'b0), .B(cskip2_inst_skip0_P), .Y(_588_) );
OAI21X1 OAI21X1_51 ( .A(cskip2_inst_skip0_P), .B(_587_), .C(_588_), .Y(w_cout_13_) );
BUFX2 BUFX2_1 ( .A(w_cout_13_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(cskip2_inst_rca0_fa0_o_sum), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(cskip2_inst_rca0_fa31_o_sum), .Y(sum[49]) );
INVX1 INVX1_58 ( .A(1'b0), .Y(_41_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_42_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_43_) );
OAI21X1 OAI21X1_52 ( .A(_41_), .B(_43_), .C(_42_), .Y(_2__1_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_37_) );
NAND3X1 NAND3X1_23 ( .A(_41_), .B(_42_), .C(_37_), .Y(_38_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_39_) );
OAI21X1 OAI21X1_53 ( .A(_43_), .B(_39_), .C(1'b0), .Y(_40_) );
NAND2X1 NAND2X1_63 ( .A(_40_), .B(_38_), .Y(_0__0_) );
INVX1 INVX1_59 ( .A(_2__3_), .Y(_48_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_49_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_50_) );
OAI21X1 OAI21X1_54 ( .A(_48_), .B(_50_), .C(_49_), .Y(_1_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_44_) );
NAND3X1 NAND3X1_24 ( .A(_48_), .B(_49_), .C(_44_), .Y(_45_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_46_) );
OAI21X1 OAI21X1_55 ( .A(_50_), .B(_46_), .C(_2__3_), .Y(_47_) );
NAND2X1 NAND2X1_65 ( .A(_47_), .B(_45_), .Y(_0__3_) );
INVX1 INVX1_60 ( .A(_2__1_), .Y(_55_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_56_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_57_) );
OAI21X1 OAI21X1_56 ( .A(_55_), .B(_57_), .C(_56_), .Y(_2__2_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_51_) );
NAND3X1 NAND3X1_25 ( .A(_55_), .B(_56_), .C(_51_), .Y(_52_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_53_) );
OAI21X1 OAI21X1_57 ( .A(_57_), .B(_53_), .C(_2__1_), .Y(_54_) );
NAND2X1 NAND2X1_67 ( .A(_54_), .B(_52_), .Y(_0__1_) );
INVX1 INVX1_61 ( .A(_2__2_), .Y(_62_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_63_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_64_) );
OAI21X1 OAI21X1_58 ( .A(_62_), .B(_64_), .C(_63_), .Y(_2__3_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_58_) );
NAND3X1 NAND3X1_26 ( .A(_62_), .B(_63_), .C(_58_), .Y(_59_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_60_) );
OAI21X1 OAI21X1_59 ( .A(_64_), .B(_60_), .C(_2__2_), .Y(_61_) );
NAND2X1 NAND2X1_69 ( .A(_61_), .B(_59_), .Y(_0__2_) );
INVX1 INVX1_62 ( .A(i_add_term1[0]), .Y(_65_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[0]), .B(_65_), .Y(_66_) );
INVX1 INVX1_63 ( .A(i_add_term2[0]), .Y(_67_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term1[0]), .B(_67_), .Y(_68_) );
INVX1 INVX1_64 ( .A(i_add_term1[1]), .Y(_69_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[1]), .B(_69_), .Y(_70_) );
INVX1 INVX1_65 ( .A(i_add_term2[1]), .Y(_71_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term1[1]), .B(_71_), .Y(_72_) );
OAI22X1 OAI22X1_7 ( .A(_66_), .B(_68_), .C(_70_), .D(_72_), .Y(_73_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_74_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_75_) );
NOR2X1 NOR2X1_74 ( .A(_74_), .B(_75_), .Y(_76_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_77_) );
NAND2X1 NAND2X1_70 ( .A(_76_), .B(_77_), .Y(_78_) );
NOR2X1 NOR2X1_75 ( .A(_73_), .B(_78_), .Y(_3_) );
INVX1 INVX1_66 ( .A(_1_), .Y(_79_) );
NAND2X1 NAND2X1_71 ( .A(1'b0), .B(_3_), .Y(_80_) );
OAI21X1 OAI21X1_60 ( .A(_3_), .B(_79_), .C(_80_), .Y(w_cout_1_) );
INVX1 INVX1_67 ( .A(w_cout_1_), .Y(_85_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_86_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_87_) );
OAI21X1 OAI21X1_61 ( .A(_85_), .B(_87_), .C(_86_), .Y(_5__1_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_81_) );
NAND3X1 NAND3X1_27 ( .A(_85_), .B(_86_), .C(_81_), .Y(_82_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_83_) );
OAI21X1 OAI21X1_62 ( .A(_87_), .B(_83_), .C(w_cout_1_), .Y(_84_) );
NAND2X1 NAND2X1_73 ( .A(_84_), .B(_82_), .Y(_0__4_) );
INVX1 INVX1_68 ( .A(_5__3_), .Y(_92_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_93_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_94_) );
OAI21X1 OAI21X1_63 ( .A(_92_), .B(_94_), .C(_93_), .Y(_4_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_88_) );
NAND3X1 NAND3X1_28 ( .A(_92_), .B(_93_), .C(_88_), .Y(_89_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_90_) );
OAI21X1 OAI21X1_64 ( .A(_94_), .B(_90_), .C(_5__3_), .Y(_91_) );
NAND2X1 NAND2X1_75 ( .A(_91_), .B(_89_), .Y(_0__7_) );
INVX1 INVX1_69 ( .A(_5__1_), .Y(_99_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_100_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_101_) );
OAI21X1 OAI21X1_65 ( .A(_99_), .B(_101_), .C(_100_), .Y(_5__2_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_95_) );
NAND3X1 NAND3X1_29 ( .A(_99_), .B(_100_), .C(_95_), .Y(_96_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_97_) );
OAI21X1 OAI21X1_66 ( .A(_101_), .B(_97_), .C(_5__1_), .Y(_98_) );
NAND2X1 NAND2X1_77 ( .A(_98_), .B(_96_), .Y(_0__5_) );
INVX1 INVX1_70 ( .A(_5__2_), .Y(_106_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_107_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_108_) );
OAI21X1 OAI21X1_67 ( .A(_106_), .B(_108_), .C(_107_), .Y(_5__3_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_102_) );
NAND3X1 NAND3X1_30 ( .A(_106_), .B(_107_), .C(_102_), .Y(_103_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_104_) );
OAI21X1 OAI21X1_68 ( .A(_108_), .B(_104_), .C(_5__2_), .Y(_105_) );
NAND2X1 NAND2X1_79 ( .A(_105_), .B(_103_), .Y(_0__6_) );
INVX1 INVX1_71 ( .A(i_add_term1[4]), .Y(_109_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[4]), .B(_109_), .Y(_110_) );
INVX1 INVX1_72 ( .A(i_add_term2[4]), .Y(_111_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term1[4]), .B(_111_), .Y(_112_) );
INVX1 INVX1_73 ( .A(i_add_term1[5]), .Y(_113_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[5]), .B(_113_), .Y(_114_) );
INVX1 INVX1_74 ( .A(i_add_term2[5]), .Y(_115_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term1[5]), .B(_115_), .Y(_116_) );
OAI22X1 OAI22X1_8 ( .A(_110_), .B(_112_), .C(_114_), .D(_116_), .Y(_117_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_118_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_119_) );
NOR2X1 NOR2X1_85 ( .A(_118_), .B(_119_), .Y(_120_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_121_) );
NAND2X1 NAND2X1_80 ( .A(_120_), .B(_121_), .Y(_122_) );
NOR2X1 NOR2X1_86 ( .A(_117_), .B(_122_), .Y(_6_) );
INVX1 INVX1_75 ( .A(_4_), .Y(_123_) );
NAND2X1 NAND2X1_81 ( .A(1'b0), .B(_6_), .Y(_124_) );
OAI21X1 OAI21X1_69 ( .A(_6_), .B(_123_), .C(_124_), .Y(w_cout_2_) );
INVX1 INVX1_76 ( .A(w_cout_2_), .Y(_129_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_130_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_131_) );
OAI21X1 OAI21X1_70 ( .A(_129_), .B(_131_), .C(_130_), .Y(_8__1_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_125_) );
NAND3X1 NAND3X1_31 ( .A(_129_), .B(_130_), .C(_125_), .Y(_126_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_127_) );
OAI21X1 OAI21X1_71 ( .A(_131_), .B(_127_), .C(w_cout_2_), .Y(_128_) );
NAND2X1 NAND2X1_83 ( .A(_128_), .B(_126_), .Y(_0__8_) );
INVX1 INVX1_77 ( .A(_8__3_), .Y(_136_) );
NAND2X1 NAND2X1_84 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_137_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_138_) );
OAI21X1 OAI21X1_72 ( .A(_136_), .B(_138_), .C(_137_), .Y(_7_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_132_) );
NAND3X1 NAND3X1_32 ( .A(_136_), .B(_137_), .C(_132_), .Y(_133_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_134_) );
OAI21X1 OAI21X1_73 ( .A(_138_), .B(_134_), .C(_8__3_), .Y(_135_) );
NAND2X1 NAND2X1_85 ( .A(_135_), .B(_133_), .Y(_0__11_) );
INVX1 INVX1_78 ( .A(_8__1_), .Y(_143_) );
NAND2X1 NAND2X1_86 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_144_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_145_) );
OAI21X1 OAI21X1_74 ( .A(_143_), .B(_145_), .C(_144_), .Y(_8__2_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_139_) );
NAND3X1 NAND3X1_33 ( .A(_143_), .B(_144_), .C(_139_), .Y(_140_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_141_) );
OAI21X1 OAI21X1_75 ( .A(_145_), .B(_141_), .C(_8__1_), .Y(_142_) );
NAND2X1 NAND2X1_87 ( .A(_142_), .B(_140_), .Y(_0__9_) );
INVX1 INVX1_79 ( .A(_8__2_), .Y(_150_) );
NAND2X1 NAND2X1_88 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_151_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_152_) );
OAI21X1 OAI21X1_76 ( .A(_150_), .B(_152_), .C(_151_), .Y(_8__3_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_146_) );
NAND3X1 NAND3X1_34 ( .A(_150_), .B(_151_), .C(_146_), .Y(_147_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_148_) );
OAI21X1 OAI21X1_77 ( .A(_152_), .B(_148_), .C(_8__2_), .Y(_149_) );
NAND2X1 NAND2X1_89 ( .A(_149_), .B(_147_), .Y(_0__10_) );
INVX1 INVX1_80 ( .A(i_add_term1[8]), .Y(_153_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[8]), .B(_153_), .Y(_154_) );
INVX1 INVX1_81 ( .A(i_add_term2[8]), .Y(_155_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term1[8]), .B(_155_), .Y(_156_) );
INVX1 INVX1_82 ( .A(i_add_term1[9]), .Y(_157_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[9]), .B(_157_), .Y(_158_) );
INVX1 INVX1_83 ( .A(i_add_term2[9]), .Y(_159_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term1[9]), .B(_159_), .Y(_160_) );
OAI22X1 OAI22X1_9 ( .A(_154_), .B(_156_), .C(_158_), .D(_160_), .Y(_161_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_162_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_163_) );
NOR2X1 NOR2X1_96 ( .A(_162_), .B(_163_), .Y(_164_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_165_) );
NAND2X1 NAND2X1_90 ( .A(_164_), .B(_165_), .Y(_166_) );
NOR2X1 NOR2X1_97 ( .A(_161_), .B(_166_), .Y(_9_) );
INVX1 INVX1_84 ( .A(_7_), .Y(_167_) );
NAND2X1 NAND2X1_91 ( .A(1'b0), .B(_9_), .Y(_168_) );
OAI21X1 OAI21X1_78 ( .A(_9_), .B(_167_), .C(_168_), .Y(w_cout_3_) );
INVX1 INVX1_85 ( .A(w_cout_3_), .Y(_173_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_174_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_175_) );
OAI21X1 OAI21X1_79 ( .A(_173_), .B(_175_), .C(_174_), .Y(_11__1_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_169_) );
NAND3X1 NAND3X1_35 ( .A(_173_), .B(_174_), .C(_169_), .Y(_170_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_171_) );
OAI21X1 OAI21X1_80 ( .A(_175_), .B(_171_), .C(w_cout_3_), .Y(_172_) );
NAND2X1 NAND2X1_93 ( .A(_172_), .B(_170_), .Y(_0__12_) );
INVX1 INVX1_86 ( .A(_11__3_), .Y(_180_) );
NAND2X1 NAND2X1_94 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_181_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_182_) );
OAI21X1 OAI21X1_81 ( .A(_180_), .B(_182_), .C(_181_), .Y(_10_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_176_) );
NAND3X1 NAND3X1_36 ( .A(_180_), .B(_181_), .C(_176_), .Y(_177_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_178_) );
OAI21X1 OAI21X1_82 ( .A(_182_), .B(_178_), .C(_11__3_), .Y(_179_) );
NAND2X1 NAND2X1_95 ( .A(_179_), .B(_177_), .Y(_0__15_) );
INVX1 INVX1_87 ( .A(_11__1_), .Y(_187_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_188_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_189_) );
OAI21X1 OAI21X1_83 ( .A(_187_), .B(_189_), .C(_188_), .Y(_11__2_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_183_) );
NAND3X1 NAND3X1_37 ( .A(_187_), .B(_188_), .C(_183_), .Y(_184_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_185_) );
OAI21X1 OAI21X1_84 ( .A(_189_), .B(_185_), .C(_11__1_), .Y(_186_) );
NAND2X1 NAND2X1_97 ( .A(_186_), .B(_184_), .Y(_0__13_) );
INVX1 INVX1_88 ( .A(_11__2_), .Y(_194_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_195_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_196_) );
OAI21X1 OAI21X1_85 ( .A(_194_), .B(_196_), .C(_195_), .Y(_11__3_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_190_) );
NAND3X1 NAND3X1_38 ( .A(_194_), .B(_195_), .C(_190_), .Y(_191_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_192_) );
OAI21X1 OAI21X1_86 ( .A(_196_), .B(_192_), .C(_11__2_), .Y(_193_) );
NAND2X1 NAND2X1_99 ( .A(_193_), .B(_191_), .Y(_0__14_) );
INVX1 INVX1_89 ( .A(i_add_term1[12]), .Y(_197_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[12]), .B(_197_), .Y(_198_) );
INVX1 INVX1_90 ( .A(i_add_term2[12]), .Y(_199_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term1[12]), .B(_199_), .Y(_200_) );
INVX1 INVX1_91 ( .A(i_add_term1[13]), .Y(_201_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term2[13]), .B(_201_), .Y(_202_) );
INVX1 INVX1_92 ( .A(i_add_term2[13]), .Y(_203_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term1[13]), .B(_203_), .Y(_204_) );
OAI22X1 OAI22X1_10 ( .A(_198_), .B(_200_), .C(_202_), .D(_204_), .Y(_205_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_206_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_207_) );
NOR2X1 NOR2X1_107 ( .A(_206_), .B(_207_), .Y(_208_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_209_) );
NAND2X1 NAND2X1_100 ( .A(_208_), .B(_209_), .Y(_210_) );
NOR2X1 NOR2X1_108 ( .A(_205_), .B(_210_), .Y(_12_) );
INVX1 INVX1_93 ( .A(_10_), .Y(_211_) );
NAND2X1 NAND2X1_101 ( .A(1'b0), .B(_12_), .Y(_212_) );
OAI21X1 OAI21X1_87 ( .A(_12_), .B(_211_), .C(_212_), .Y(w_cout_4_) );
INVX1 INVX1_94 ( .A(w_cout_4_), .Y(_217_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_218_) );
NOR2X1 NOR2X1_109 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_219_) );
OAI21X1 OAI21X1_88 ( .A(_217_), .B(_219_), .C(_218_), .Y(_14__1_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_213_) );
NAND3X1 NAND3X1_39 ( .A(_217_), .B(_218_), .C(_213_), .Y(_214_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_215_) );
OAI21X1 OAI21X1_89 ( .A(_219_), .B(_215_), .C(w_cout_4_), .Y(_216_) );
NAND2X1 NAND2X1_103 ( .A(_216_), .B(_214_), .Y(_0__16_) );
INVX1 INVX1_95 ( .A(_14__3_), .Y(_224_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_225_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_226_) );
OAI21X1 OAI21X1_90 ( .A(_224_), .B(_226_), .C(_225_), .Y(_13_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_220_) );
NAND3X1 NAND3X1_40 ( .A(_224_), .B(_225_), .C(_220_), .Y(_221_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_222_) );
OAI21X1 OAI21X1_91 ( .A(_226_), .B(_222_), .C(_14__3_), .Y(_223_) );
NAND2X1 NAND2X1_105 ( .A(_223_), .B(_221_), .Y(_0__19_) );
INVX1 INVX1_96 ( .A(_14__1_), .Y(_231_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_232_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_233_) );
OAI21X1 OAI21X1_92 ( .A(_231_), .B(_233_), .C(_232_), .Y(_14__2_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_227_) );
NAND3X1 NAND3X1_41 ( .A(_231_), .B(_232_), .C(_227_), .Y(_228_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_229_) );
OAI21X1 OAI21X1_93 ( .A(_233_), .B(_229_), .C(_14__1_), .Y(_230_) );
NAND2X1 NAND2X1_107 ( .A(_230_), .B(_228_), .Y(_0__17_) );
INVX1 INVX1_97 ( .A(_14__2_), .Y(_238_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_239_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_240_) );
OAI21X1 OAI21X1_94 ( .A(_238_), .B(_240_), .C(_239_), .Y(_14__3_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_234_) );
NAND3X1 NAND3X1_42 ( .A(_238_), .B(_239_), .C(_234_), .Y(_235_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_236_) );
OAI21X1 OAI21X1_95 ( .A(_240_), .B(_236_), .C(_14__2_), .Y(_237_) );
NAND2X1 NAND2X1_109 ( .A(_237_), .B(_235_), .Y(_0__18_) );
INVX1 INVX1_98 ( .A(i_add_term1[16]), .Y(_241_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term2[16]), .B(_241_), .Y(_242_) );
INVX1 INVX1_99 ( .A(i_add_term2[16]), .Y(_243_) );
NOR2X1 NOR2X1_114 ( .A(i_add_term1[16]), .B(_243_), .Y(_244_) );
INVX1 INVX1_100 ( .A(i_add_term1[17]), .Y(_245_) );
NOR2X1 NOR2X1_115 ( .A(i_add_term2[17]), .B(_245_), .Y(_246_) );
INVX1 INVX1_101 ( .A(i_add_term2[17]), .Y(_247_) );
NOR2X1 NOR2X1_116 ( .A(i_add_term1[17]), .B(_247_), .Y(_248_) );
OAI22X1 OAI22X1_11 ( .A(_242_), .B(_244_), .C(_246_), .D(_248_), .Y(_249_) );
NOR2X1 NOR2X1_117 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_250_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_251_) );
NOR2X1 NOR2X1_118 ( .A(_250_), .B(_251_), .Y(_252_) );
XOR2X1 XOR2X1_11 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_253_) );
NAND2X1 NAND2X1_110 ( .A(_252_), .B(_253_), .Y(_254_) );
NOR2X1 NOR2X1_119 ( .A(_249_), .B(_254_), .Y(_15_) );
INVX1 INVX1_102 ( .A(_13_), .Y(_255_) );
NAND2X1 NAND2X1_111 ( .A(1'b0), .B(_15_), .Y(_256_) );
OAI21X1 OAI21X1_96 ( .A(_15_), .B(_255_), .C(_256_), .Y(w_cout_5_) );
INVX1 INVX1_103 ( .A(w_cout_5_), .Y(_261_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_262_) );
NOR2X1 NOR2X1_120 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_263_) );
OAI21X1 OAI21X1_97 ( .A(_261_), .B(_263_), .C(_262_), .Y(_17__1_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_257_) );
NAND3X1 NAND3X1_43 ( .A(_261_), .B(_262_), .C(_257_), .Y(_258_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_259_) );
OAI21X1 OAI21X1_98 ( .A(_263_), .B(_259_), .C(w_cout_5_), .Y(_260_) );
NAND2X1 NAND2X1_113 ( .A(_260_), .B(_258_), .Y(_0__20_) );
INVX1 INVX1_104 ( .A(_17__3_), .Y(_268_) );
NAND2X1 NAND2X1_114 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_269_) );
NOR2X1 NOR2X1_121 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_270_) );
OAI21X1 OAI21X1_99 ( .A(_268_), .B(_270_), .C(_269_), .Y(_16_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_264_) );
NAND3X1 NAND3X1_44 ( .A(_268_), .B(_269_), .C(_264_), .Y(_265_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_266_) );
OAI21X1 OAI21X1_100 ( .A(_270_), .B(_266_), .C(_17__3_), .Y(_267_) );
NAND2X1 NAND2X1_115 ( .A(_267_), .B(_265_), .Y(_0__23_) );
INVX1 INVX1_105 ( .A(_17__1_), .Y(_275_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_276_) );
NOR2X1 NOR2X1_122 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_277_) );
OAI21X1 OAI21X1_101 ( .A(_275_), .B(_277_), .C(_276_), .Y(_17__2_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_271_) );
NAND3X1 NAND3X1_45 ( .A(_275_), .B(_276_), .C(_271_), .Y(_272_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_273_) );
OAI21X1 OAI21X1_102 ( .A(_277_), .B(_273_), .C(_17__1_), .Y(_274_) );
NAND2X1 NAND2X1_117 ( .A(_274_), .B(_272_), .Y(_0__21_) );
INVX1 INVX1_106 ( .A(_17__2_), .Y(_282_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_283_) );
NOR2X1 NOR2X1_123 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_284_) );
OAI21X1 OAI21X1_103 ( .A(_282_), .B(_284_), .C(_283_), .Y(_17__3_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_278_) );
NAND3X1 NAND3X1_46 ( .A(_282_), .B(_283_), .C(_278_), .Y(_279_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_280_) );
OAI21X1 OAI21X1_104 ( .A(_284_), .B(_280_), .C(_17__2_), .Y(_281_) );
NAND2X1 NAND2X1_119 ( .A(_281_), .B(_279_), .Y(_0__22_) );
INVX1 INVX1_107 ( .A(i_add_term1[20]), .Y(_285_) );
NOR2X1 NOR2X1_124 ( .A(i_add_term2[20]), .B(_285_), .Y(_286_) );
INVX1 INVX1_108 ( .A(i_add_term2[20]), .Y(_287_) );
NOR2X1 NOR2X1_125 ( .A(i_add_term1[20]), .B(_287_), .Y(_288_) );
INVX1 INVX1_109 ( .A(i_add_term1[21]), .Y(_289_) );
NOR2X1 NOR2X1_126 ( .A(i_add_term2[21]), .B(_289_), .Y(_290_) );
INVX1 INVX1_110 ( .A(i_add_term2[21]), .Y(_291_) );
NOR2X1 NOR2X1_127 ( .A(i_add_term1[21]), .B(_291_), .Y(_292_) );
OAI22X1 OAI22X1_12 ( .A(_286_), .B(_288_), .C(_290_), .D(_292_), .Y(_293_) );
NOR2X1 NOR2X1_128 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_294_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_295_) );
NOR2X1 NOR2X1_129 ( .A(_294_), .B(_295_), .Y(_296_) );
XOR2X1 XOR2X1_12 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_297_) );
NAND2X1 NAND2X1_120 ( .A(_296_), .B(_297_), .Y(_298_) );
NOR2X1 NOR2X1_130 ( .A(_293_), .B(_298_), .Y(_18_) );
INVX1 INVX1_111 ( .A(_16_), .Y(_299_) );
NAND2X1 NAND2X1_121 ( .A(1'b0), .B(_18_), .Y(_300_) );
OAI21X1 OAI21X1_105 ( .A(_18_), .B(_299_), .C(_300_), .Y(w_cout_6_) );
INVX1 INVX1_112 ( .A(w_cout_6_), .Y(_305_) );
NAND2X1 NAND2X1_122 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_306_) );
NOR2X1 NOR2X1_131 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_307_) );
OAI21X1 OAI21X1_106 ( .A(_305_), .B(_307_), .C(_306_), .Y(_20__1_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_301_) );
NAND3X1 NAND3X1_47 ( .A(_305_), .B(_306_), .C(_301_), .Y(_302_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_303_) );
OAI21X1 OAI21X1_107 ( .A(_307_), .B(_303_), .C(w_cout_6_), .Y(_304_) );
NAND2X1 NAND2X1_123 ( .A(_304_), .B(_302_), .Y(_0__24_) );
INVX1 INVX1_113 ( .A(_20__3_), .Y(_312_) );
NAND2X1 NAND2X1_124 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_313_) );
NOR2X1 NOR2X1_132 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_314_) );
OAI21X1 OAI21X1_108 ( .A(_312_), .B(_314_), .C(_313_), .Y(_19_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_308_) );
NAND3X1 NAND3X1_48 ( .A(_312_), .B(_313_), .C(_308_), .Y(_309_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_310_) );
OAI21X1 OAI21X1_109 ( .A(_314_), .B(_310_), .C(_20__3_), .Y(_311_) );
NAND2X1 NAND2X1_125 ( .A(_311_), .B(_309_), .Y(_0__27_) );
INVX1 INVX1_114 ( .A(_20__1_), .Y(_319_) );
NAND2X1 NAND2X1_126 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_320_) );
NOR2X1 NOR2X1_133 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_321_) );
OAI21X1 OAI21X1_110 ( .A(_319_), .B(_321_), .C(_320_), .Y(_20__2_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_315_) );
NAND3X1 NAND3X1_49 ( .A(_319_), .B(_320_), .C(_315_), .Y(_316_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_317_) );
OAI21X1 OAI21X1_111 ( .A(_321_), .B(_317_), .C(_20__1_), .Y(_318_) );
NAND2X1 NAND2X1_127 ( .A(_318_), .B(_316_), .Y(_0__25_) );
INVX1 INVX1_115 ( .A(_20__2_), .Y(_326_) );
NAND2X1 NAND2X1_128 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_327_) );
NOR2X1 NOR2X1_134 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_328_) );
OAI21X1 OAI21X1_112 ( .A(_326_), .B(_328_), .C(_327_), .Y(_20__3_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_322_) );
NAND3X1 NAND3X1_50 ( .A(_326_), .B(_327_), .C(_322_), .Y(_323_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_324_) );
OAI21X1 OAI21X1_113 ( .A(_328_), .B(_324_), .C(_20__2_), .Y(_325_) );
NAND2X1 NAND2X1_129 ( .A(_325_), .B(_323_), .Y(_0__26_) );
BUFX2 BUFX2_52 ( .A(cskip2_inst_rca0_fa0_o_sum), .Y(_0__48_) );
BUFX2 BUFX2_53 ( .A(cskip2_inst_rca0_fa31_o_sum), .Y(_0__49_) );
BUFX2 BUFX2_54 ( .A(1'b0), .Y(w_cout_0_) );
BUFX2 BUFX2_55 ( .A(cskip2_inst_cin), .Y(w_cout_12_) );
endmodule
