module csa_7bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [6:0] i_add_term1;
input [6:0] i_add_term2;
output [6:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

INVX1 INVX1_1 ( .A(gnd), .Y(_13_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_14_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_15_) );
NAND3X1 NAND3X1_1 ( .A(_13_), .B(_15_), .C(_14_), .Y(_16_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_10_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_11_) );
OAI21X1 OAI21X1_1 ( .A(_10_), .B(_11_), .C(gnd), .Y(_12_) );
NAND2X1 NAND2X1_2 ( .A(_12_), .B(_16_), .Y(csa_inst_rca0_0_fa0_o_sum) );
OAI21X1 OAI21X1_2 ( .A(_13_), .B(_10_), .C(_15_), .Y(csa_inst_rca0_0_fa0_o_carry) );
INVX1 INVX1_2 ( .A(csa_inst_rca0_0_fa0_o_carry), .Y(_20_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_21_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_22_) );
NAND3X1 NAND3X1_2 ( .A(_20_), .B(_22_), .C(_21_), .Y(_23_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_17_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_18_) );
OAI21X1 OAI21X1_3 ( .A(_17_), .B(_18_), .C(csa_inst_rca0_0_fa0_o_carry), .Y(_19_) );
NAND2X1 NAND2X1_4 ( .A(_19_), .B(_23_), .Y(csa_inst_rca0_0_fa1_o_sum) );
OAI21X1 OAI21X1_4 ( .A(_20_), .B(_17_), .C(_22_), .Y(csa_inst_rca0_0_fa1_o_carry) );
INVX1 INVX1_3 ( .A(csa_inst_rca0_0_fa1_o_carry), .Y(_27_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_28_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_29_) );
NAND3X1 NAND3X1_3 ( .A(_27_), .B(_29_), .C(_28_), .Y(_30_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_24_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_25_) );
OAI21X1 OAI21X1_5 ( .A(_24_), .B(_25_), .C(csa_inst_rca0_0_fa1_o_carry), .Y(_26_) );
NAND2X1 NAND2X1_6 ( .A(_26_), .B(_30_), .Y(csa_inst_rca0_0_fa2_o_sum) );
OAI21X1 OAI21X1_6 ( .A(_27_), .B(_24_), .C(_29_), .Y(csa_inst_cout0_0) );
INVX1 INVX1_4 ( .A(vdd), .Y(_34_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_35_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_36_) );
NAND3X1 NAND3X1_4 ( .A(_34_), .B(_36_), .C(_35_), .Y(_37_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_31_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_32_) );
OAI21X1 OAI21X1_7 ( .A(_31_), .B(_32_), .C(vdd), .Y(_33_) );
NAND2X1 NAND2X1_8 ( .A(_33_), .B(_37_), .Y(csa_inst_rca0_1_fa0_o_sum) );
OAI21X1 OAI21X1_8 ( .A(_34_), .B(_31_), .C(_36_), .Y(csa_inst_rca0_1_fa0_o_carry) );
INVX1 INVX1_5 ( .A(csa_inst_rca0_1_fa0_o_carry), .Y(_41_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_42_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_43_) );
NAND3X1 NAND3X1_5 ( .A(_41_), .B(_43_), .C(_42_), .Y(_44_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_38_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_39_) );
OAI21X1 OAI21X1_9 ( .A(_38_), .B(_39_), .C(csa_inst_rca0_1_fa0_o_carry), .Y(_40_) );
NAND2X1 NAND2X1_10 ( .A(_40_), .B(_44_), .Y(csa_inst_rca0_1_fa1_o_sum) );
OAI21X1 OAI21X1_10 ( .A(_41_), .B(_38_), .C(_43_), .Y(csa_inst_rca0_1_fa1_o_carry) );
INVX1 INVX1_6 ( .A(csa_inst_rca0_1_fa1_o_carry), .Y(_48_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_49_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_50_) );
NAND3X1 NAND3X1_6 ( .A(_48_), .B(_50_), .C(_49_), .Y(_51_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_45_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_46_) );
OAI21X1 OAI21X1_11 ( .A(_45_), .B(_46_), .C(csa_inst_rca0_1_fa1_o_carry), .Y(_47_) );
NAND2X1 NAND2X1_12 ( .A(_47_), .B(_51_), .Y(csa_inst_rca0_1_fa2_o_sum) );
OAI21X1 OAI21X1_12 ( .A(_48_), .B(_45_), .C(_50_), .Y(csa_inst_cout0_1) );
INVX1 INVX1_7 ( .A(gnd), .Y(_55_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_56_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_57_) );
NAND3X1 NAND3X1_7 ( .A(_55_), .B(_57_), .C(_56_), .Y(_58_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_52_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_53_) );
OAI21X1 OAI21X1_13 ( .A(_52_), .B(_53_), .C(gnd), .Y(_54_) );
NAND2X1 NAND2X1_14 ( .A(_54_), .B(_58_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_14 ( .A(_55_), .B(_52_), .C(_57_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_8 ( .A(rca_inst_fa3_i_carry), .Y(_62_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_63_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_64_) );
NAND3X1 NAND3X1_8 ( .A(_62_), .B(_64_), .C(_63_), .Y(_65_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_59_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_60_) );
OAI21X1 OAI21X1_15 ( .A(_59_), .B(_60_), .C(rca_inst_fa3_i_carry), .Y(_61_) );
NAND2X1 NAND2X1_16 ( .A(_61_), .B(_65_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_16 ( .A(_62_), .B(_59_), .C(_64_), .Y(csa_inst_cin) );
INVX1 INVX1_9 ( .A(rca_inst_fa0_o_carry), .Y(_69_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_70_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_71_) );
NAND3X1 NAND3X1_9 ( .A(_69_), .B(_71_), .C(_70_), .Y(_72_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_66_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_67_) );
OAI21X1 OAI21X1_17 ( .A(_66_), .B(_67_), .C(rca_inst_fa0_o_carry), .Y(_68_) );
NAND2X1 NAND2X1_18 ( .A(_68_), .B(_72_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_18 ( .A(_69_), .B(_66_), .C(_71_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_10 ( .A(rca_inst_fa_1__o_carry), .Y(_76_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_77_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_78_) );
NAND3X1 NAND3X1_10 ( .A(_76_), .B(_78_), .C(_77_), .Y(_79_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_73_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_74_) );
OAI21X1 OAI21X1_19 ( .A(_73_), .B(_74_), .C(rca_inst_fa_1__o_carry), .Y(_75_) );
NAND2X1 NAND2X1_20 ( .A(_75_), .B(_79_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_20 ( .A(_76_), .B(_73_), .C(_78_), .Y(rca_inst_fa3_i_carry) );
BUFX2 BUFX2_1 ( .A(_0_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_1__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_1__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_1__6_), .Y(sum[6]) );
INVX1 INVX1_11 ( .A(csa_inst_cout0_0), .Y(_2_) );
NAND2X1 NAND2X1_21 ( .A(csa_inst_cout0_1), .B(csa_inst_cin), .Y(_3_) );
OAI21X1 OAI21X1_21 ( .A(csa_inst_cin), .B(_2_), .C(_3_), .Y(_0_) );
INVX1 INVX1_12 ( .A(csa_inst_rca0_0_fa0_o_sum), .Y(_4_) );
NAND2X1 NAND2X1_22 ( .A(csa_inst_rca0_1_fa0_o_sum), .B(csa_inst_cin), .Y(_5_) );
OAI21X1 OAI21X1_22 ( .A(csa_inst_cin), .B(_4_), .C(_5_), .Y(_1__4_) );
INVX1 INVX1_13 ( .A(csa_inst_rca0_0_fa1_o_sum), .Y(_6_) );
NAND2X1 NAND2X1_23 ( .A(csa_inst_cin), .B(csa_inst_rca0_1_fa1_o_sum), .Y(_7_) );
OAI21X1 OAI21X1_23 ( .A(csa_inst_cin), .B(_6_), .C(_7_), .Y(_1__5_) );
INVX1 INVX1_14 ( .A(csa_inst_rca0_0_fa2_o_sum), .Y(_8_) );
NAND2X1 NAND2X1_24 ( .A(csa_inst_cin), .B(csa_inst_rca0_1_fa2_o_sum), .Y(_9_) );
OAI21X1 OAI21X1_24 ( .A(csa_inst_cin), .B(_8_), .C(_9_), .Y(_1__6_) );
BUFX2 BUFX2_9 ( .A(rca_inst_fa0_o_sum), .Y(_1__0_) );
BUFX2 BUFX2_10 ( .A(rca_inst_fa_1__o_sum), .Y(_1__1_) );
BUFX2 BUFX2_11 ( .A(rca_inst_fa_2__o_sum), .Y(_1__2_) );
BUFX2 BUFX2_12 ( .A(rca_inst_fa3_o_sum), .Y(_1__3_) );
endmodule
