module CSkipA_52bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [51:0] i_add_term1;
input [51:0] i_add_term2;
output [51:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

AND2X2 AND2X2_1 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_321_) );
OAI21X1 OAI21X1_1 ( .A(_320_), .B(_321_), .C(_11__1_), .Y(_322_) );
NAND2X1 NAND2X1_1 ( .A(_322_), .B(_326_), .Y(_0__17_) );
OAI21X1 OAI21X1_2 ( .A(_323_), .B(_320_), .C(_325_), .Y(_11__2_) );
INVX1 INVX1_1 ( .A(_11__2_), .Y(_330_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_331_) );
NAND2X1 NAND2X1_2 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_332_) );
NAND3X1 NAND3X1_1 ( .A(_330_), .B(_332_), .C(_331_), .Y(_333_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_327_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_328_) );
OAI21X1 OAI21X1_3 ( .A(_327_), .B(_328_), .C(_11__2_), .Y(_329_) );
NAND2X1 NAND2X1_3 ( .A(_329_), .B(_333_), .Y(_0__18_) );
OAI21X1 OAI21X1_4 ( .A(_330_), .B(_327_), .C(_332_), .Y(_11__3_) );
INVX1 INVX1_2 ( .A(_11__3_), .Y(_337_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_338_) );
NAND2X1 NAND2X1_4 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_339_) );
NAND3X1 NAND3X1_2 ( .A(_337_), .B(_339_), .C(_338_), .Y(_340_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_334_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_335_) );
OAI21X1 OAI21X1_5 ( .A(_334_), .B(_335_), .C(_11__3_), .Y(_336_) );
NAND2X1 NAND2X1_5 ( .A(_336_), .B(_340_), .Y(_0__19_) );
OAI21X1 OAI21X1_6 ( .A(_337_), .B(_334_), .C(_339_), .Y(_10_) );
INVX1 INVX1_3 ( .A(w_cout_4_), .Y(_344_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_345_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_346_) );
NAND3X1 NAND3X1_3 ( .A(_344_), .B(_346_), .C(_345_), .Y(_347_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_341_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_342_) );
OAI21X1 OAI21X1_7 ( .A(_341_), .B(_342_), .C(w_cout_4_), .Y(_343_) );
NAND2X1 NAND2X1_7 ( .A(_343_), .B(_347_), .Y(_0__20_) );
OAI21X1 OAI21X1_8 ( .A(_344_), .B(_341_), .C(_346_), .Y(_14__1_) );
INVX1 INVX1_4 ( .A(_14__1_), .Y(_351_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_352_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_353_) );
NAND3X1 NAND3X1_4 ( .A(_351_), .B(_353_), .C(_352_), .Y(_354_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_348_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_349_) );
OAI21X1 OAI21X1_9 ( .A(_348_), .B(_349_), .C(_14__1_), .Y(_350_) );
NAND2X1 NAND2X1_9 ( .A(_350_), .B(_354_), .Y(_0__21_) );
OAI21X1 OAI21X1_10 ( .A(_351_), .B(_348_), .C(_353_), .Y(_14__2_) );
INVX1 INVX1_5 ( .A(_14__2_), .Y(_358_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_359_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_360_) );
NAND3X1 NAND3X1_5 ( .A(_358_), .B(_360_), .C(_359_), .Y(_361_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_355_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_356_) );
OAI21X1 OAI21X1_11 ( .A(_355_), .B(_356_), .C(_14__2_), .Y(_357_) );
NAND2X1 NAND2X1_11 ( .A(_357_), .B(_361_), .Y(_0__22_) );
OAI21X1 OAI21X1_12 ( .A(_358_), .B(_355_), .C(_360_), .Y(_14__3_) );
INVX1 INVX1_6 ( .A(_14__3_), .Y(_365_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_366_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_367_) );
NAND3X1 NAND3X1_6 ( .A(_365_), .B(_367_), .C(_366_), .Y(_368_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_362_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_363_) );
OAI21X1 OAI21X1_13 ( .A(_362_), .B(_363_), .C(_14__3_), .Y(_364_) );
NAND2X1 NAND2X1_13 ( .A(_364_), .B(_368_), .Y(_0__23_) );
OAI21X1 OAI21X1_14 ( .A(_365_), .B(_362_), .C(_367_), .Y(_13_) );
INVX1 INVX1_7 ( .A(w_cout_5_), .Y(_372_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_373_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_374_) );
NAND3X1 NAND3X1_7 ( .A(_372_), .B(_374_), .C(_373_), .Y(_375_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_369_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_370_) );
OAI21X1 OAI21X1_15 ( .A(_369_), .B(_370_), .C(w_cout_5_), .Y(_371_) );
NAND2X1 NAND2X1_15 ( .A(_371_), .B(_375_), .Y(_0__24_) );
OAI21X1 OAI21X1_16 ( .A(_372_), .B(_369_), .C(_374_), .Y(_17__1_) );
INVX1 INVX1_8 ( .A(_17__1_), .Y(_379_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_380_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_381_) );
NAND3X1 NAND3X1_8 ( .A(_379_), .B(_381_), .C(_380_), .Y(_382_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_376_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_377_) );
OAI21X1 OAI21X1_17 ( .A(_376_), .B(_377_), .C(_17__1_), .Y(_378_) );
NAND2X1 NAND2X1_17 ( .A(_378_), .B(_382_), .Y(_0__25_) );
OAI21X1 OAI21X1_18 ( .A(_379_), .B(_376_), .C(_381_), .Y(_17__2_) );
INVX1 INVX1_9 ( .A(_17__2_), .Y(_386_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_387_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_388_) );
NAND3X1 NAND3X1_9 ( .A(_386_), .B(_388_), .C(_387_), .Y(_389_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_383_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_384_) );
OAI21X1 OAI21X1_19 ( .A(_383_), .B(_384_), .C(_17__2_), .Y(_385_) );
NAND2X1 NAND2X1_19 ( .A(_385_), .B(_389_), .Y(_0__26_) );
OAI21X1 OAI21X1_20 ( .A(_386_), .B(_383_), .C(_388_), .Y(_17__3_) );
INVX1 INVX1_10 ( .A(_17__3_), .Y(_393_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_394_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_395_) );
NAND3X1 NAND3X1_10 ( .A(_393_), .B(_395_), .C(_394_), .Y(_396_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_390_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_391_) );
OAI21X1 OAI21X1_21 ( .A(_390_), .B(_391_), .C(_17__3_), .Y(_392_) );
NAND2X1 NAND2X1_21 ( .A(_392_), .B(_396_), .Y(_0__27_) );
OAI21X1 OAI21X1_22 ( .A(_393_), .B(_390_), .C(_395_), .Y(_16_) );
INVX1 INVX1_11 ( .A(w_cout_6_), .Y(_400_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_401_) );
NAND2X1 NAND2X1_22 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_402_) );
NAND3X1 NAND3X1_11 ( .A(_400_), .B(_402_), .C(_401_), .Y(_403_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_397_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_398_) );
OAI21X1 OAI21X1_23 ( .A(_397_), .B(_398_), .C(w_cout_6_), .Y(_399_) );
NAND2X1 NAND2X1_23 ( .A(_399_), .B(_403_), .Y(_0__28_) );
OAI21X1 OAI21X1_24 ( .A(_400_), .B(_397_), .C(_402_), .Y(_20__1_) );
INVX1 INVX1_12 ( .A(_20__1_), .Y(_407_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_408_) );
NAND2X1 NAND2X1_24 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_409_) );
NAND3X1 NAND3X1_12 ( .A(_407_), .B(_409_), .C(_408_), .Y(_410_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_404_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_405_) );
OAI21X1 OAI21X1_25 ( .A(_404_), .B(_405_), .C(_20__1_), .Y(_406_) );
NAND2X1 NAND2X1_25 ( .A(_406_), .B(_410_), .Y(_0__29_) );
OAI21X1 OAI21X1_26 ( .A(_407_), .B(_404_), .C(_409_), .Y(_20__2_) );
INVX1 INVX1_13 ( .A(_20__2_), .Y(_414_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_415_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_416_) );
NAND3X1 NAND3X1_13 ( .A(_414_), .B(_416_), .C(_415_), .Y(_417_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_411_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_412_) );
OAI21X1 OAI21X1_27 ( .A(_411_), .B(_412_), .C(_20__2_), .Y(_413_) );
NAND2X1 NAND2X1_27 ( .A(_413_), .B(_417_), .Y(_0__30_) );
OAI21X1 OAI21X1_28 ( .A(_414_), .B(_411_), .C(_416_), .Y(_20__3_) );
INVX1 INVX1_14 ( .A(_20__3_), .Y(_421_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_422_) );
NAND2X1 NAND2X1_28 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_423_) );
NAND3X1 NAND3X1_14 ( .A(_421_), .B(_423_), .C(_422_), .Y(_424_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_418_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_419_) );
OAI21X1 OAI21X1_29 ( .A(_418_), .B(_419_), .C(_20__3_), .Y(_420_) );
NAND2X1 NAND2X1_29 ( .A(_420_), .B(_424_), .Y(_0__31_) );
OAI21X1 OAI21X1_30 ( .A(_421_), .B(_418_), .C(_423_), .Y(_19_) );
INVX1 INVX1_15 ( .A(w_cout_7_), .Y(_428_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_429_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_430_) );
NAND3X1 NAND3X1_15 ( .A(_428_), .B(_430_), .C(_429_), .Y(_431_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_425_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_426_) );
OAI21X1 OAI21X1_31 ( .A(_425_), .B(_426_), .C(w_cout_7_), .Y(_427_) );
NAND2X1 NAND2X1_31 ( .A(_427_), .B(_431_), .Y(_0__32_) );
OAI21X1 OAI21X1_32 ( .A(_428_), .B(_425_), .C(_430_), .Y(_23__1_) );
INVX1 INVX1_16 ( .A(_23__1_), .Y(_435_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_436_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_437_) );
NAND3X1 NAND3X1_16 ( .A(_435_), .B(_437_), .C(_436_), .Y(_438_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_432_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_433_) );
OAI21X1 OAI21X1_33 ( .A(_432_), .B(_433_), .C(_23__1_), .Y(_434_) );
NAND2X1 NAND2X1_33 ( .A(_434_), .B(_438_), .Y(_0__33_) );
OAI21X1 OAI21X1_34 ( .A(_435_), .B(_432_), .C(_437_), .Y(_23__2_) );
INVX1 INVX1_17 ( .A(_23__2_), .Y(_442_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_443_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_444_) );
NAND3X1 NAND3X1_17 ( .A(_442_), .B(_444_), .C(_443_), .Y(_445_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_439_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_440_) );
OAI21X1 OAI21X1_35 ( .A(_439_), .B(_440_), .C(_23__2_), .Y(_441_) );
NAND2X1 NAND2X1_35 ( .A(_441_), .B(_445_), .Y(_0__34_) );
OAI21X1 OAI21X1_36 ( .A(_442_), .B(_439_), .C(_444_), .Y(_23__3_) );
INVX1 INVX1_18 ( .A(_23__3_), .Y(_449_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_450_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_451_) );
NAND3X1 NAND3X1_18 ( .A(_449_), .B(_451_), .C(_450_), .Y(_452_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_446_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_447_) );
OAI21X1 OAI21X1_37 ( .A(_446_), .B(_447_), .C(_23__3_), .Y(_448_) );
NAND2X1 NAND2X1_37 ( .A(_448_), .B(_452_), .Y(_0__35_) );
OAI21X1 OAI21X1_38 ( .A(_449_), .B(_446_), .C(_451_), .Y(_22_) );
INVX1 INVX1_19 ( .A(w_cout_8_), .Y(_456_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_457_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_458_) );
NAND3X1 NAND3X1_19 ( .A(_456_), .B(_458_), .C(_457_), .Y(_459_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_453_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_454_) );
OAI21X1 OAI21X1_39 ( .A(_453_), .B(_454_), .C(w_cout_8_), .Y(_455_) );
NAND2X1 NAND2X1_39 ( .A(_455_), .B(_459_), .Y(_0__36_) );
OAI21X1 OAI21X1_40 ( .A(_456_), .B(_453_), .C(_458_), .Y(_26__1_) );
INVX1 INVX1_20 ( .A(_26__1_), .Y(_463_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_464_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_465_) );
NAND3X1 NAND3X1_20 ( .A(_463_), .B(_465_), .C(_464_), .Y(_466_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_460_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_461_) );
OAI21X1 OAI21X1_41 ( .A(_460_), .B(_461_), .C(_26__1_), .Y(_462_) );
NAND2X1 NAND2X1_41 ( .A(_462_), .B(_466_), .Y(_0__37_) );
OAI21X1 OAI21X1_42 ( .A(_463_), .B(_460_), .C(_465_), .Y(_26__2_) );
INVX1 INVX1_21 ( .A(_26__2_), .Y(_470_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_471_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_472_) );
NAND3X1 NAND3X1_21 ( .A(_470_), .B(_472_), .C(_471_), .Y(_473_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_467_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_468_) );
OAI21X1 OAI21X1_43 ( .A(_467_), .B(_468_), .C(_26__2_), .Y(_469_) );
NAND2X1 NAND2X1_43 ( .A(_469_), .B(_473_), .Y(_0__38_) );
OAI21X1 OAI21X1_44 ( .A(_470_), .B(_467_), .C(_472_), .Y(_26__3_) );
INVX1 INVX1_22 ( .A(_26__3_), .Y(_477_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_478_) );
NAND2X1 NAND2X1_44 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_479_) );
NAND3X1 NAND3X1_22 ( .A(_477_), .B(_479_), .C(_478_), .Y(_480_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_474_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_475_) );
OAI21X1 OAI21X1_45 ( .A(_474_), .B(_475_), .C(_26__3_), .Y(_476_) );
NAND2X1 NAND2X1_45 ( .A(_476_), .B(_480_), .Y(_0__39_) );
OAI21X1 OAI21X1_46 ( .A(_477_), .B(_474_), .C(_479_), .Y(_25_) );
INVX1 INVX1_23 ( .A(w_cout_9_), .Y(_484_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_485_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_486_) );
NAND3X1 NAND3X1_23 ( .A(_484_), .B(_486_), .C(_485_), .Y(_487_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_481_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_482_) );
OAI21X1 OAI21X1_47 ( .A(_481_), .B(_482_), .C(w_cout_9_), .Y(_483_) );
NAND2X1 NAND2X1_47 ( .A(_483_), .B(_487_), .Y(_0__40_) );
OAI21X1 OAI21X1_48 ( .A(_484_), .B(_481_), .C(_486_), .Y(_29__1_) );
INVX1 INVX1_24 ( .A(_29__1_), .Y(_491_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_492_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_493_) );
NAND3X1 NAND3X1_24 ( .A(_491_), .B(_493_), .C(_492_), .Y(_494_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_488_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_489_) );
OAI21X1 OAI21X1_49 ( .A(_488_), .B(_489_), .C(_29__1_), .Y(_490_) );
NAND2X1 NAND2X1_49 ( .A(_490_), .B(_494_), .Y(_0__41_) );
OAI21X1 OAI21X1_50 ( .A(_491_), .B(_488_), .C(_493_), .Y(_29__2_) );
INVX1 INVX1_25 ( .A(_29__2_), .Y(_498_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_499_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_500_) );
NAND3X1 NAND3X1_25 ( .A(_498_), .B(_500_), .C(_499_), .Y(_501_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_495_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_496_) );
OAI21X1 OAI21X1_51 ( .A(_495_), .B(_496_), .C(_29__2_), .Y(_497_) );
NAND2X1 NAND2X1_51 ( .A(_497_), .B(_501_), .Y(_0__42_) );
OAI21X1 OAI21X1_52 ( .A(_498_), .B(_495_), .C(_500_), .Y(_29__3_) );
INVX1 INVX1_26 ( .A(_29__3_), .Y(_505_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_506_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_507_) );
NAND3X1 NAND3X1_26 ( .A(_505_), .B(_507_), .C(_506_), .Y(_508_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_502_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_503_) );
OAI21X1 OAI21X1_53 ( .A(_502_), .B(_503_), .C(_29__3_), .Y(_504_) );
NAND2X1 NAND2X1_53 ( .A(_504_), .B(_508_), .Y(_0__43_) );
OAI21X1 OAI21X1_54 ( .A(_505_), .B(_502_), .C(_507_), .Y(_28_) );
INVX1 INVX1_27 ( .A(w_cout_10_), .Y(_512_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_513_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_514_) );
NAND3X1 NAND3X1_27 ( .A(_512_), .B(_514_), .C(_513_), .Y(_515_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_509_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_510_) );
OAI21X1 OAI21X1_55 ( .A(_509_), .B(_510_), .C(w_cout_10_), .Y(_511_) );
NAND2X1 NAND2X1_55 ( .A(_511_), .B(_515_), .Y(_0__44_) );
OAI21X1 OAI21X1_56 ( .A(_512_), .B(_509_), .C(_514_), .Y(_32__1_) );
INVX1 INVX1_28 ( .A(_32__1_), .Y(_519_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_520_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_521_) );
NAND3X1 NAND3X1_28 ( .A(_519_), .B(_521_), .C(_520_), .Y(_522_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_516_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_517_) );
OAI21X1 OAI21X1_57 ( .A(_516_), .B(_517_), .C(_32__1_), .Y(_518_) );
NAND2X1 NAND2X1_57 ( .A(_518_), .B(_522_), .Y(_0__45_) );
OAI21X1 OAI21X1_58 ( .A(_519_), .B(_516_), .C(_521_), .Y(_32__2_) );
INVX1 INVX1_29 ( .A(_32__2_), .Y(_526_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_527_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_528_) );
NAND3X1 NAND3X1_29 ( .A(_526_), .B(_528_), .C(_527_), .Y(_529_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_523_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_524_) );
OAI21X1 OAI21X1_59 ( .A(_523_), .B(_524_), .C(_32__2_), .Y(_525_) );
NAND2X1 NAND2X1_59 ( .A(_525_), .B(_529_), .Y(_0__46_) );
OAI21X1 OAI21X1_60 ( .A(_526_), .B(_523_), .C(_528_), .Y(_32__3_) );
INVX1 INVX1_30 ( .A(_32__3_), .Y(_533_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_534_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_535_) );
NAND3X1 NAND3X1_30 ( .A(_533_), .B(_535_), .C(_534_), .Y(_536_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_530_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_531_) );
OAI21X1 OAI21X1_61 ( .A(_530_), .B(_531_), .C(_32__3_), .Y(_532_) );
NAND2X1 NAND2X1_61 ( .A(_532_), .B(_536_), .Y(_0__47_) );
OAI21X1 OAI21X1_62 ( .A(_533_), .B(_530_), .C(_535_), .Y(_31_) );
INVX1 INVX1_31 ( .A(w_cout_11_), .Y(_540_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_541_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_542_) );
NAND3X1 NAND3X1_31 ( .A(_540_), .B(_542_), .C(_541_), .Y(_543_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_537_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_538_) );
OAI21X1 OAI21X1_63 ( .A(_537_), .B(_538_), .C(w_cout_11_), .Y(_539_) );
NAND2X1 NAND2X1_63 ( .A(_539_), .B(_543_), .Y(_0__48_) );
OAI21X1 OAI21X1_64 ( .A(_540_), .B(_537_), .C(_542_), .Y(_35__1_) );
INVX1 INVX1_32 ( .A(_35__1_), .Y(_547_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_548_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_549_) );
NAND3X1 NAND3X1_32 ( .A(_547_), .B(_549_), .C(_548_), .Y(_550_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_544_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_545_) );
OAI21X1 OAI21X1_65 ( .A(_544_), .B(_545_), .C(_35__1_), .Y(_546_) );
NAND2X1 NAND2X1_65 ( .A(_546_), .B(_550_), .Y(_0__49_) );
OAI21X1 OAI21X1_66 ( .A(_547_), .B(_544_), .C(_549_), .Y(_35__2_) );
INVX1 INVX1_33 ( .A(_35__2_), .Y(_554_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_555_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_556_) );
NAND3X1 NAND3X1_33 ( .A(_554_), .B(_556_), .C(_555_), .Y(_557_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_551_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_552_) );
OAI21X1 OAI21X1_67 ( .A(_551_), .B(_552_), .C(_35__2_), .Y(_553_) );
NAND2X1 NAND2X1_67 ( .A(_553_), .B(_557_), .Y(_0__50_) );
OAI21X1 OAI21X1_68 ( .A(_554_), .B(_551_), .C(_556_), .Y(_35__3_) );
INVX1 INVX1_34 ( .A(_35__3_), .Y(_561_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_562_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_563_) );
NAND3X1 NAND3X1_34 ( .A(_561_), .B(_563_), .C(_562_), .Y(_564_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_558_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_559_) );
OAI21X1 OAI21X1_69 ( .A(_558_), .B(_559_), .C(_35__3_), .Y(_560_) );
NAND2X1 NAND2X1_69 ( .A(_560_), .B(_564_), .Y(_0__51_) );
OAI21X1 OAI21X1_70 ( .A(_561_), .B(_558_), .C(_563_), .Y(_34_) );
INVX1 INVX1_35 ( .A(gnd), .Y(_568_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_569_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_570_) );
NAND3X1 NAND3X1_35 ( .A(_568_), .B(_570_), .C(_569_), .Y(_571_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_565_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_566_) );
OAI21X1 OAI21X1_71 ( .A(_565_), .B(_566_), .C(gnd), .Y(_567_) );
NAND2X1 NAND2X1_71 ( .A(_567_), .B(_571_), .Y(_0__0_) );
OAI21X1 OAI21X1_72 ( .A(_568_), .B(_565_), .C(_570_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_36 ( .A(rca_inst_w_CARRY_1_), .Y(_575_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_576_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_577_) );
NAND3X1 NAND3X1_36 ( .A(_575_), .B(_577_), .C(_576_), .Y(_578_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_572_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_573_) );
OAI21X1 OAI21X1_73 ( .A(_572_), .B(_573_), .C(rca_inst_w_CARRY_1_), .Y(_574_) );
NAND2X1 NAND2X1_73 ( .A(_574_), .B(_578_), .Y(_0__1_) );
OAI21X1 OAI21X1_74 ( .A(_575_), .B(_572_), .C(_577_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_37 ( .A(rca_inst_w_CARRY_2_), .Y(_582_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_583_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_584_) );
NAND3X1 NAND3X1_37 ( .A(_582_), .B(_584_), .C(_583_), .Y(_585_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_579_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_580_) );
OAI21X1 OAI21X1_75 ( .A(_579_), .B(_580_), .C(rca_inst_w_CARRY_2_), .Y(_581_) );
NAND2X1 NAND2X1_75 ( .A(_581_), .B(_585_), .Y(_0__2_) );
OAI21X1 OAI21X1_76 ( .A(_582_), .B(_579_), .C(_584_), .Y(rca_inst_w_CARRY_3_) );
INVX1 INVX1_38 ( .A(rca_inst_w_CARRY_3_), .Y(_589_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_590_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_591_) );
NAND3X1 NAND3X1_38 ( .A(_589_), .B(_591_), .C(_590_), .Y(_592_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_586_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_587_) );
OAI21X1 OAI21X1_77 ( .A(_586_), .B(_587_), .C(rca_inst_w_CARRY_3_), .Y(_588_) );
NAND2X1 NAND2X1_77 ( .A(_588_), .B(_592_), .Y(_0__3_) );
OAI21X1 OAI21X1_78 ( .A(_589_), .B(_586_), .C(_591_), .Y(cout0) );
INVX1 INVX1_39 ( .A(i_add_term1[0]), .Y(_593_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[0]), .B(_593_), .Y(_594_) );
INVX1 INVX1_40 ( .A(i_add_term2[0]), .Y(_595_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term1[0]), .B(_595_), .Y(_596_) );
INVX1 INVX1_41 ( .A(i_add_term1[1]), .Y(_597_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[1]), .B(_597_), .Y(_598_) );
INVX1 INVX1_42 ( .A(i_add_term2[1]), .Y(_599_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term1[1]), .B(_599_), .Y(_600_) );
OAI22X1 OAI22X1_1 ( .A(_594_), .B(_596_), .C(_598_), .D(_600_), .Y(_601_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_602_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_603_) );
NOR2X1 NOR2X1_44 ( .A(_602_), .B(_603_), .Y(_604_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_605_) );
NAND2X1 NAND2X1_78 ( .A(_604_), .B(_605_), .Y(_606_) );
NOR2X1 NOR2X1_45 ( .A(_601_), .B(_606_), .Y(skip0_P) );
INVX1 INVX1_43 ( .A(cout0), .Y(_607_) );
NAND2X1 NAND2X1_79 ( .A(gnd), .B(skip0_P), .Y(_608_) );
OAI21X1 OAI21X1_79 ( .A(skip0_P), .B(_607_), .C(_608_), .Y(skip0_cin_next) );
BUFX2 BUFX2_1 ( .A(w_cout_12_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
INVX1 INVX1_44 ( .A(i_add_term1[4]), .Y(_37_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[4]), .B(_37_), .Y(_38_) );
INVX1 INVX1_45 ( .A(i_add_term2[4]), .Y(_39_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term1[4]), .B(_39_), .Y(_40_) );
INVX1 INVX1_46 ( .A(i_add_term1[5]), .Y(_41_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[5]), .B(_41_), .Y(_42_) );
INVX1 INVX1_47 ( .A(i_add_term2[5]), .Y(_43_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term1[5]), .B(_43_), .Y(_44_) );
OAI22X1 OAI22X1_2 ( .A(_38_), .B(_40_), .C(_42_), .D(_44_), .Y(_45_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_46_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_47_) );
NOR2X1 NOR2X1_51 ( .A(_46_), .B(_47_), .Y(_48_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_49_) );
NAND2X1 NAND2X1_80 ( .A(_48_), .B(_49_), .Y(_50_) );
NOR2X1 NOR2X1_52 ( .A(_45_), .B(_50_), .Y(_3_) );
INVX1 INVX1_48 ( .A(_1_), .Y(_51_) );
NAND2X1 NAND2X1_81 ( .A(gnd), .B(_3_), .Y(_52_) );
OAI21X1 OAI21X1_80 ( .A(_3_), .B(_51_), .C(_52_), .Y(w_cout_1_) );
INVX1 INVX1_49 ( .A(i_add_term1[8]), .Y(_53_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[8]), .B(_53_), .Y(_54_) );
INVX1 INVX1_50 ( .A(i_add_term2[8]), .Y(_55_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term1[8]), .B(_55_), .Y(_56_) );
INVX1 INVX1_51 ( .A(i_add_term1[9]), .Y(_57_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[9]), .B(_57_), .Y(_58_) );
INVX1 INVX1_52 ( .A(i_add_term2[9]), .Y(_59_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term1[9]), .B(_59_), .Y(_60_) );
OAI22X1 OAI22X1_3 ( .A(_54_), .B(_56_), .C(_58_), .D(_60_), .Y(_61_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_62_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_63_) );
NOR2X1 NOR2X1_58 ( .A(_62_), .B(_63_), .Y(_64_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_65_) );
NAND2X1 NAND2X1_82 ( .A(_64_), .B(_65_), .Y(_66_) );
NOR2X1 NOR2X1_59 ( .A(_61_), .B(_66_), .Y(_6_) );
INVX1 INVX1_53 ( .A(_4_), .Y(_67_) );
NAND2X1 NAND2X1_83 ( .A(gnd), .B(_6_), .Y(_68_) );
OAI21X1 OAI21X1_81 ( .A(_6_), .B(_67_), .C(_68_), .Y(w_cout_2_) );
INVX1 INVX1_54 ( .A(i_add_term1[12]), .Y(_69_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[12]), .B(_69_), .Y(_70_) );
INVX1 INVX1_55 ( .A(i_add_term2[12]), .Y(_71_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term1[12]), .B(_71_), .Y(_72_) );
INVX1 INVX1_56 ( .A(i_add_term1[13]), .Y(_73_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[13]), .B(_73_), .Y(_74_) );
INVX1 INVX1_57 ( .A(i_add_term2[13]), .Y(_75_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term1[13]), .B(_75_), .Y(_76_) );
OAI22X1 OAI22X1_4 ( .A(_70_), .B(_72_), .C(_74_), .D(_76_), .Y(_77_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_78_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_79_) );
NOR2X1 NOR2X1_65 ( .A(_78_), .B(_79_), .Y(_80_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_81_) );
NAND2X1 NAND2X1_84 ( .A(_80_), .B(_81_), .Y(_82_) );
NOR2X1 NOR2X1_66 ( .A(_77_), .B(_82_), .Y(_9_) );
INVX1 INVX1_58 ( .A(_7_), .Y(_83_) );
NAND2X1 NAND2X1_85 ( .A(gnd), .B(_9_), .Y(_84_) );
OAI21X1 OAI21X1_82 ( .A(_9_), .B(_83_), .C(_84_), .Y(w_cout_3_) );
INVX1 INVX1_59 ( .A(i_add_term1[16]), .Y(_85_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[16]), .B(_85_), .Y(_86_) );
INVX1 INVX1_60 ( .A(i_add_term2[16]), .Y(_87_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term1[16]), .B(_87_), .Y(_88_) );
INVX1 INVX1_61 ( .A(i_add_term1[17]), .Y(_89_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[17]), .B(_89_), .Y(_90_) );
INVX1 INVX1_62 ( .A(i_add_term2[17]), .Y(_91_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term1[17]), .B(_91_), .Y(_92_) );
OAI22X1 OAI22X1_5 ( .A(_86_), .B(_88_), .C(_90_), .D(_92_), .Y(_93_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_94_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_95_) );
NOR2X1 NOR2X1_72 ( .A(_94_), .B(_95_), .Y(_96_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_97_) );
NAND2X1 NAND2X1_86 ( .A(_96_), .B(_97_), .Y(_98_) );
NOR2X1 NOR2X1_73 ( .A(_93_), .B(_98_), .Y(_12_) );
INVX1 INVX1_63 ( .A(_10_), .Y(_99_) );
NAND2X1 NAND2X1_87 ( .A(gnd), .B(_12_), .Y(_100_) );
OAI21X1 OAI21X1_83 ( .A(_12_), .B(_99_), .C(_100_), .Y(w_cout_4_) );
INVX1 INVX1_64 ( .A(i_add_term1[20]), .Y(_101_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[20]), .B(_101_), .Y(_102_) );
INVX1 INVX1_65 ( .A(i_add_term2[20]), .Y(_103_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term1[20]), .B(_103_), .Y(_104_) );
INVX1 INVX1_66 ( .A(i_add_term1[21]), .Y(_105_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[21]), .B(_105_), .Y(_106_) );
INVX1 INVX1_67 ( .A(i_add_term2[21]), .Y(_107_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term1[21]), .B(_107_), .Y(_108_) );
OAI22X1 OAI22X1_6 ( .A(_102_), .B(_104_), .C(_106_), .D(_108_), .Y(_109_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_110_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_111_) );
NOR2X1 NOR2X1_79 ( .A(_110_), .B(_111_), .Y(_112_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_113_) );
NAND2X1 NAND2X1_88 ( .A(_112_), .B(_113_), .Y(_114_) );
NOR2X1 NOR2X1_80 ( .A(_109_), .B(_114_), .Y(_15_) );
INVX1 INVX1_68 ( .A(_13_), .Y(_115_) );
NAND2X1 NAND2X1_89 ( .A(gnd), .B(_15_), .Y(_116_) );
OAI21X1 OAI21X1_84 ( .A(_15_), .B(_115_), .C(_116_), .Y(w_cout_5_) );
INVX1 INVX1_69 ( .A(i_add_term1[24]), .Y(_117_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[24]), .B(_117_), .Y(_118_) );
INVX1 INVX1_70 ( .A(i_add_term2[24]), .Y(_119_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term1[24]), .B(_119_), .Y(_120_) );
INVX1 INVX1_71 ( .A(i_add_term1[25]), .Y(_121_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[25]), .B(_121_), .Y(_122_) );
INVX1 INVX1_72 ( .A(i_add_term2[25]), .Y(_123_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term1[25]), .B(_123_), .Y(_124_) );
OAI22X1 OAI22X1_7 ( .A(_118_), .B(_120_), .C(_122_), .D(_124_), .Y(_125_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_126_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_127_) );
NOR2X1 NOR2X1_86 ( .A(_126_), .B(_127_), .Y(_128_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_129_) );
NAND2X1 NAND2X1_90 ( .A(_128_), .B(_129_), .Y(_130_) );
NOR2X1 NOR2X1_87 ( .A(_125_), .B(_130_), .Y(_18_) );
INVX1 INVX1_73 ( .A(_16_), .Y(_131_) );
NAND2X1 NAND2X1_91 ( .A(gnd), .B(_18_), .Y(_132_) );
OAI21X1 OAI21X1_85 ( .A(_18_), .B(_131_), .C(_132_), .Y(w_cout_6_) );
INVX1 INVX1_74 ( .A(i_add_term1[28]), .Y(_133_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[28]), .B(_133_), .Y(_134_) );
INVX1 INVX1_75 ( .A(i_add_term2[28]), .Y(_135_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term1[28]), .B(_135_), .Y(_136_) );
INVX1 INVX1_76 ( .A(i_add_term1[29]), .Y(_137_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[29]), .B(_137_), .Y(_138_) );
INVX1 INVX1_77 ( .A(i_add_term2[29]), .Y(_139_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term1[29]), .B(_139_), .Y(_140_) );
OAI22X1 OAI22X1_8 ( .A(_134_), .B(_136_), .C(_138_), .D(_140_), .Y(_141_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_142_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_143_) );
NOR2X1 NOR2X1_93 ( .A(_142_), .B(_143_), .Y(_144_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_145_) );
NAND2X1 NAND2X1_92 ( .A(_144_), .B(_145_), .Y(_146_) );
NOR2X1 NOR2X1_94 ( .A(_141_), .B(_146_), .Y(_21_) );
INVX1 INVX1_78 ( .A(_19_), .Y(_147_) );
NAND2X1 NAND2X1_93 ( .A(gnd), .B(_21_), .Y(_148_) );
OAI21X1 OAI21X1_86 ( .A(_21_), .B(_147_), .C(_148_), .Y(w_cout_7_) );
INVX1 INVX1_79 ( .A(i_add_term1[32]), .Y(_149_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[32]), .B(_149_), .Y(_150_) );
INVX1 INVX1_80 ( .A(i_add_term2[32]), .Y(_151_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term1[32]), .B(_151_), .Y(_152_) );
INVX1 INVX1_81 ( .A(i_add_term1[33]), .Y(_153_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[33]), .B(_153_), .Y(_154_) );
INVX1 INVX1_82 ( .A(i_add_term2[33]), .Y(_155_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term1[33]), .B(_155_), .Y(_156_) );
OAI22X1 OAI22X1_9 ( .A(_150_), .B(_152_), .C(_154_), .D(_156_), .Y(_157_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_158_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_159_) );
NOR2X1 NOR2X1_100 ( .A(_158_), .B(_159_), .Y(_160_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_161_) );
NAND2X1 NAND2X1_94 ( .A(_160_), .B(_161_), .Y(_162_) );
NOR2X1 NOR2X1_101 ( .A(_157_), .B(_162_), .Y(_24_) );
INVX1 INVX1_83 ( .A(_22_), .Y(_163_) );
NAND2X1 NAND2X1_95 ( .A(gnd), .B(_24_), .Y(_164_) );
OAI21X1 OAI21X1_87 ( .A(_24_), .B(_163_), .C(_164_), .Y(w_cout_8_) );
INVX1 INVX1_84 ( .A(i_add_term1[36]), .Y(_165_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[36]), .B(_165_), .Y(_166_) );
INVX1 INVX1_85 ( .A(i_add_term2[36]), .Y(_167_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term1[36]), .B(_167_), .Y(_168_) );
INVX1 INVX1_86 ( .A(i_add_term1[37]), .Y(_169_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term2[37]), .B(_169_), .Y(_170_) );
INVX1 INVX1_87 ( .A(i_add_term2[37]), .Y(_171_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term1[37]), .B(_171_), .Y(_172_) );
OAI22X1 OAI22X1_10 ( .A(_166_), .B(_168_), .C(_170_), .D(_172_), .Y(_173_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_174_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_175_) );
NOR2X1 NOR2X1_107 ( .A(_174_), .B(_175_), .Y(_176_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_177_) );
NAND2X1 NAND2X1_96 ( .A(_176_), .B(_177_), .Y(_178_) );
NOR2X1 NOR2X1_108 ( .A(_173_), .B(_178_), .Y(_27_) );
INVX1 INVX1_88 ( .A(_25_), .Y(_179_) );
NAND2X1 NAND2X1_97 ( .A(gnd), .B(_27_), .Y(_180_) );
OAI21X1 OAI21X1_88 ( .A(_27_), .B(_179_), .C(_180_), .Y(w_cout_9_) );
INVX1 INVX1_89 ( .A(i_add_term1[40]), .Y(_181_) );
NOR2X1 NOR2X1_109 ( .A(i_add_term2[40]), .B(_181_), .Y(_182_) );
INVX1 INVX1_90 ( .A(i_add_term2[40]), .Y(_183_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term1[40]), .B(_183_), .Y(_184_) );
INVX1 INVX1_91 ( .A(i_add_term1[41]), .Y(_185_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term2[41]), .B(_185_), .Y(_186_) );
INVX1 INVX1_92 ( .A(i_add_term2[41]), .Y(_187_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term1[41]), .B(_187_), .Y(_188_) );
OAI22X1 OAI22X1_11 ( .A(_182_), .B(_184_), .C(_186_), .D(_188_), .Y(_189_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_190_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_191_) );
NOR2X1 NOR2X1_114 ( .A(_190_), .B(_191_), .Y(_192_) );
XOR2X1 XOR2X1_11 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_193_) );
NAND2X1 NAND2X1_98 ( .A(_192_), .B(_193_), .Y(_194_) );
NOR2X1 NOR2X1_115 ( .A(_189_), .B(_194_), .Y(_30_) );
INVX1 INVX1_93 ( .A(_28_), .Y(_195_) );
NAND2X1 NAND2X1_99 ( .A(gnd), .B(_30_), .Y(_196_) );
OAI21X1 OAI21X1_89 ( .A(_30_), .B(_195_), .C(_196_), .Y(w_cout_10_) );
INVX1 INVX1_94 ( .A(i_add_term1[44]), .Y(_197_) );
NOR2X1 NOR2X1_116 ( .A(i_add_term2[44]), .B(_197_), .Y(_198_) );
INVX1 INVX1_95 ( .A(i_add_term2[44]), .Y(_199_) );
NOR2X1 NOR2X1_117 ( .A(i_add_term1[44]), .B(_199_), .Y(_200_) );
INVX1 INVX1_96 ( .A(i_add_term1[45]), .Y(_201_) );
NOR2X1 NOR2X1_118 ( .A(i_add_term2[45]), .B(_201_), .Y(_202_) );
INVX1 INVX1_97 ( .A(i_add_term2[45]), .Y(_203_) );
NOR2X1 NOR2X1_119 ( .A(i_add_term1[45]), .B(_203_), .Y(_204_) );
OAI22X1 OAI22X1_12 ( .A(_198_), .B(_200_), .C(_202_), .D(_204_), .Y(_205_) );
NOR2X1 NOR2X1_120 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_206_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_207_) );
NOR2X1 NOR2X1_121 ( .A(_206_), .B(_207_), .Y(_208_) );
XOR2X1 XOR2X1_12 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_209_) );
NAND2X1 NAND2X1_100 ( .A(_208_), .B(_209_), .Y(_210_) );
NOR2X1 NOR2X1_122 ( .A(_205_), .B(_210_), .Y(_33_) );
INVX1 INVX1_98 ( .A(_31_), .Y(_211_) );
NAND2X1 NAND2X1_101 ( .A(gnd), .B(_33_), .Y(_212_) );
OAI21X1 OAI21X1_90 ( .A(_33_), .B(_211_), .C(_212_), .Y(w_cout_11_) );
INVX1 INVX1_99 ( .A(i_add_term1[48]), .Y(_213_) );
NOR2X1 NOR2X1_123 ( .A(i_add_term2[48]), .B(_213_), .Y(_214_) );
INVX1 INVX1_100 ( .A(i_add_term2[48]), .Y(_215_) );
NOR2X1 NOR2X1_124 ( .A(i_add_term1[48]), .B(_215_), .Y(_216_) );
INVX1 INVX1_101 ( .A(i_add_term1[49]), .Y(_217_) );
NOR2X1 NOR2X1_125 ( .A(i_add_term2[49]), .B(_217_), .Y(_218_) );
INVX1 INVX1_102 ( .A(i_add_term2[49]), .Y(_219_) );
NOR2X1 NOR2X1_126 ( .A(i_add_term1[49]), .B(_219_), .Y(_220_) );
OAI22X1 OAI22X1_13 ( .A(_214_), .B(_216_), .C(_218_), .D(_220_), .Y(_221_) );
NOR2X1 NOR2X1_127 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_222_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_223_) );
NOR2X1 NOR2X1_128 ( .A(_222_), .B(_223_), .Y(_224_) );
XOR2X1 XOR2X1_13 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_225_) );
NAND2X1 NAND2X1_102 ( .A(_224_), .B(_225_), .Y(_226_) );
NOR2X1 NOR2X1_129 ( .A(_221_), .B(_226_), .Y(_36_) );
INVX1 INVX1_103 ( .A(_34_), .Y(_227_) );
NAND2X1 NAND2X1_103 ( .A(gnd), .B(_36_), .Y(_228_) );
OAI21X1 OAI21X1_91 ( .A(_36_), .B(_227_), .C(_228_), .Y(w_cout_12_) );
INVX1 INVX1_104 ( .A(skip0_cin_next), .Y(_232_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_233_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_234_) );
NAND3X1 NAND3X1_39 ( .A(_232_), .B(_234_), .C(_233_), .Y(_235_) );
NOR2X1 NOR2X1_130 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_229_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_230_) );
OAI21X1 OAI21X1_92 ( .A(_229_), .B(_230_), .C(skip0_cin_next), .Y(_231_) );
NAND2X1 NAND2X1_105 ( .A(_231_), .B(_235_), .Y(_0__4_) );
OAI21X1 OAI21X1_93 ( .A(_232_), .B(_229_), .C(_234_), .Y(_2__1_) );
INVX1 INVX1_105 ( .A(_2__1_), .Y(_239_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_240_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_241_) );
NAND3X1 NAND3X1_40 ( .A(_239_), .B(_241_), .C(_240_), .Y(_242_) );
NOR2X1 NOR2X1_131 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_236_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_237_) );
OAI21X1 OAI21X1_94 ( .A(_236_), .B(_237_), .C(_2__1_), .Y(_238_) );
NAND2X1 NAND2X1_107 ( .A(_238_), .B(_242_), .Y(_0__5_) );
OAI21X1 OAI21X1_95 ( .A(_239_), .B(_236_), .C(_241_), .Y(_2__2_) );
INVX1 INVX1_106 ( .A(_2__2_), .Y(_246_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_247_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_248_) );
NAND3X1 NAND3X1_41 ( .A(_246_), .B(_248_), .C(_247_), .Y(_249_) );
NOR2X1 NOR2X1_132 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_243_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_244_) );
OAI21X1 OAI21X1_96 ( .A(_243_), .B(_244_), .C(_2__2_), .Y(_245_) );
NAND2X1 NAND2X1_109 ( .A(_245_), .B(_249_), .Y(_0__6_) );
OAI21X1 OAI21X1_97 ( .A(_246_), .B(_243_), .C(_248_), .Y(_2__3_) );
INVX1 INVX1_107 ( .A(_2__3_), .Y(_253_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_254_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_255_) );
NAND3X1 NAND3X1_42 ( .A(_253_), .B(_255_), .C(_254_), .Y(_256_) );
NOR2X1 NOR2X1_133 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_250_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_251_) );
OAI21X1 OAI21X1_98 ( .A(_250_), .B(_251_), .C(_2__3_), .Y(_252_) );
NAND2X1 NAND2X1_111 ( .A(_252_), .B(_256_), .Y(_0__7_) );
OAI21X1 OAI21X1_99 ( .A(_253_), .B(_250_), .C(_255_), .Y(_1_) );
INVX1 INVX1_108 ( .A(w_cout_1_), .Y(_260_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_261_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_262_) );
NAND3X1 NAND3X1_43 ( .A(_260_), .B(_262_), .C(_261_), .Y(_263_) );
NOR2X1 NOR2X1_134 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_257_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_258_) );
OAI21X1 OAI21X1_100 ( .A(_257_), .B(_258_), .C(w_cout_1_), .Y(_259_) );
NAND2X1 NAND2X1_113 ( .A(_259_), .B(_263_), .Y(_0__8_) );
OAI21X1 OAI21X1_101 ( .A(_260_), .B(_257_), .C(_262_), .Y(_5__1_) );
INVX1 INVX1_109 ( .A(_5__1_), .Y(_267_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_268_) );
NAND2X1 NAND2X1_114 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_269_) );
NAND3X1 NAND3X1_44 ( .A(_267_), .B(_269_), .C(_268_), .Y(_270_) );
NOR2X1 NOR2X1_135 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_264_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_265_) );
OAI21X1 OAI21X1_102 ( .A(_264_), .B(_265_), .C(_5__1_), .Y(_266_) );
NAND2X1 NAND2X1_115 ( .A(_266_), .B(_270_), .Y(_0__9_) );
OAI21X1 OAI21X1_103 ( .A(_267_), .B(_264_), .C(_269_), .Y(_5__2_) );
INVX1 INVX1_110 ( .A(_5__2_), .Y(_274_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_275_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_276_) );
NAND3X1 NAND3X1_45 ( .A(_274_), .B(_276_), .C(_275_), .Y(_277_) );
NOR2X1 NOR2X1_136 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_271_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_272_) );
OAI21X1 OAI21X1_104 ( .A(_271_), .B(_272_), .C(_5__2_), .Y(_273_) );
NAND2X1 NAND2X1_117 ( .A(_273_), .B(_277_), .Y(_0__10_) );
OAI21X1 OAI21X1_105 ( .A(_274_), .B(_271_), .C(_276_), .Y(_5__3_) );
INVX1 INVX1_111 ( .A(_5__3_), .Y(_281_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_282_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_283_) );
NAND3X1 NAND3X1_46 ( .A(_281_), .B(_283_), .C(_282_), .Y(_284_) );
NOR2X1 NOR2X1_137 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_278_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_279_) );
OAI21X1 OAI21X1_106 ( .A(_278_), .B(_279_), .C(_5__3_), .Y(_280_) );
NAND2X1 NAND2X1_119 ( .A(_280_), .B(_284_), .Y(_0__11_) );
OAI21X1 OAI21X1_107 ( .A(_281_), .B(_278_), .C(_283_), .Y(_4_) );
INVX1 INVX1_112 ( .A(w_cout_2_), .Y(_288_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_289_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_290_) );
NAND3X1 NAND3X1_47 ( .A(_288_), .B(_290_), .C(_289_), .Y(_291_) );
NOR2X1 NOR2X1_138 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_285_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_286_) );
OAI21X1 OAI21X1_108 ( .A(_285_), .B(_286_), .C(w_cout_2_), .Y(_287_) );
NAND2X1 NAND2X1_121 ( .A(_287_), .B(_291_), .Y(_0__12_) );
OAI21X1 OAI21X1_109 ( .A(_288_), .B(_285_), .C(_290_), .Y(_8__1_) );
INVX1 INVX1_113 ( .A(_8__1_), .Y(_295_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_296_) );
NAND2X1 NAND2X1_122 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_297_) );
NAND3X1 NAND3X1_48 ( .A(_295_), .B(_297_), .C(_296_), .Y(_298_) );
NOR2X1 NOR2X1_139 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_292_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_293_) );
OAI21X1 OAI21X1_110 ( .A(_292_), .B(_293_), .C(_8__1_), .Y(_294_) );
NAND2X1 NAND2X1_123 ( .A(_294_), .B(_298_), .Y(_0__13_) );
OAI21X1 OAI21X1_111 ( .A(_295_), .B(_292_), .C(_297_), .Y(_8__2_) );
INVX1 INVX1_114 ( .A(_8__2_), .Y(_302_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_303_) );
NAND2X1 NAND2X1_124 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_304_) );
NAND3X1 NAND3X1_49 ( .A(_302_), .B(_304_), .C(_303_), .Y(_305_) );
NOR2X1 NOR2X1_140 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_299_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_300_) );
OAI21X1 OAI21X1_112 ( .A(_299_), .B(_300_), .C(_8__2_), .Y(_301_) );
NAND2X1 NAND2X1_125 ( .A(_301_), .B(_305_), .Y(_0__14_) );
OAI21X1 OAI21X1_113 ( .A(_302_), .B(_299_), .C(_304_), .Y(_8__3_) );
INVX1 INVX1_115 ( .A(_8__3_), .Y(_309_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_310_) );
NAND2X1 NAND2X1_126 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_311_) );
NAND3X1 NAND3X1_50 ( .A(_309_), .B(_311_), .C(_310_), .Y(_312_) );
NOR2X1 NOR2X1_141 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_306_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_307_) );
OAI21X1 OAI21X1_114 ( .A(_306_), .B(_307_), .C(_8__3_), .Y(_308_) );
NAND2X1 NAND2X1_127 ( .A(_308_), .B(_312_), .Y(_0__15_) );
OAI21X1 OAI21X1_115 ( .A(_309_), .B(_306_), .C(_311_), .Y(_7_) );
INVX1 INVX1_116 ( .A(w_cout_3_), .Y(_316_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_317_) );
NAND2X1 NAND2X1_128 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_318_) );
NAND3X1 NAND3X1_51 ( .A(_316_), .B(_318_), .C(_317_), .Y(_319_) );
NOR2X1 NOR2X1_142 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_313_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_314_) );
OAI21X1 OAI21X1_116 ( .A(_313_), .B(_314_), .C(w_cout_3_), .Y(_315_) );
NAND2X1 NAND2X1_129 ( .A(_315_), .B(_319_), .Y(_0__16_) );
OAI21X1 OAI21X1_117 ( .A(_316_), .B(_313_), .C(_318_), .Y(_11__1_) );
INVX1 INVX1_117 ( .A(_11__1_), .Y(_323_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_324_) );
NAND2X1 NAND2X1_130 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_325_) );
NAND3X1 NAND3X1_52 ( .A(_323_), .B(_325_), .C(_324_), .Y(_326_) );
NOR2X1 NOR2X1_143 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_320_) );
BUFX2 BUFX2_54 ( .A(skip0_cin_next), .Y(_2__0_) );
BUFX2 BUFX2_55 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_56 ( .A(w_cout_1_), .Y(_5__0_) );
BUFX2 BUFX2_57 ( .A(_4_), .Y(_5__4_) );
BUFX2 BUFX2_58 ( .A(w_cout_2_), .Y(_8__0_) );
BUFX2 BUFX2_59 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_60 ( .A(w_cout_3_), .Y(_11__0_) );
BUFX2 BUFX2_61 ( .A(_10_), .Y(_11__4_) );
BUFX2 BUFX2_62 ( .A(w_cout_4_), .Y(_14__0_) );
BUFX2 BUFX2_63 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_64 ( .A(w_cout_5_), .Y(_17__0_) );
BUFX2 BUFX2_65 ( .A(_16_), .Y(_17__4_) );
BUFX2 BUFX2_66 ( .A(w_cout_6_), .Y(_20__0_) );
BUFX2 BUFX2_67 ( .A(_19_), .Y(_20__4_) );
BUFX2 BUFX2_68 ( .A(w_cout_7_), .Y(_23__0_) );
BUFX2 BUFX2_69 ( .A(_22_), .Y(_23__4_) );
BUFX2 BUFX2_70 ( .A(w_cout_8_), .Y(_26__0_) );
BUFX2 BUFX2_71 ( .A(_25_), .Y(_26__4_) );
BUFX2 BUFX2_72 ( .A(w_cout_9_), .Y(_29__0_) );
BUFX2 BUFX2_73 ( .A(_28_), .Y(_29__4_) );
BUFX2 BUFX2_74 ( .A(w_cout_10_), .Y(_32__0_) );
BUFX2 BUFX2_75 ( .A(_31_), .Y(_32__4_) );
BUFX2 BUFX2_76 ( .A(w_cout_11_), .Y(_35__0_) );
BUFX2 BUFX2_77 ( .A(_34_), .Y(_35__4_) );
BUFX2 BUFX2_78 ( .A(gnd), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_79 ( .A(cout0), .Y(rca_inst_w_CARRY_4_) );
BUFX2 BUFX2_80 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
