module csa_15bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_3_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_19_) );
NAND2X1 NAND2X1_1 ( .A(_2_), .B(1'b0), .Y(_20_) );
OAI21X1 OAI21X1_1 ( .A(1'b0), .B(_19_), .C(_20_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3__3_), .Y(_21_) );
NAND2X1 NAND2X1_2 ( .A(_4__3_), .B(1'b0), .Y(_22_) );
OAI21X1 OAI21X1_2 ( .A(1'b0), .B(_21_), .C(_22_), .Y(_0__6_) );
INVX1 INVX1_3 ( .A(_3__0_), .Y(_23_) );
NAND2X1 NAND2X1_3 ( .A(1'b0), .B(_4__0_), .Y(_24_) );
OAI21X1 OAI21X1_3 ( .A(1'b0), .B(_23_), .C(_24_), .Y(_0__3_) );
INVX1 INVX1_4 ( .A(_3__1_), .Y(_25_) );
NAND2X1 NAND2X1_4 ( .A(1'b0), .B(_4__1_), .Y(_26_) );
OAI21X1 OAI21X1_4 ( .A(1'b0), .B(_25_), .C(_26_), .Y(_0__4_) );
INVX1 INVX1_5 ( .A(_3__2_), .Y(_27_) );
NAND2X1 NAND2X1_5 ( .A(1'b0), .B(_4__2_), .Y(_28_) );
OAI21X1 OAI21X1_5 ( .A(1'b0), .B(_27_), .C(_28_), .Y(_0__5_) );
INVX1 INVX1_6 ( .A(_7_), .Y(_29_) );
NAND2X1 NAND2X1_6 ( .A(_8_), .B(w_cout_1_), .Y(_30_) );
OAI21X1 OAI21X1_6 ( .A(w_cout_1_), .B(_29_), .C(_30_), .Y(w_cout_2_) );
INVX1 INVX1_7 ( .A(_9__3_), .Y(_31_) );
NAND2X1 NAND2X1_7 ( .A(_10__3_), .B(w_cout_1_), .Y(_32_) );
OAI21X1 OAI21X1_7 ( .A(w_cout_1_), .B(_31_), .C(_32_), .Y(_0__10_) );
INVX1 INVX1_8 ( .A(_9__0_), .Y(_33_) );
NAND2X1 NAND2X1_8 ( .A(w_cout_1_), .B(_10__0_), .Y(_34_) );
OAI21X1 OAI21X1_8 ( .A(w_cout_1_), .B(_33_), .C(_34_), .Y(_0__7_) );
INVX1 INVX1_9 ( .A(_9__1_), .Y(_35_) );
NAND2X1 NAND2X1_9 ( .A(w_cout_1_), .B(_10__1_), .Y(_36_) );
OAI21X1 OAI21X1_9 ( .A(w_cout_1_), .B(_35_), .C(_36_), .Y(_0__8_) );
INVX1 INVX1_10 ( .A(_9__2_), .Y(_37_) );
NAND2X1 NAND2X1_10 ( .A(w_cout_1_), .B(_10__2_), .Y(_38_) );
OAI21X1 OAI21X1_10 ( .A(w_cout_1_), .B(_37_), .C(_38_), .Y(_0__9_) );
INVX1 INVX1_11 ( .A(_13_), .Y(_39_) );
NAND2X1 NAND2X1_11 ( .A(_14_), .B(w_cout_2_), .Y(_40_) );
OAI21X1 OAI21X1_11 ( .A(w_cout_2_), .B(_39_), .C(_40_), .Y(w_cout_3_) );
INVX1 INVX1_12 ( .A(_15__3_), .Y(_41_) );
NAND2X1 NAND2X1_12 ( .A(_16__3_), .B(w_cout_2_), .Y(_42_) );
OAI21X1 OAI21X1_12 ( .A(w_cout_2_), .B(_41_), .C(_42_), .Y(_0__14_) );
INVX1 INVX1_13 ( .A(_15__0_), .Y(_43_) );
NAND2X1 NAND2X1_13 ( .A(w_cout_2_), .B(_16__0_), .Y(_44_) );
OAI21X1 OAI21X1_13 ( .A(w_cout_2_), .B(_43_), .C(_44_), .Y(_0__11_) );
INVX1 INVX1_14 ( .A(_15__1_), .Y(_45_) );
NAND2X1 NAND2X1_14 ( .A(w_cout_2_), .B(_16__1_), .Y(_46_) );
OAI21X1 OAI21X1_14 ( .A(w_cout_2_), .B(_45_), .C(_46_), .Y(_0__12_) );
INVX1 INVX1_15 ( .A(_15__2_), .Y(_47_) );
NAND2X1 NAND2X1_15 ( .A(w_cout_2_), .B(_16__2_), .Y(_48_) );
OAI21X1 OAI21X1_15 ( .A(w_cout_2_), .B(_47_), .C(_48_), .Y(_0__13_) );
INVX1 INVX1_16 ( .A(1'b0), .Y(_52_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_53_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_54_) );
NAND3X1 NAND3X1_1 ( .A(_52_), .B(_54_), .C(_53_), .Y(_55_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_49_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_50_) );
OAI21X1 OAI21X1_16 ( .A(_49_), .B(_50_), .C(1'b0), .Y(_51_) );
NAND2X1 NAND2X1_17 ( .A(_51_), .B(_55_), .Y(_3__0_) );
OAI21X1 OAI21X1_17 ( .A(_52_), .B(_49_), .C(_54_), .Y(_5__1_) );
INVX1 INVX1_17 ( .A(_5__1_), .Y(_59_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_60_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_61_) );
NAND3X1 NAND3X1_2 ( .A(_59_), .B(_61_), .C(_60_), .Y(_62_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_56_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_57_) );
OAI21X1 OAI21X1_18 ( .A(_56_), .B(_57_), .C(_5__1_), .Y(_58_) );
NAND2X1 NAND2X1_19 ( .A(_58_), .B(_62_), .Y(_3__1_) );
OAI21X1 OAI21X1_19 ( .A(_59_), .B(_56_), .C(_61_), .Y(_5__2_) );
INVX1 INVX1_18 ( .A(_5__2_), .Y(_66_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_67_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_68_) );
NAND3X1 NAND3X1_3 ( .A(_66_), .B(_68_), .C(_67_), .Y(_69_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_63_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_64_) );
OAI21X1 OAI21X1_20 ( .A(_63_), .B(_64_), .C(_5__2_), .Y(_65_) );
NAND2X1 NAND2X1_21 ( .A(_65_), .B(_69_), .Y(_3__2_) );
OAI21X1 OAI21X1_21 ( .A(_66_), .B(_63_), .C(_68_), .Y(_5__3_) );
INVX1 INVX1_19 ( .A(_5__3_), .Y(_73_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_74_) );
NAND2X1 NAND2X1_22 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_75_) );
NAND3X1 NAND3X1_4 ( .A(_73_), .B(_75_), .C(_74_), .Y(_76_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_70_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_71_) );
OAI21X1 OAI21X1_22 ( .A(_70_), .B(_71_), .C(_5__3_), .Y(_72_) );
NAND2X1 NAND2X1_23 ( .A(_72_), .B(_76_), .Y(_3__3_) );
OAI21X1 OAI21X1_23 ( .A(_73_), .B(_70_), .C(_75_), .Y(_1_) );
INVX1 INVX1_20 ( .A(1'b1), .Y(_80_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_81_) );
NAND2X1 NAND2X1_24 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_82_) );
NAND3X1 NAND3X1_5 ( .A(_80_), .B(_82_), .C(_81_), .Y(_83_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_77_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_78_) );
OAI21X1 OAI21X1_24 ( .A(_77_), .B(_78_), .C(1'b1), .Y(_79_) );
NAND2X1 NAND2X1_25 ( .A(_79_), .B(_83_), .Y(_4__0_) );
OAI21X1 OAI21X1_25 ( .A(_80_), .B(_77_), .C(_82_), .Y(_6__1_) );
INVX1 INVX1_21 ( .A(_6__1_), .Y(_87_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_88_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_89_) );
NAND3X1 NAND3X1_6 ( .A(_87_), .B(_89_), .C(_88_), .Y(_90_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_84_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_85_) );
OAI21X1 OAI21X1_26 ( .A(_84_), .B(_85_), .C(_6__1_), .Y(_86_) );
NAND2X1 NAND2X1_27 ( .A(_86_), .B(_90_), .Y(_4__1_) );
OAI21X1 OAI21X1_27 ( .A(_87_), .B(_84_), .C(_89_), .Y(_6__2_) );
INVX1 INVX1_22 ( .A(_6__2_), .Y(_94_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_95_) );
NAND2X1 NAND2X1_28 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_96_) );
NAND3X1 NAND3X1_7 ( .A(_94_), .B(_96_), .C(_95_), .Y(_97_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_91_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_92_) );
OAI21X1 OAI21X1_28 ( .A(_91_), .B(_92_), .C(_6__2_), .Y(_93_) );
NAND2X1 NAND2X1_29 ( .A(_93_), .B(_97_), .Y(_4__2_) );
OAI21X1 OAI21X1_29 ( .A(_94_), .B(_91_), .C(_96_), .Y(_6__3_) );
INVX1 INVX1_23 ( .A(_6__3_), .Y(_101_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_102_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_103_) );
NAND3X1 NAND3X1_8 ( .A(_101_), .B(_103_), .C(_102_), .Y(_104_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_98_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_99_) );
OAI21X1 OAI21X1_30 ( .A(_98_), .B(_99_), .C(_6__3_), .Y(_100_) );
NAND2X1 NAND2X1_31 ( .A(_100_), .B(_104_), .Y(_4__3_) );
OAI21X1 OAI21X1_31 ( .A(_101_), .B(_98_), .C(_103_), .Y(_2_) );
INVX1 INVX1_24 ( .A(1'b0), .Y(_108_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_109_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_110_) );
NAND3X1 NAND3X1_9 ( .A(_108_), .B(_110_), .C(_109_), .Y(_111_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_105_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_106_) );
OAI21X1 OAI21X1_32 ( .A(_105_), .B(_106_), .C(1'b0), .Y(_107_) );
NAND2X1 NAND2X1_33 ( .A(_107_), .B(_111_), .Y(_9__0_) );
OAI21X1 OAI21X1_33 ( .A(_108_), .B(_105_), .C(_110_), .Y(_11__1_) );
INVX1 INVX1_25 ( .A(_11__1_), .Y(_115_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_116_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_117_) );
NAND3X1 NAND3X1_10 ( .A(_115_), .B(_117_), .C(_116_), .Y(_118_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_112_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_113_) );
OAI21X1 OAI21X1_34 ( .A(_112_), .B(_113_), .C(_11__1_), .Y(_114_) );
NAND2X1 NAND2X1_35 ( .A(_114_), .B(_118_), .Y(_9__1_) );
OAI21X1 OAI21X1_35 ( .A(_115_), .B(_112_), .C(_117_), .Y(_11__2_) );
INVX1 INVX1_26 ( .A(_11__2_), .Y(_122_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_123_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_124_) );
NAND3X1 NAND3X1_11 ( .A(_122_), .B(_124_), .C(_123_), .Y(_125_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_119_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_120_) );
OAI21X1 OAI21X1_36 ( .A(_119_), .B(_120_), .C(_11__2_), .Y(_121_) );
NAND2X1 NAND2X1_37 ( .A(_121_), .B(_125_), .Y(_9__2_) );
OAI21X1 OAI21X1_37 ( .A(_122_), .B(_119_), .C(_124_), .Y(_11__3_) );
INVX1 INVX1_27 ( .A(_11__3_), .Y(_129_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_130_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_131_) );
NAND3X1 NAND3X1_12 ( .A(_129_), .B(_131_), .C(_130_), .Y(_132_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_126_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_127_) );
OAI21X1 OAI21X1_38 ( .A(_126_), .B(_127_), .C(_11__3_), .Y(_128_) );
NAND2X1 NAND2X1_39 ( .A(_128_), .B(_132_), .Y(_9__3_) );
OAI21X1 OAI21X1_39 ( .A(_129_), .B(_126_), .C(_131_), .Y(_7_) );
INVX1 INVX1_28 ( .A(1'b1), .Y(_136_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_137_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_138_) );
NAND3X1 NAND3X1_13 ( .A(_136_), .B(_138_), .C(_137_), .Y(_139_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_133_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_134_) );
OAI21X1 OAI21X1_40 ( .A(_133_), .B(_134_), .C(1'b1), .Y(_135_) );
NAND2X1 NAND2X1_41 ( .A(_135_), .B(_139_), .Y(_10__0_) );
OAI21X1 OAI21X1_41 ( .A(_136_), .B(_133_), .C(_138_), .Y(_12__1_) );
INVX1 INVX1_29 ( .A(_12__1_), .Y(_143_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_144_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_145_) );
NAND3X1 NAND3X1_14 ( .A(_143_), .B(_145_), .C(_144_), .Y(_146_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_140_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_141_) );
OAI21X1 OAI21X1_42 ( .A(_140_), .B(_141_), .C(_12__1_), .Y(_142_) );
NAND2X1 NAND2X1_43 ( .A(_142_), .B(_146_), .Y(_10__1_) );
OAI21X1 OAI21X1_43 ( .A(_143_), .B(_140_), .C(_145_), .Y(_12__2_) );
INVX1 INVX1_30 ( .A(_12__2_), .Y(_150_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_151_) );
NAND2X1 NAND2X1_44 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_152_) );
NAND3X1 NAND3X1_15 ( .A(_150_), .B(_152_), .C(_151_), .Y(_153_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_147_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_148_) );
OAI21X1 OAI21X1_44 ( .A(_147_), .B(_148_), .C(_12__2_), .Y(_149_) );
NAND2X1 NAND2X1_45 ( .A(_149_), .B(_153_), .Y(_10__2_) );
OAI21X1 OAI21X1_45 ( .A(_150_), .B(_147_), .C(_152_), .Y(_12__3_) );
INVX1 INVX1_31 ( .A(_12__3_), .Y(_157_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_158_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_159_) );
NAND3X1 NAND3X1_16 ( .A(_157_), .B(_159_), .C(_158_), .Y(_160_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_154_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_155_) );
OAI21X1 OAI21X1_46 ( .A(_154_), .B(_155_), .C(_12__3_), .Y(_156_) );
NAND2X1 NAND2X1_47 ( .A(_156_), .B(_160_), .Y(_10__3_) );
OAI21X1 OAI21X1_47 ( .A(_157_), .B(_154_), .C(_159_), .Y(_8_) );
INVX1 INVX1_32 ( .A(1'b0), .Y(_164_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_165_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_166_) );
NAND3X1 NAND3X1_17 ( .A(_164_), .B(_166_), .C(_165_), .Y(_167_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_161_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_162_) );
OAI21X1 OAI21X1_48 ( .A(_161_), .B(_162_), .C(1'b0), .Y(_163_) );
NAND2X1 NAND2X1_49 ( .A(_163_), .B(_167_), .Y(_15__0_) );
OAI21X1 OAI21X1_49 ( .A(_164_), .B(_161_), .C(_166_), .Y(_17__1_) );
INVX1 INVX1_33 ( .A(_17__1_), .Y(_171_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_172_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_173_) );
NAND3X1 NAND3X1_18 ( .A(_171_), .B(_173_), .C(_172_), .Y(_174_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_168_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_169_) );
OAI21X1 OAI21X1_50 ( .A(_168_), .B(_169_), .C(_17__1_), .Y(_170_) );
NAND2X1 NAND2X1_51 ( .A(_170_), .B(_174_), .Y(_15__1_) );
OAI21X1 OAI21X1_51 ( .A(_171_), .B(_168_), .C(_173_), .Y(_17__2_) );
INVX1 INVX1_34 ( .A(_17__2_), .Y(_178_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_179_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_180_) );
NAND3X1 NAND3X1_19 ( .A(_178_), .B(_180_), .C(_179_), .Y(_181_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_175_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_176_) );
OAI21X1 OAI21X1_52 ( .A(_175_), .B(_176_), .C(_17__2_), .Y(_177_) );
NAND2X1 NAND2X1_53 ( .A(_177_), .B(_181_), .Y(_15__2_) );
OAI21X1 OAI21X1_53 ( .A(_178_), .B(_175_), .C(_180_), .Y(_17__3_) );
INVX1 INVX1_35 ( .A(_17__3_), .Y(_185_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_186_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_187_) );
NAND3X1 NAND3X1_20 ( .A(_185_), .B(_187_), .C(_186_), .Y(_188_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_182_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_183_) );
OAI21X1 OAI21X1_54 ( .A(_182_), .B(_183_), .C(_17__3_), .Y(_184_) );
NAND2X1 NAND2X1_55 ( .A(_184_), .B(_188_), .Y(_15__3_) );
OAI21X1 OAI21X1_55 ( .A(_185_), .B(_182_), .C(_187_), .Y(_13_) );
INVX1 INVX1_36 ( .A(1'b1), .Y(_192_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_193_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_194_) );
NAND3X1 NAND3X1_21 ( .A(_192_), .B(_194_), .C(_193_), .Y(_195_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_189_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_190_) );
OAI21X1 OAI21X1_56 ( .A(_189_), .B(_190_), .C(1'b1), .Y(_191_) );
NAND2X1 NAND2X1_57 ( .A(_191_), .B(_195_), .Y(_16__0_) );
OAI21X1 OAI21X1_57 ( .A(_192_), .B(_189_), .C(_194_), .Y(_18__1_) );
INVX1 INVX1_37 ( .A(_18__1_), .Y(_199_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_200_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_201_) );
NAND3X1 NAND3X1_22 ( .A(_199_), .B(_201_), .C(_200_), .Y(_202_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_196_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_197_) );
OAI21X1 OAI21X1_58 ( .A(_196_), .B(_197_), .C(_18__1_), .Y(_198_) );
NAND2X1 NAND2X1_59 ( .A(_198_), .B(_202_), .Y(_16__1_) );
OAI21X1 OAI21X1_59 ( .A(_199_), .B(_196_), .C(_201_), .Y(_18__2_) );
INVX1 INVX1_38 ( .A(_18__2_), .Y(_206_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_207_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_208_) );
NAND3X1 NAND3X1_23 ( .A(_206_), .B(_208_), .C(_207_), .Y(_209_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_203_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_204_) );
OAI21X1 OAI21X1_60 ( .A(_203_), .B(_204_), .C(_18__2_), .Y(_205_) );
NAND2X1 NAND2X1_61 ( .A(_205_), .B(_209_), .Y(_16__2_) );
OAI21X1 OAI21X1_61 ( .A(_206_), .B(_203_), .C(_208_), .Y(_18__3_) );
INVX1 INVX1_39 ( .A(_18__3_), .Y(_213_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_214_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_215_) );
NAND3X1 NAND3X1_24 ( .A(_213_), .B(_215_), .C(_214_), .Y(_216_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_210_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_211_) );
OAI21X1 OAI21X1_62 ( .A(_210_), .B(_211_), .C(_18__3_), .Y(_212_) );
NAND2X1 NAND2X1_63 ( .A(_212_), .B(_216_), .Y(_16__3_) );
OAI21X1 OAI21X1_63 ( .A(_213_), .B(_210_), .C(_215_), .Y(_14_) );
INVX1 INVX1_40 ( .A(1'b0), .Y(_220_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_221_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_222_) );
NAND3X1 NAND3X1_25 ( .A(_220_), .B(_222_), .C(_221_), .Y(_223_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_217_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_218_) );
OAI21X1 OAI21X1_64 ( .A(_217_), .B(_218_), .C(1'b0), .Y(_219_) );
NAND2X1 NAND2X1_65 ( .A(_219_), .B(_223_), .Y(_0__0_) );
OAI21X1 OAI21X1_65 ( .A(_220_), .B(_217_), .C(_222_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_41 ( .A(rca_inst_w_CARRY_1_), .Y(_227_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_228_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_229_) );
NAND3X1 NAND3X1_26 ( .A(_227_), .B(_229_), .C(_228_), .Y(_230_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_224_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_225_) );
OAI21X1 OAI21X1_66 ( .A(_224_), .B(_225_), .C(rca_inst_w_CARRY_1_), .Y(_226_) );
NAND2X1 NAND2X1_67 ( .A(_226_), .B(_230_), .Y(_0__1_) );
OAI21X1 OAI21X1_67 ( .A(_227_), .B(_224_), .C(_229_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_42 ( .A(rca_inst_w_CARRY_2_), .Y(_234_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_235_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_236_) );
NAND3X1 NAND3X1_27 ( .A(_234_), .B(_236_), .C(_235_), .Y(_237_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_231_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_232_) );
OAI21X1 OAI21X1_68 ( .A(_231_), .B(_232_), .C(rca_inst_w_CARRY_2_), .Y(_233_) );
NAND2X1 NAND2X1_69 ( .A(_233_), .B(_237_), .Y(_0__2_) );
BUFX2 BUFX2_17 ( .A(1'b0), .Y(_5__0_) );
BUFX2 BUFX2_18 ( .A(_1_), .Y(_5__4_) );
BUFX2 BUFX2_19 ( .A(1'b1), .Y(_6__0_) );
BUFX2 BUFX2_20 ( .A(_2_), .Y(_6__4_) );
BUFX2 BUFX2_21 ( .A(1'b0), .Y(_11__0_) );
BUFX2 BUFX2_22 ( .A(_7_), .Y(_11__4_) );
BUFX2 BUFX2_23 ( .A(1'b1), .Y(_12__0_) );
BUFX2 BUFX2_24 ( .A(_8_), .Y(_12__4_) );
BUFX2 BUFX2_25 ( .A(1'b0), .Y(_17__0_) );
BUFX2 BUFX2_26 ( .A(_13_), .Y(_17__4_) );
BUFX2 BUFX2_27 ( .A(1'b1), .Y(_18__0_) );
BUFX2 BUFX2_28 ( .A(_14_), .Y(_18__4_) );
BUFX2 BUFX2_29 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_30 ( .A(1'b0), .Y(w_cout_0_) );
endmodule
