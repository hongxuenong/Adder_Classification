module CSkipA_19bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_5_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(cskip3_inst_rca0_fa0_o_sum), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(cskip3_inst_rca0_fa1_o_sum), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(cskip3_inst_rca0_fa2_o_sum), .Y(sum[18]) );
INVX1 INVX1_1 ( .A(1'b0), .Y(_16_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_17_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_18_) );
NAND3X1 NAND3X1_1 ( .A(_16_), .B(_18_), .C(_17_), .Y(_19_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_13_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_14_) );
OAI21X1 OAI21X1_1 ( .A(_13_), .B(_14_), .C(1'b0), .Y(_15_) );
NAND2X1 NAND2X1_2 ( .A(_15_), .B(_19_), .Y(_0__0_) );
OAI21X1 OAI21X1_2 ( .A(_16_), .B(_13_), .C(_18_), .Y(_2__1_) );
INVX1 INVX1_2 ( .A(_2__3_), .Y(_23_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_24_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_25_) );
NAND3X1 NAND3X1_2 ( .A(_23_), .B(_25_), .C(_24_), .Y(_26_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_20_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_21_) );
OAI21X1 OAI21X1_3 ( .A(_20_), .B(_21_), .C(_2__3_), .Y(_22_) );
NAND2X1 NAND2X1_4 ( .A(_22_), .B(_26_), .Y(_0__3_) );
OAI21X1 OAI21X1_4 ( .A(_23_), .B(_20_), .C(_25_), .Y(_1_) );
INVX1 INVX1_3 ( .A(_2__1_), .Y(_30_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_31_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_32_) );
NAND3X1 NAND3X1_3 ( .A(_30_), .B(_32_), .C(_31_), .Y(_33_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_27_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_28_) );
OAI21X1 OAI21X1_5 ( .A(_27_), .B(_28_), .C(_2__1_), .Y(_29_) );
NAND2X1 NAND2X1_6 ( .A(_29_), .B(_33_), .Y(_0__1_) );
OAI21X1 OAI21X1_6 ( .A(_30_), .B(_27_), .C(_32_), .Y(_2__2_) );
INVX1 INVX1_4 ( .A(_2__2_), .Y(_37_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_38_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_39_) );
NAND3X1 NAND3X1_4 ( .A(_37_), .B(_39_), .C(_38_), .Y(_40_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_34_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_35_) );
OAI21X1 OAI21X1_7 ( .A(_34_), .B(_35_), .C(_2__2_), .Y(_36_) );
NAND2X1 NAND2X1_8 ( .A(_36_), .B(_40_), .Y(_0__2_) );
OAI21X1 OAI21X1_8 ( .A(_37_), .B(_34_), .C(_39_), .Y(_2__3_) );
INVX1 INVX1_5 ( .A(i_add_term1[0]), .Y(_41_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[0]), .B(_41_), .Y(_42_) );
INVX1 INVX1_6 ( .A(i_add_term2[0]), .Y(_43_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term1[0]), .B(_43_), .Y(_44_) );
INVX1 INVX1_7 ( .A(i_add_term1[1]), .Y(_45_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[1]), .B(_45_), .Y(_46_) );
INVX1 INVX1_8 ( .A(i_add_term2[1]), .Y(_47_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term1[1]), .B(_47_), .Y(_48_) );
OAI22X1 OAI22X1_1 ( .A(_42_), .B(_44_), .C(_46_), .D(_48_), .Y(_49_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_50_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_51_) );
NOR2X1 NOR2X1_10 ( .A(_50_), .B(_51_), .Y(_52_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_53_) );
NAND2X1 NAND2X1_9 ( .A(_52_), .B(_53_), .Y(_54_) );
NOR2X1 NOR2X1_11 ( .A(_49_), .B(_54_), .Y(_3_) );
INVX1 INVX1_9 ( .A(_1_), .Y(_55_) );
NAND2X1 NAND2X1_10 ( .A(1'b0), .B(_3_), .Y(_56_) );
OAI21X1 OAI21X1_9 ( .A(_3_), .B(_55_), .C(_56_), .Y(w_cout_1_) );
INVX1 INVX1_10 ( .A(w_cout_1_), .Y(_60_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_61_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_62_) );
NAND3X1 NAND3X1_5 ( .A(_60_), .B(_62_), .C(_61_), .Y(_63_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_57_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_58_) );
OAI21X1 OAI21X1_10 ( .A(_57_), .B(_58_), .C(w_cout_1_), .Y(_59_) );
NAND2X1 NAND2X1_12 ( .A(_59_), .B(_63_), .Y(_0__4_) );
OAI21X1 OAI21X1_11 ( .A(_60_), .B(_57_), .C(_62_), .Y(_5__1_) );
INVX1 INVX1_11 ( .A(_5__3_), .Y(_67_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_68_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_69_) );
NAND3X1 NAND3X1_6 ( .A(_67_), .B(_69_), .C(_68_), .Y(_70_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_64_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_65_) );
OAI21X1 OAI21X1_12 ( .A(_64_), .B(_65_), .C(_5__3_), .Y(_66_) );
NAND2X1 NAND2X1_14 ( .A(_66_), .B(_70_), .Y(_0__7_) );
OAI21X1 OAI21X1_13 ( .A(_67_), .B(_64_), .C(_69_), .Y(_4_) );
INVX1 INVX1_12 ( .A(_5__1_), .Y(_74_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_75_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_76_) );
NAND3X1 NAND3X1_7 ( .A(_74_), .B(_76_), .C(_75_), .Y(_77_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_71_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_72_) );
OAI21X1 OAI21X1_14 ( .A(_71_), .B(_72_), .C(_5__1_), .Y(_73_) );
NAND2X1 NAND2X1_16 ( .A(_73_), .B(_77_), .Y(_0__5_) );
OAI21X1 OAI21X1_15 ( .A(_74_), .B(_71_), .C(_76_), .Y(_5__2_) );
INVX1 INVX1_13 ( .A(_5__2_), .Y(_81_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_82_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_83_) );
NAND3X1 NAND3X1_8 ( .A(_81_), .B(_83_), .C(_82_), .Y(_84_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_78_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_79_) );
OAI21X1 OAI21X1_16 ( .A(_78_), .B(_79_), .C(_5__2_), .Y(_80_) );
NAND2X1 NAND2X1_18 ( .A(_80_), .B(_84_), .Y(_0__6_) );
OAI21X1 OAI21X1_17 ( .A(_81_), .B(_78_), .C(_83_), .Y(_5__3_) );
INVX1 INVX1_14 ( .A(i_add_term1[4]), .Y(_85_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[4]), .B(_85_), .Y(_86_) );
INVX1 INVX1_15 ( .A(i_add_term2[4]), .Y(_87_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term1[4]), .B(_87_), .Y(_88_) );
INVX1 INVX1_16 ( .A(i_add_term1[5]), .Y(_89_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[5]), .B(_89_), .Y(_90_) );
INVX1 INVX1_17 ( .A(i_add_term2[5]), .Y(_91_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term1[5]), .B(_91_), .Y(_92_) );
OAI22X1 OAI22X1_2 ( .A(_86_), .B(_88_), .C(_90_), .D(_92_), .Y(_93_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_94_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_95_) );
NOR2X1 NOR2X1_21 ( .A(_94_), .B(_95_), .Y(_96_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_97_) );
NAND2X1 NAND2X1_19 ( .A(_96_), .B(_97_), .Y(_98_) );
NOR2X1 NOR2X1_22 ( .A(_93_), .B(_98_), .Y(_6_) );
INVX1 INVX1_18 ( .A(_4_), .Y(_99_) );
NAND2X1 NAND2X1_20 ( .A(1'b0), .B(_6_), .Y(_100_) );
OAI21X1 OAI21X1_18 ( .A(_6_), .B(_99_), .C(_100_), .Y(w_cout_2_) );
INVX1 INVX1_19 ( .A(w_cout_2_), .Y(_104_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_105_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_106_) );
NAND3X1 NAND3X1_9 ( .A(_104_), .B(_106_), .C(_105_), .Y(_107_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_101_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_102_) );
OAI21X1 OAI21X1_19 ( .A(_101_), .B(_102_), .C(w_cout_2_), .Y(_103_) );
NAND2X1 NAND2X1_22 ( .A(_103_), .B(_107_), .Y(_0__8_) );
OAI21X1 OAI21X1_20 ( .A(_104_), .B(_101_), .C(_106_), .Y(_8__1_) );
INVX1 INVX1_20 ( .A(_8__3_), .Y(_111_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_112_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_113_) );
NAND3X1 NAND3X1_10 ( .A(_111_), .B(_113_), .C(_112_), .Y(_114_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_108_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_109_) );
OAI21X1 OAI21X1_21 ( .A(_108_), .B(_109_), .C(_8__3_), .Y(_110_) );
NAND2X1 NAND2X1_24 ( .A(_110_), .B(_114_), .Y(_0__11_) );
OAI21X1 OAI21X1_22 ( .A(_111_), .B(_108_), .C(_113_), .Y(_7_) );
INVX1 INVX1_21 ( .A(_8__1_), .Y(_118_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_119_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_120_) );
NAND3X1 NAND3X1_11 ( .A(_118_), .B(_120_), .C(_119_), .Y(_121_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_115_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_116_) );
OAI21X1 OAI21X1_23 ( .A(_115_), .B(_116_), .C(_8__1_), .Y(_117_) );
NAND2X1 NAND2X1_26 ( .A(_117_), .B(_121_), .Y(_0__9_) );
OAI21X1 OAI21X1_24 ( .A(_118_), .B(_115_), .C(_120_), .Y(_8__2_) );
INVX1 INVX1_22 ( .A(_8__2_), .Y(_125_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_126_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_127_) );
NAND3X1 NAND3X1_12 ( .A(_125_), .B(_127_), .C(_126_), .Y(_128_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_122_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_123_) );
OAI21X1 OAI21X1_25 ( .A(_122_), .B(_123_), .C(_8__2_), .Y(_124_) );
NAND2X1 NAND2X1_28 ( .A(_124_), .B(_128_), .Y(_0__10_) );
OAI21X1 OAI21X1_26 ( .A(_125_), .B(_122_), .C(_127_), .Y(_8__3_) );
INVX1 INVX1_23 ( .A(i_add_term1[8]), .Y(_129_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[8]), .B(_129_), .Y(_130_) );
INVX1 INVX1_24 ( .A(i_add_term2[8]), .Y(_131_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term1[8]), .B(_131_), .Y(_132_) );
INVX1 INVX1_25 ( .A(i_add_term1[9]), .Y(_133_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[9]), .B(_133_), .Y(_134_) );
INVX1 INVX1_26 ( .A(i_add_term2[9]), .Y(_135_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term1[9]), .B(_135_), .Y(_136_) );
OAI22X1 OAI22X1_3 ( .A(_130_), .B(_132_), .C(_134_), .D(_136_), .Y(_137_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_138_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_139_) );
NOR2X1 NOR2X1_32 ( .A(_138_), .B(_139_), .Y(_140_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_141_) );
NAND2X1 NAND2X1_29 ( .A(_140_), .B(_141_), .Y(_142_) );
NOR2X1 NOR2X1_33 ( .A(_137_), .B(_142_), .Y(_9_) );
INVX1 INVX1_27 ( .A(_7_), .Y(_143_) );
NAND2X1 NAND2X1_30 ( .A(1'b0), .B(_9_), .Y(_144_) );
OAI21X1 OAI21X1_27 ( .A(_9_), .B(_143_), .C(_144_), .Y(w_cout_3_) );
INVX1 INVX1_28 ( .A(w_cout_3_), .Y(_148_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_149_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_150_) );
NAND3X1 NAND3X1_13 ( .A(_148_), .B(_150_), .C(_149_), .Y(_151_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_145_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_146_) );
OAI21X1 OAI21X1_28 ( .A(_145_), .B(_146_), .C(w_cout_3_), .Y(_147_) );
NAND2X1 NAND2X1_32 ( .A(_147_), .B(_151_), .Y(_0__12_) );
OAI21X1 OAI21X1_29 ( .A(_148_), .B(_145_), .C(_150_), .Y(_11__1_) );
INVX1 INVX1_29 ( .A(_11__3_), .Y(_155_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_156_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_157_) );
NAND3X1 NAND3X1_14 ( .A(_155_), .B(_157_), .C(_156_), .Y(_158_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_152_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_153_) );
OAI21X1 OAI21X1_30 ( .A(_152_), .B(_153_), .C(_11__3_), .Y(_154_) );
NAND2X1 NAND2X1_34 ( .A(_154_), .B(_158_), .Y(_0__15_) );
OAI21X1 OAI21X1_31 ( .A(_155_), .B(_152_), .C(_157_), .Y(_10_) );
INVX1 INVX1_30 ( .A(_11__1_), .Y(_162_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_163_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_164_) );
NAND3X1 NAND3X1_15 ( .A(_162_), .B(_164_), .C(_163_), .Y(_165_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_159_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_160_) );
OAI21X1 OAI21X1_32 ( .A(_159_), .B(_160_), .C(_11__1_), .Y(_161_) );
NAND2X1 NAND2X1_36 ( .A(_161_), .B(_165_), .Y(_0__13_) );
OAI21X1 OAI21X1_33 ( .A(_162_), .B(_159_), .C(_164_), .Y(_11__2_) );
INVX1 INVX1_31 ( .A(_11__2_), .Y(_169_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_170_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_171_) );
NAND3X1 NAND3X1_16 ( .A(_169_), .B(_171_), .C(_170_), .Y(_172_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_166_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_167_) );
OAI21X1 OAI21X1_34 ( .A(_166_), .B(_167_), .C(_11__2_), .Y(_168_) );
NAND2X1 NAND2X1_38 ( .A(_168_), .B(_172_), .Y(_0__14_) );
OAI21X1 OAI21X1_35 ( .A(_169_), .B(_166_), .C(_171_), .Y(_11__3_) );
INVX1 INVX1_32 ( .A(i_add_term1[12]), .Y(_173_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[12]), .B(_173_), .Y(_174_) );
INVX1 INVX1_33 ( .A(i_add_term2[12]), .Y(_175_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term1[12]), .B(_175_), .Y(_176_) );
INVX1 INVX1_34 ( .A(i_add_term1[13]), .Y(_177_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[13]), .B(_177_), .Y(_178_) );
INVX1 INVX1_35 ( .A(i_add_term2[13]), .Y(_179_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term1[13]), .B(_179_), .Y(_180_) );
OAI22X1 OAI22X1_4 ( .A(_174_), .B(_176_), .C(_178_), .D(_180_), .Y(_181_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_182_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_183_) );
NOR2X1 NOR2X1_43 ( .A(_182_), .B(_183_), .Y(_184_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_185_) );
NAND2X1 NAND2X1_39 ( .A(_184_), .B(_185_), .Y(_186_) );
NOR2X1 NOR2X1_44 ( .A(_181_), .B(_186_), .Y(_12_) );
INVX1 INVX1_36 ( .A(_10_), .Y(_187_) );
NAND2X1 NAND2X1_40 ( .A(1'b0), .B(_12_), .Y(_188_) );
OAI21X1 OAI21X1_36 ( .A(_12_), .B(_187_), .C(_188_), .Y(cskip3_inst_cin) );
INVX1 INVX1_37 ( .A(cskip3_inst_cin), .Y(_192_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_193_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_194_) );
NAND3X1 NAND3X1_17 ( .A(_192_), .B(_194_), .C(_193_), .Y(_195_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_189_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_190_) );
OAI21X1 OAI21X1_37 ( .A(_189_), .B(_190_), .C(cskip3_inst_cin), .Y(_191_) );
NAND2X1 NAND2X1_42 ( .A(_191_), .B(_195_), .Y(cskip3_inst_rca0_fa0_o_sum) );
OAI21X1 OAI21X1_38 ( .A(_192_), .B(_189_), .C(_194_), .Y(cskip3_inst_rca0_fa0_o_carry) );
INVX1 INVX1_38 ( .A(cskip3_inst_rca0_fa0_o_carry), .Y(_199_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_200_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_201_) );
NAND3X1 NAND3X1_18 ( .A(_199_), .B(_201_), .C(_200_), .Y(_202_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_196_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_197_) );
OAI21X1 OAI21X1_39 ( .A(_196_), .B(_197_), .C(cskip3_inst_rca0_fa0_o_carry), .Y(_198_) );
NAND2X1 NAND2X1_44 ( .A(_198_), .B(_202_), .Y(cskip3_inst_rca0_fa1_o_sum) );
OAI21X1 OAI21X1_40 ( .A(_199_), .B(_196_), .C(_201_), .Y(cskip3_inst_rca0_fa1_o_carry) );
INVX1 INVX1_39 ( .A(cskip3_inst_rca0_fa1_o_carry), .Y(_206_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_207_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_208_) );
NAND3X1 NAND3X1_19 ( .A(_206_), .B(_208_), .C(_207_), .Y(_209_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_203_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_204_) );
OAI21X1 OAI21X1_41 ( .A(_203_), .B(_204_), .C(cskip3_inst_rca0_fa1_o_carry), .Y(_205_) );
NAND2X1 NAND2X1_46 ( .A(_205_), .B(_209_), .Y(cskip3_inst_rca0_fa2_o_sum) );
OAI21X1 OAI21X1_42 ( .A(_206_), .B(_203_), .C(_208_), .Y(cskip3_inst_cout0) );
OR2X2 OR2X2_20 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_213_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_214_) );
NAND2X1 NAND2X1_48 ( .A(_214_), .B(_213_), .Y(_210_) );
XNOR2X1 XNOR2X1_1 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_211_) );
XNOR2X1 XNOR2X1_2 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_212_) );
NOR3X1 NOR3X1_1 ( .A(_210_), .B(_211_), .C(_212_), .Y(cskip3_inst_skip0_P) );
INVX1 INVX1_40 ( .A(cskip3_inst_cout0), .Y(_215_) );
NAND2X1 NAND2X1_49 ( .A(1'b0), .B(cskip3_inst_skip0_P), .Y(_216_) );
OAI21X1 OAI21X1_43 ( .A(cskip3_inst_skip0_P), .B(_215_), .C(_216_), .Y(w_cout_5_) );
BUFX2 BUFX2_21 ( .A(cskip3_inst_rca0_fa0_o_sum), .Y(_0__16_) );
BUFX2 BUFX2_22 ( .A(cskip3_inst_rca0_fa1_o_sum), .Y(_0__17_) );
BUFX2 BUFX2_23 ( .A(cskip3_inst_rca0_fa2_o_sum), .Y(_0__18_) );
BUFX2 BUFX2_24 ( .A(1'b0), .Y(w_cout_0_) );
BUFX2 BUFX2_25 ( .A(cskip3_inst_cin), .Y(w_cout_4_) );
endmodule
