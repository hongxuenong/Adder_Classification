module CSkipA_51bit ( gnd, vdd, i_add_term1, i_add_term2, sum, cout);

input gnd, vdd;
output cout;
input [50:0] i_add_term1;
input [50:0] i_add_term2;
output [50:0] sum;

NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_322_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_323_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_323_), .C(_20__2_), .Y(_324_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_328_), .Y(_0__26_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_322_), .C(_327_), .Y(_20__3_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[24]), .Y(_329_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(_329_), .Y(_330_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .Y(_331_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[24]), .B(_331_), .Y(_332_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[25]), .Y(_333_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(_333_), .Y(_334_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .Y(_335_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[25]), .B(_335_), .Y(_336_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_332_), .C(_334_), .D(_336_), .Y(_337_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_338_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_339_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_339_), .Y(_340_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_341_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_341_), .Y(_342_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_342_), .Y(_21_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_343_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_21_), .Y(_344_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_343_), .C(_344_), .Y(w_cout_7_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .Y(_348_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_349_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_350_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_350_), .C(_349_), .Y(_351_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_345_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_346_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_346_), .C(w_cout_7_), .Y(_347_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_351_), .Y(_0__28_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_345_), .C(_350_), .Y(_23__1_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_23__3_), .Y(_355_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_356_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_357_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_357_), .C(_356_), .Y(_358_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_352_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_353_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_353_), .C(_23__3_), .Y(_354_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_358_), .Y(_0__31_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_352_), .C(_357_), .Y(_22_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_23__1_), .Y(_362_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_363_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_364_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_364_), .C(_363_), .Y(_365_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_359_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_360_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_360_), .C(_23__1_), .Y(_361_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_365_), .Y(_0__29_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_359_), .C(_364_), .Y(_23__2_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_23__2_), .Y(_369_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_370_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_371_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_371_), .C(_370_), .Y(_372_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_366_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_367_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_367_), .C(_23__2_), .Y(_368_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_372_), .Y(_0__30_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_366_), .C(_371_), .Y(_23__3_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[28]), .Y(_373_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(_373_), .Y(_374_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .Y(_375_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[28]), .B(_375_), .Y(_376_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[29]), .Y(_377_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(_377_), .Y(_378_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .Y(_379_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[29]), .B(_379_), .Y(_380_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_376_), .C(_378_), .D(_380_), .Y(_381_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_382_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_383_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_382_), .B(_383_), .Y(_384_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_385_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_385_), .Y(_386_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_386_), .Y(_24_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_387_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_24_), .Y(_388_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_387_), .C(_388_), .Y(w_cout_8_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .Y(_392_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_393_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_394_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_392_), .B(_394_), .C(_393_), .Y(_395_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_389_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_390_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_390_), .C(w_cout_8_), .Y(_391_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_395_), .Y(_0__32_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_392_), .B(_389_), .C(_394_), .Y(_26__1_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_26__3_), .Y(_399_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_400_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_401_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_401_), .C(_400_), .Y(_402_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_396_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_397_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_397_), .C(_26__3_), .Y(_398_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_402_), .Y(_0__35_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_396_), .C(_401_), .Y(_25_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_26__1_), .Y(_406_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_407_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_408_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_406_), .B(_408_), .C(_407_), .Y(_409_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_403_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_404_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_404_), .C(_26__1_), .Y(_405_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_409_), .Y(_0__33_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_406_), .B(_403_), .C(_408_), .Y(_26__2_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_26__2_), .Y(_413_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_414_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_415_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_415_), .C(_414_), .Y(_416_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_410_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_411_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(_411_), .C(_26__2_), .Y(_412_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_416_), .Y(_0__34_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_410_), .C(_415_), .Y(_26__3_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[32]), .Y(_417_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(_417_), .Y(_418_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .Y(_419_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[32]), .B(_419_), .Y(_420_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[33]), .Y(_421_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(_421_), .Y(_422_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .Y(_423_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[33]), .B(_423_), .Y(_424_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_420_), .C(_422_), .D(_424_), .Y(_425_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_426_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_427_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_427_), .Y(_428_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_429_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_429_), .Y(_430_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(_430_), .Y(_27_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(_431_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_27_), .Y(_432_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_431_), .C(_432_), .Y(w_cout_9_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .Y(_436_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_437_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_438_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_438_), .C(_437_), .Y(_439_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_433_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_434_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_434_), .C(w_cout_9_), .Y(_435_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_439_), .Y(_0__36_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_433_), .C(_438_), .Y(_29__1_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_29__3_), .Y(_443_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_444_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_445_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_445_), .C(_444_), .Y(_446_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_440_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_441_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_441_), .C(_29__3_), .Y(_442_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_446_), .Y(_0__39_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_440_), .C(_445_), .Y(_28_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_29__1_), .Y(_450_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_451_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_452_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_452_), .C(_451_), .Y(_453_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_447_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_448_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_448_), .C(_29__1_), .Y(_449_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_453_), .Y(_0__37_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_447_), .C(_452_), .Y(_29__2_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_29__2_), .Y(_457_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_458_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_459_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_459_), .C(_458_), .Y(_460_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_454_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_455_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_454_), .B(_455_), .C(_29__2_), .Y(_456_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_456_), .B(_460_), .Y(_0__38_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_454_), .C(_459_), .Y(_29__3_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[36]), .Y(_461_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(_461_), .Y(_462_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .Y(_463_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[36]), .B(_463_), .Y(_464_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[37]), .Y(_465_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(_465_), .Y(_466_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .Y(_467_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[37]), .B(_467_), .Y(_468_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_462_), .B(_464_), .C(_466_), .D(_468_), .Y(_469_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_470_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_471_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_470_), .B(_471_), .Y(_472_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_473_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_473_), .Y(_474_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_474_), .Y(_30_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_28_), .Y(_475_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_30_), .Y(_476_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_475_), .C(_476_), .Y(w_cout_10_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .Y(_480_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_481_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_482_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_482_), .C(_481_), .Y(_483_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_477_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_478_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_477_), .B(_478_), .C(w_cout_10_), .Y(_479_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_483_), .Y(_0__40_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_477_), .C(_482_), .Y(_32__1_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_32__3_), .Y(_487_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_488_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_489_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_489_), .C(_488_), .Y(_490_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_484_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_485_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_484_), .B(_485_), .C(_32__3_), .Y(_486_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_490_), .Y(_0__43_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_484_), .C(_489_), .Y(_31_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_32__1_), .Y(_494_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_495_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_496_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_496_), .C(_495_), .Y(_497_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_491_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_492_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_492_), .C(_32__1_), .Y(_493_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_497_), .Y(_0__41_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_491_), .C(_496_), .Y(_32__2_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_32__2_), .Y(_501_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_502_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_503_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_501_), .B(_503_), .C(_502_), .Y(_504_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_498_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_499_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_499_), .C(_32__2_), .Y(_500_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_504_), .Y(_0__42_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_501_), .B(_498_), .C(_503_), .Y(_32__3_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[40]), .Y(_505_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(_505_), .Y(_506_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .Y(_507_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[40]), .B(_507_), .Y(_508_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[41]), .Y(_509_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(_509_), .Y(_510_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .Y(_511_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[41]), .B(_511_), .Y(_512_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_508_), .C(_510_), .D(_512_), .Y(_513_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_514_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_515_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_515_), .Y(_516_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_517_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_517_), .Y(_518_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_518_), .Y(_33_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_31_), .Y(_519_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_33_), .Y(_520_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_519_), .C(_520_), .Y(w_cout_11_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .Y(_524_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_525_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_526_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_526_), .C(_525_), .Y(_527_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_521_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_522_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_522_), .C(w_cout_11_), .Y(_523_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_527_), .Y(_0__44_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_521_), .C(_526_), .Y(_35__1_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_35__3_), .Y(_531_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_532_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_533_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_533_), .C(_532_), .Y(_534_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_528_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_529_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_529_), .C(_35__3_), .Y(_530_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_534_), .Y(_0__47_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_528_), .C(_533_), .Y(_34_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_35__1_), .Y(_538_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_539_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_540_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_540_), .C(_539_), .Y(_541_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_535_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_536_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_536_), .C(_35__1_), .Y(_537_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_541_), .Y(_0__45_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_535_), .C(_540_), .Y(_35__2_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_35__2_), .Y(_545_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_546_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_547_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_547_), .C(_546_), .Y(_548_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_542_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_543_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_542_), .B(_543_), .C(_35__2_), .Y(_544_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_548_), .Y(_0__46_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_542_), .C(_547_), .Y(_35__3_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[44]), .Y(_549_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(_549_), .Y(_550_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .Y(_551_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[44]), .B(_551_), .Y(_552_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[45]), .Y(_553_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(_553_), .Y(_554_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .Y(_555_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[45]), .B(_555_), .Y(_556_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_550_), .B(_552_), .C(_554_), .D(_556_), .Y(_557_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_558_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_559_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_559_), .Y(_560_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_561_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_560_), .B(_561_), .Y(_562_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_557_), .B(_562_), .Y(_36_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_34_), .Y(_563_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_36_), .Y(_564_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_563_), .C(_564_), .Y(cskip3_inst_cin) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_cin), .Y(_568_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_569_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_570_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_570_), .C(_569_), .Y(_571_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_565_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_566_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_566_), .C(cskip3_inst_cin), .Y(_567_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_567_), .B(_571_), .Y(cskip3_inst_rca0_fa0_o_sum) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_565_), .C(_570_), .Y(cskip3_inst_rca0_fa0_o_carry) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_rca0_fa0_o_carry), .Y(_575_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_576_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_577_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_577_), .C(_576_), .Y(_578_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_572_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_573_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_573_), .C(cskip3_inst_rca0_fa0_o_carry), .Y(_574_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_574_), .B(_578_), .Y(cskip3_inst_rca0_fa1_o_sum) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_572_), .C(_577_), .Y(cskip3_inst_rca0_fa1_o_carry) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_rca0_fa1_o_carry), .Y(_582_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_583_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_584_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_584_), .C(_583_), .Y(_585_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_579_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_580_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_580_), .C(cskip3_inst_rca0_fa1_o_carry), .Y(_581_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_581_), .B(_585_), .Y(cskip3_inst_rca0_fa2_o_sum) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_579_), .C(_584_), .Y(cskip3_inst_cout0) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_589_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_590_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_590_), .B(_589_), .Y(_586_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_587_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_588_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_586_), .B(_587_), .C(_588_), .Y(cskip3_inst_skip0_P) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_cout0), .Y(_591_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(cskip3_inst_skip0_P), .Y(_592_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_skip0_P), .B(_591_), .C(_592_), .Y(w_cout_13_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(w_cout_13_), .Y(cout) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_rca0_fa0_o_sum), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_rca0_fa1_o_sum), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_rca0_fa2_o_sum), .Y(sum[50]) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_40_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_41_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_42_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_42_), .C(_41_), .Y(_43_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_37_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_38_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_38_), .C(gnd), .Y(_39_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_43_), .Y(_0__0_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_37_), .C(_42_), .Y(_2__1_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_2__3_), .Y(_47_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_48_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_49_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_49_), .C(_48_), .Y(_50_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_44_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_45_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_45_), .C(_2__3_), .Y(_46_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_50_), .Y(_0__3_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_44_), .C(_49_), .Y(_1_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_2__1_), .Y(_54_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_55_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_56_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_56_), .C(_55_), .Y(_57_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_51_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_52_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_52_), .C(_2__1_), .Y(_53_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_57_), .Y(_0__1_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_51_), .C(_56_), .Y(_2__2_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_2__2_), .Y(_61_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_62_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_63_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_63_), .C(_62_), .Y(_64_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_58_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_59_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_59_), .C(_2__2_), .Y(_60_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_64_), .Y(_0__2_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_58_), .C(_63_), .Y(_2__3_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .Y(_65_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(_65_), .Y(_66_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .Y(_67_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .B(_67_), .Y(_68_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .Y(_69_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(_69_), .Y(_70_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .Y(_71_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .B(_71_), .Y(_72_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_68_), .C(_70_), .D(_72_), .Y(_73_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_74_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_75_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_75_), .Y(_76_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_77_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_77_), .Y(_78_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_78_), .Y(_3_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_79_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_3_), .Y(_80_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_79_), .C(_80_), .Y(w_cout_1_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .Y(_84_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_85_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_86_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_86_), .C(_85_), .Y(_87_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_81_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_82_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_82_), .C(w_cout_1_), .Y(_83_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_87_), .Y(_0__4_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_81_), .C(_86_), .Y(_5__1_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_5__3_), .Y(_91_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_92_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_93_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_93_), .C(_92_), .Y(_94_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_88_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_89_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_89_), .C(_5__3_), .Y(_90_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_94_), .Y(_0__7_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_88_), .C(_93_), .Y(_4_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_5__1_), .Y(_98_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_99_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_100_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_100_), .C(_99_), .Y(_101_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_95_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_96_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_96_), .C(_5__1_), .Y(_97_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_101_), .Y(_0__5_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_95_), .C(_100_), .Y(_5__2_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_5__2_), .Y(_105_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_106_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_107_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_107_), .C(_106_), .Y(_108_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_102_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_103_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_103_), .C(_5__2_), .Y(_104_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_108_), .Y(_0__6_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_102_), .C(_107_), .Y(_5__3_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[4]), .Y(_109_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(_109_), .Y(_110_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .Y(_111_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[4]), .B(_111_), .Y(_112_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[5]), .Y(_113_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(_113_), .Y(_114_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .Y(_115_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[5]), .B(_115_), .Y(_116_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_112_), .C(_114_), .D(_116_), .Y(_117_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_118_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_119_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_119_), .Y(_120_) );
XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_121_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_121_), .Y(_122_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_122_), .Y(_6_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(_123_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_6_), .Y(_124_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_123_), .C(_124_), .Y(w_cout_2_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .Y(_128_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_129_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_130_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_130_), .C(_129_), .Y(_131_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_125_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_126_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_126_), .C(w_cout_2_), .Y(_127_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_131_), .Y(_0__8_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_125_), .C(_130_), .Y(_8__1_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_8__3_), .Y(_135_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_136_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_137_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_137_), .C(_136_), .Y(_138_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_132_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_133_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_133_), .C(_8__3_), .Y(_134_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_138_), .Y(_0__11_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_132_), .C(_137_), .Y(_7_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_8__1_), .Y(_142_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_143_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_144_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_144_), .C(_143_), .Y(_145_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_139_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_140_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_140_), .C(_8__1_), .Y(_141_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_145_), .Y(_0__9_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_139_), .C(_144_), .Y(_8__2_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_8__2_), .Y(_149_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_150_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_151_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_151_), .C(_150_), .Y(_152_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_146_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_147_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_147_), .C(_8__2_), .Y(_148_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_152_), .Y(_0__10_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_146_), .C(_151_), .Y(_8__3_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[8]), .Y(_153_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(_153_), .Y(_154_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .Y(_155_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[8]), .B(_155_), .Y(_156_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[9]), .Y(_157_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(_157_), .Y(_158_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .Y(_159_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[9]), .B(_159_), .Y(_160_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_156_), .C(_158_), .D(_160_), .Y(_161_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_162_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_163_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_163_), .Y(_164_) );
XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_165_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_165_), .Y(_166_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_166_), .Y(_9_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_167_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_9_), .Y(_168_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_167_), .C(_168_), .Y(w_cout_3_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .Y(_172_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_173_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_174_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_174_), .C(_173_), .Y(_175_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_169_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_170_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_170_), .C(w_cout_3_), .Y(_171_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_175_), .Y(_0__12_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_169_), .C(_174_), .Y(_11__1_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_11__3_), .Y(_179_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_180_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_181_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_181_), .C(_180_), .Y(_182_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_176_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_177_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_177_), .C(_11__3_), .Y(_178_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_182_), .Y(_0__15_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_176_), .C(_181_), .Y(_10_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(_11__1_), .Y(_186_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_187_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_188_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_188_), .C(_187_), .Y(_189_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_183_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_184_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_184_), .C(_11__1_), .Y(_185_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_189_), .Y(_0__13_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_183_), .C(_188_), .Y(_11__2_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_11__2_), .Y(_193_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_194_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_195_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_195_), .C(_194_), .Y(_196_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_190_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_191_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_191_), .C(_11__2_), .Y(_192_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(_196_), .Y(_0__14_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_190_), .C(_195_), .Y(_11__3_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[12]), .Y(_197_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(_197_), .Y(_198_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .Y(_199_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[12]), .B(_199_), .Y(_200_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[13]), .Y(_201_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(_201_), .Y(_202_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .Y(_203_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[13]), .B(_203_), .Y(_204_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_200_), .C(_202_), .D(_204_), .Y(_205_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_206_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_207_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_207_), .Y(_208_) );
XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_209_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_209_), .Y(_210_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_210_), .Y(_12_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(_211_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_12_), .Y(_212_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_211_), .C(_212_), .Y(w_cout_4_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .Y(_216_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_217_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_218_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_218_), .C(_217_), .Y(_219_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_213_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_214_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_214_), .C(w_cout_4_), .Y(_215_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_219_), .Y(_0__16_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_213_), .C(_218_), .Y(_14__1_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(_14__3_), .Y(_223_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_224_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_225_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_225_), .C(_224_), .Y(_226_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_220_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_221_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_221_), .C(_14__3_), .Y(_222_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_226_), .Y(_0__19_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_220_), .C(_225_), .Y(_13_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(_14__1_), .Y(_230_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_231_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_232_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_232_), .C(_231_), .Y(_233_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_227_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_228_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_228_), .C(_14__1_), .Y(_229_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_233_), .Y(_0__17_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_227_), .C(_232_), .Y(_14__2_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_14__2_), .Y(_237_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_238_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_239_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_239_), .C(_238_), .Y(_240_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_234_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_235_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_235_), .C(_14__2_), .Y(_236_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_240_), .Y(_0__18_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_234_), .C(_239_), .Y(_14__3_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[16]), .Y(_241_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(_241_), .Y(_242_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .Y(_243_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[16]), .B(_243_), .Y(_244_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[17]), .Y(_245_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(_245_), .Y(_246_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .Y(_247_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[17]), .B(_247_), .Y(_248_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_244_), .C(_246_), .D(_248_), .Y(_249_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_250_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_251_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_251_), .Y(_252_) );
XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_253_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_253_), .Y(_254_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_254_), .Y(_15_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_255_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_15_), .Y(_256_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_255_), .C(_256_), .Y(w_cout_5_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .Y(_260_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_261_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_262_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_262_), .C(_261_), .Y(_263_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_257_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_258_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_258_), .C(w_cout_5_), .Y(_259_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_263_), .Y(_0__20_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_257_), .C(_262_), .Y(_17__1_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(_17__3_), .Y(_267_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_268_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_269_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_269_), .C(_268_), .Y(_270_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_264_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_265_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_265_), .C(_17__3_), .Y(_266_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_270_), .Y(_0__23_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_264_), .C(_269_), .Y(_16_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(_17__1_), .Y(_274_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_275_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_276_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_276_), .C(_275_), .Y(_277_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_271_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_272_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_272_), .C(_17__1_), .Y(_273_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_277_), .Y(_0__21_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_271_), .C(_276_), .Y(_17__2_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_17__2_), .Y(_281_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_282_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_283_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_283_), .C(_282_), .Y(_284_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_278_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_279_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_279_), .C(_17__2_), .Y(_280_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_284_), .Y(_0__22_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_278_), .C(_283_), .Y(_17__3_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[20]), .Y(_285_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(_285_), .Y(_286_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .Y(_287_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[20]), .B(_287_), .Y(_288_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[21]), .Y(_289_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(_289_), .Y(_290_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .Y(_291_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[21]), .B(_291_), .Y(_292_) );
OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_288_), .C(_290_), .D(_292_), .Y(_293_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_294_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_295_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_295_), .Y(_296_) );
XOR2X1 XOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_297_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_297_), .Y(_298_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_298_), .Y(_18_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_299_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_18_), .Y(_300_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_299_), .C(_300_), .Y(w_cout_6_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .Y(_304_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_305_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_306_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_306_), .C(_305_), .Y(_307_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_301_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_302_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_302_), .C(w_cout_6_), .Y(_303_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_307_), .Y(_0__24_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_301_), .C(_306_), .Y(_20__1_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(_20__3_), .Y(_311_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_312_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_313_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_313_), .C(_312_), .Y(_314_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_308_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_309_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_309_), .C(_20__3_), .Y(_310_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_314_), .Y(_0__27_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_308_), .C(_313_), .Y(_19_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_20__1_), .Y(_318_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_319_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_320_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_320_), .C(_319_), .Y(_321_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_315_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_316_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_316_), .C(_20__1_), .Y(_317_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_321_), .Y(_0__25_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_315_), .C(_320_), .Y(_20__2_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(_20__2_), .Y(_325_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_326_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_327_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_327_), .C(_326_), .Y(_328_) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_rca0_fa0_o_sum), .Y(_0__48_) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_rca0_fa1_o_sum), .Y(_0__49_) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_rca0_fa2_o_sum), .Y(_0__50_) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(cskip3_inst_cin), .Y(w_cout_12_) );
endmodule
