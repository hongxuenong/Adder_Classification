module CSkipA_32bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [31:0] i_add_term1;
input [31:0] i_add_term2;
output [31:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX2 BUFX2_1 ( .A(w_cout_7_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
INVX1 INVX1_1 ( .A(skip0_cin_next), .Y(_25_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_26_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_27_) );
NAND3X1 NAND3X1_1 ( .A(_25_), .B(_27_), .C(_26_), .Y(_28_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_22_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_23_) );
OAI21X1 OAI21X1_1 ( .A(_22_), .B(_23_), .C(skip0_cin_next), .Y(_24_) );
NAND2X1 NAND2X1_2 ( .A(_24_), .B(_28_), .Y(_0__4_) );
OAI21X1 OAI21X1_2 ( .A(_25_), .B(_22_), .C(_27_), .Y(_2__1_) );
INVX1 INVX1_2 ( .A(_2__3_), .Y(_32_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_33_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_34_) );
NAND3X1 NAND3X1_2 ( .A(_32_), .B(_34_), .C(_33_), .Y(_35_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_29_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_30_) );
OAI21X1 OAI21X1_3 ( .A(_29_), .B(_30_), .C(_2__3_), .Y(_31_) );
NAND2X1 NAND2X1_4 ( .A(_31_), .B(_35_), .Y(_0__7_) );
OAI21X1 OAI21X1_4 ( .A(_32_), .B(_29_), .C(_34_), .Y(_1_) );
INVX1 INVX1_3 ( .A(_2__1_), .Y(_39_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_40_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_41_) );
NAND3X1 NAND3X1_3 ( .A(_39_), .B(_41_), .C(_40_), .Y(_42_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_36_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_37_) );
OAI21X1 OAI21X1_5 ( .A(_36_), .B(_37_), .C(_2__1_), .Y(_38_) );
NAND2X1 NAND2X1_6 ( .A(_38_), .B(_42_), .Y(_0__5_) );
OAI21X1 OAI21X1_6 ( .A(_39_), .B(_36_), .C(_41_), .Y(_2__2_) );
INVX1 INVX1_4 ( .A(_2__2_), .Y(_46_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_47_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_48_) );
NAND3X1 NAND3X1_4 ( .A(_46_), .B(_48_), .C(_47_), .Y(_49_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_43_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_44_) );
OAI21X1 OAI21X1_7 ( .A(_43_), .B(_44_), .C(_2__2_), .Y(_45_) );
NAND2X1 NAND2X1_8 ( .A(_45_), .B(_49_), .Y(_0__6_) );
OAI21X1 OAI21X1_8 ( .A(_46_), .B(_43_), .C(_48_), .Y(_2__3_) );
INVX1 INVX1_5 ( .A(i_add_term1[4]), .Y(_50_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[4]), .B(_50_), .Y(_51_) );
INVX1 INVX1_6 ( .A(i_add_term2[4]), .Y(_52_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term1[4]), .B(_52_), .Y(_53_) );
INVX1 INVX1_7 ( .A(i_add_term1[5]), .Y(_54_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[5]), .B(_54_), .Y(_55_) );
INVX1 INVX1_8 ( .A(i_add_term2[5]), .Y(_56_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term1[5]), .B(_56_), .Y(_57_) );
OAI22X1 OAI22X1_1 ( .A(_51_), .B(_53_), .C(_55_), .D(_57_), .Y(_58_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_59_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_60_) );
NOR2X1 NOR2X1_10 ( .A(_59_), .B(_60_), .Y(_61_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_62_) );
NAND2X1 NAND2X1_9 ( .A(_61_), .B(_62_), .Y(_63_) );
NOR2X1 NOR2X1_11 ( .A(_58_), .B(_63_), .Y(_3_) );
INVX1 INVX1_9 ( .A(_1_), .Y(_64_) );
NAND2X1 NAND2X1_10 ( .A(gnd), .B(_3_), .Y(_65_) );
OAI21X1 OAI21X1_9 ( .A(_3_), .B(_64_), .C(_65_), .Y(w_cout_1_) );
INVX1 INVX1_10 ( .A(w_cout_1_), .Y(_69_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_70_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_71_) );
NAND3X1 NAND3X1_5 ( .A(_69_), .B(_71_), .C(_70_), .Y(_72_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_66_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_67_) );
OAI21X1 OAI21X1_10 ( .A(_66_), .B(_67_), .C(w_cout_1_), .Y(_68_) );
NAND2X1 NAND2X1_12 ( .A(_68_), .B(_72_), .Y(_0__8_) );
OAI21X1 OAI21X1_11 ( .A(_69_), .B(_66_), .C(_71_), .Y(_5__1_) );
INVX1 INVX1_11 ( .A(_5__3_), .Y(_76_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_77_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_78_) );
NAND3X1 NAND3X1_6 ( .A(_76_), .B(_78_), .C(_77_), .Y(_79_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_73_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_74_) );
OAI21X1 OAI21X1_12 ( .A(_73_), .B(_74_), .C(_5__3_), .Y(_75_) );
NAND2X1 NAND2X1_14 ( .A(_75_), .B(_79_), .Y(_0__11_) );
OAI21X1 OAI21X1_13 ( .A(_76_), .B(_73_), .C(_78_), .Y(_4_) );
INVX1 INVX1_12 ( .A(_5__1_), .Y(_83_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_84_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_85_) );
NAND3X1 NAND3X1_7 ( .A(_83_), .B(_85_), .C(_84_), .Y(_86_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_80_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_81_) );
OAI21X1 OAI21X1_14 ( .A(_80_), .B(_81_), .C(_5__1_), .Y(_82_) );
NAND2X1 NAND2X1_16 ( .A(_82_), .B(_86_), .Y(_0__9_) );
OAI21X1 OAI21X1_15 ( .A(_83_), .B(_80_), .C(_85_), .Y(_5__2_) );
INVX1 INVX1_13 ( .A(_5__2_), .Y(_90_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_91_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_92_) );
NAND3X1 NAND3X1_8 ( .A(_90_), .B(_92_), .C(_91_), .Y(_93_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_87_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_88_) );
OAI21X1 OAI21X1_16 ( .A(_87_), .B(_88_), .C(_5__2_), .Y(_89_) );
NAND2X1 NAND2X1_18 ( .A(_89_), .B(_93_), .Y(_0__10_) );
OAI21X1 OAI21X1_17 ( .A(_90_), .B(_87_), .C(_92_), .Y(_5__3_) );
INVX1 INVX1_14 ( .A(i_add_term1[8]), .Y(_94_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[8]), .B(_94_), .Y(_95_) );
INVX1 INVX1_15 ( .A(i_add_term2[8]), .Y(_96_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term1[8]), .B(_96_), .Y(_97_) );
INVX1 INVX1_16 ( .A(i_add_term1[9]), .Y(_98_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[9]), .B(_98_), .Y(_99_) );
INVX1 INVX1_17 ( .A(i_add_term2[9]), .Y(_100_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term1[9]), .B(_100_), .Y(_101_) );
OAI22X1 OAI22X1_2 ( .A(_95_), .B(_97_), .C(_99_), .D(_101_), .Y(_102_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_103_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_104_) );
NOR2X1 NOR2X1_21 ( .A(_103_), .B(_104_), .Y(_105_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_106_) );
NAND2X1 NAND2X1_19 ( .A(_105_), .B(_106_), .Y(_107_) );
NOR2X1 NOR2X1_22 ( .A(_102_), .B(_107_), .Y(_6_) );
INVX1 INVX1_18 ( .A(_4_), .Y(_108_) );
NAND2X1 NAND2X1_20 ( .A(gnd), .B(_6_), .Y(_109_) );
OAI21X1 OAI21X1_18 ( .A(_6_), .B(_108_), .C(_109_), .Y(w_cout_2_) );
INVX1 INVX1_19 ( .A(w_cout_2_), .Y(_113_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_114_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_115_) );
NAND3X1 NAND3X1_9 ( .A(_113_), .B(_115_), .C(_114_), .Y(_116_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_110_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_111_) );
OAI21X1 OAI21X1_19 ( .A(_110_), .B(_111_), .C(w_cout_2_), .Y(_112_) );
NAND2X1 NAND2X1_22 ( .A(_112_), .B(_116_), .Y(_0__12_) );
OAI21X1 OAI21X1_20 ( .A(_113_), .B(_110_), .C(_115_), .Y(_8__1_) );
INVX1 INVX1_20 ( .A(_8__3_), .Y(_120_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_121_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_122_) );
NAND3X1 NAND3X1_10 ( .A(_120_), .B(_122_), .C(_121_), .Y(_123_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_117_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_118_) );
OAI21X1 OAI21X1_21 ( .A(_117_), .B(_118_), .C(_8__3_), .Y(_119_) );
NAND2X1 NAND2X1_24 ( .A(_119_), .B(_123_), .Y(_0__15_) );
OAI21X1 OAI21X1_22 ( .A(_120_), .B(_117_), .C(_122_), .Y(_7_) );
INVX1 INVX1_21 ( .A(_8__1_), .Y(_127_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_128_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_129_) );
NAND3X1 NAND3X1_11 ( .A(_127_), .B(_129_), .C(_128_), .Y(_130_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_124_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_125_) );
OAI21X1 OAI21X1_23 ( .A(_124_), .B(_125_), .C(_8__1_), .Y(_126_) );
NAND2X1 NAND2X1_26 ( .A(_126_), .B(_130_), .Y(_0__13_) );
OAI21X1 OAI21X1_24 ( .A(_127_), .B(_124_), .C(_129_), .Y(_8__2_) );
INVX1 INVX1_22 ( .A(_8__2_), .Y(_134_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_135_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_136_) );
NAND3X1 NAND3X1_12 ( .A(_134_), .B(_136_), .C(_135_), .Y(_137_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_131_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_132_) );
OAI21X1 OAI21X1_25 ( .A(_131_), .B(_132_), .C(_8__2_), .Y(_133_) );
NAND2X1 NAND2X1_28 ( .A(_133_), .B(_137_), .Y(_0__14_) );
OAI21X1 OAI21X1_26 ( .A(_134_), .B(_131_), .C(_136_), .Y(_8__3_) );
INVX1 INVX1_23 ( .A(i_add_term1[12]), .Y(_138_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[12]), .B(_138_), .Y(_139_) );
INVX1 INVX1_24 ( .A(i_add_term2[12]), .Y(_140_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term1[12]), .B(_140_), .Y(_141_) );
INVX1 INVX1_25 ( .A(i_add_term1[13]), .Y(_142_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[13]), .B(_142_), .Y(_143_) );
INVX1 INVX1_26 ( .A(i_add_term2[13]), .Y(_144_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term1[13]), .B(_144_), .Y(_145_) );
OAI22X1 OAI22X1_3 ( .A(_139_), .B(_141_), .C(_143_), .D(_145_), .Y(_146_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_147_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_148_) );
NOR2X1 NOR2X1_32 ( .A(_147_), .B(_148_), .Y(_149_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_150_) );
NAND2X1 NAND2X1_29 ( .A(_149_), .B(_150_), .Y(_151_) );
NOR2X1 NOR2X1_33 ( .A(_146_), .B(_151_), .Y(_9_) );
INVX1 INVX1_27 ( .A(_7_), .Y(_152_) );
NAND2X1 NAND2X1_30 ( .A(gnd), .B(_9_), .Y(_153_) );
OAI21X1 OAI21X1_27 ( .A(_9_), .B(_152_), .C(_153_), .Y(w_cout_3_) );
INVX1 INVX1_28 ( .A(w_cout_3_), .Y(_157_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_158_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_159_) );
NAND3X1 NAND3X1_13 ( .A(_157_), .B(_159_), .C(_158_), .Y(_160_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_154_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_155_) );
OAI21X1 OAI21X1_28 ( .A(_154_), .B(_155_), .C(w_cout_3_), .Y(_156_) );
NAND2X1 NAND2X1_32 ( .A(_156_), .B(_160_), .Y(_0__16_) );
OAI21X1 OAI21X1_29 ( .A(_157_), .B(_154_), .C(_159_), .Y(_11__1_) );
INVX1 INVX1_29 ( .A(_11__3_), .Y(_164_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_165_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_166_) );
NAND3X1 NAND3X1_14 ( .A(_164_), .B(_166_), .C(_165_), .Y(_167_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_161_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_162_) );
OAI21X1 OAI21X1_30 ( .A(_161_), .B(_162_), .C(_11__3_), .Y(_163_) );
NAND2X1 NAND2X1_34 ( .A(_163_), .B(_167_), .Y(_0__19_) );
OAI21X1 OAI21X1_31 ( .A(_164_), .B(_161_), .C(_166_), .Y(_10_) );
INVX1 INVX1_30 ( .A(_11__1_), .Y(_171_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_172_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_173_) );
NAND3X1 NAND3X1_15 ( .A(_171_), .B(_173_), .C(_172_), .Y(_174_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_168_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_169_) );
OAI21X1 OAI21X1_32 ( .A(_168_), .B(_169_), .C(_11__1_), .Y(_170_) );
NAND2X1 NAND2X1_36 ( .A(_170_), .B(_174_), .Y(_0__17_) );
OAI21X1 OAI21X1_33 ( .A(_171_), .B(_168_), .C(_173_), .Y(_11__2_) );
INVX1 INVX1_31 ( .A(_11__2_), .Y(_178_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_179_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_180_) );
NAND3X1 NAND3X1_16 ( .A(_178_), .B(_180_), .C(_179_), .Y(_181_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_175_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_176_) );
OAI21X1 OAI21X1_34 ( .A(_175_), .B(_176_), .C(_11__2_), .Y(_177_) );
NAND2X1 NAND2X1_38 ( .A(_177_), .B(_181_), .Y(_0__18_) );
OAI21X1 OAI21X1_35 ( .A(_178_), .B(_175_), .C(_180_), .Y(_11__3_) );
INVX1 INVX1_32 ( .A(i_add_term1[16]), .Y(_182_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[16]), .B(_182_), .Y(_183_) );
INVX1 INVX1_33 ( .A(i_add_term2[16]), .Y(_184_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term1[16]), .B(_184_), .Y(_185_) );
INVX1 INVX1_34 ( .A(i_add_term1[17]), .Y(_186_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[17]), .B(_186_), .Y(_187_) );
INVX1 INVX1_35 ( .A(i_add_term2[17]), .Y(_188_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term1[17]), .B(_188_), .Y(_189_) );
OAI22X1 OAI22X1_4 ( .A(_183_), .B(_185_), .C(_187_), .D(_189_), .Y(_190_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_191_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_192_) );
NOR2X1 NOR2X1_43 ( .A(_191_), .B(_192_), .Y(_193_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_194_) );
NAND2X1 NAND2X1_39 ( .A(_193_), .B(_194_), .Y(_195_) );
NOR2X1 NOR2X1_44 ( .A(_190_), .B(_195_), .Y(_12_) );
INVX1 INVX1_36 ( .A(_10_), .Y(_196_) );
NAND2X1 NAND2X1_40 ( .A(gnd), .B(_12_), .Y(_197_) );
OAI21X1 OAI21X1_36 ( .A(_12_), .B(_196_), .C(_197_), .Y(w_cout_4_) );
INVX1 INVX1_37 ( .A(w_cout_4_), .Y(_201_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_202_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_203_) );
NAND3X1 NAND3X1_17 ( .A(_201_), .B(_203_), .C(_202_), .Y(_204_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_198_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_199_) );
OAI21X1 OAI21X1_37 ( .A(_198_), .B(_199_), .C(w_cout_4_), .Y(_200_) );
NAND2X1 NAND2X1_42 ( .A(_200_), .B(_204_), .Y(_0__20_) );
OAI21X1 OAI21X1_38 ( .A(_201_), .B(_198_), .C(_203_), .Y(_14__1_) );
INVX1 INVX1_38 ( .A(_14__3_), .Y(_208_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_209_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_210_) );
NAND3X1 NAND3X1_18 ( .A(_208_), .B(_210_), .C(_209_), .Y(_211_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_205_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_206_) );
OAI21X1 OAI21X1_39 ( .A(_205_), .B(_206_), .C(_14__3_), .Y(_207_) );
NAND2X1 NAND2X1_44 ( .A(_207_), .B(_211_), .Y(_0__23_) );
OAI21X1 OAI21X1_40 ( .A(_208_), .B(_205_), .C(_210_), .Y(_13_) );
INVX1 INVX1_39 ( .A(_14__1_), .Y(_215_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_216_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_217_) );
NAND3X1 NAND3X1_19 ( .A(_215_), .B(_217_), .C(_216_), .Y(_218_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_212_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_213_) );
OAI21X1 OAI21X1_41 ( .A(_212_), .B(_213_), .C(_14__1_), .Y(_214_) );
NAND2X1 NAND2X1_46 ( .A(_214_), .B(_218_), .Y(_0__21_) );
OAI21X1 OAI21X1_42 ( .A(_215_), .B(_212_), .C(_217_), .Y(_14__2_) );
INVX1 INVX1_40 ( .A(_14__2_), .Y(_222_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_223_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_224_) );
NAND3X1 NAND3X1_20 ( .A(_222_), .B(_224_), .C(_223_), .Y(_225_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_219_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_220_) );
OAI21X1 OAI21X1_43 ( .A(_219_), .B(_220_), .C(_14__2_), .Y(_221_) );
NAND2X1 NAND2X1_48 ( .A(_221_), .B(_225_), .Y(_0__22_) );
OAI21X1 OAI21X1_44 ( .A(_222_), .B(_219_), .C(_224_), .Y(_14__3_) );
INVX1 INVX1_41 ( .A(i_add_term1[20]), .Y(_226_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[20]), .B(_226_), .Y(_227_) );
INVX1 INVX1_42 ( .A(i_add_term2[20]), .Y(_228_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term1[20]), .B(_228_), .Y(_229_) );
INVX1 INVX1_43 ( .A(i_add_term1[21]), .Y(_230_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[21]), .B(_230_), .Y(_231_) );
INVX1 INVX1_44 ( .A(i_add_term2[21]), .Y(_232_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term1[21]), .B(_232_), .Y(_233_) );
OAI22X1 OAI22X1_5 ( .A(_227_), .B(_229_), .C(_231_), .D(_233_), .Y(_234_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_235_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_236_) );
NOR2X1 NOR2X1_54 ( .A(_235_), .B(_236_), .Y(_237_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_238_) );
NAND2X1 NAND2X1_49 ( .A(_237_), .B(_238_), .Y(_239_) );
NOR2X1 NOR2X1_55 ( .A(_234_), .B(_239_), .Y(_15_) );
INVX1 INVX1_45 ( .A(_13_), .Y(_240_) );
NAND2X1 NAND2X1_50 ( .A(gnd), .B(_15_), .Y(_241_) );
OAI21X1 OAI21X1_45 ( .A(_15_), .B(_240_), .C(_241_), .Y(w_cout_5_) );
INVX1 INVX1_46 ( .A(w_cout_5_), .Y(_245_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_246_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_247_) );
NAND3X1 NAND3X1_21 ( .A(_245_), .B(_247_), .C(_246_), .Y(_248_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_242_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_243_) );
OAI21X1 OAI21X1_46 ( .A(_242_), .B(_243_), .C(w_cout_5_), .Y(_244_) );
NAND2X1 NAND2X1_52 ( .A(_244_), .B(_248_), .Y(_0__24_) );
OAI21X1 OAI21X1_47 ( .A(_245_), .B(_242_), .C(_247_), .Y(_17__1_) );
INVX1 INVX1_47 ( .A(_17__3_), .Y(_252_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_253_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_254_) );
NAND3X1 NAND3X1_22 ( .A(_252_), .B(_254_), .C(_253_), .Y(_255_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_249_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_250_) );
OAI21X1 OAI21X1_48 ( .A(_249_), .B(_250_), .C(_17__3_), .Y(_251_) );
NAND2X1 NAND2X1_54 ( .A(_251_), .B(_255_), .Y(_0__27_) );
OAI21X1 OAI21X1_49 ( .A(_252_), .B(_249_), .C(_254_), .Y(_16_) );
INVX1 INVX1_48 ( .A(_17__1_), .Y(_259_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_260_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_261_) );
NAND3X1 NAND3X1_23 ( .A(_259_), .B(_261_), .C(_260_), .Y(_262_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_256_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_257_) );
OAI21X1 OAI21X1_50 ( .A(_256_), .B(_257_), .C(_17__1_), .Y(_258_) );
NAND2X1 NAND2X1_56 ( .A(_258_), .B(_262_), .Y(_0__25_) );
OAI21X1 OAI21X1_51 ( .A(_259_), .B(_256_), .C(_261_), .Y(_17__2_) );
INVX1 INVX1_49 ( .A(_17__2_), .Y(_266_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_267_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_268_) );
NAND3X1 NAND3X1_24 ( .A(_266_), .B(_268_), .C(_267_), .Y(_269_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_263_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_264_) );
OAI21X1 OAI21X1_52 ( .A(_263_), .B(_264_), .C(_17__2_), .Y(_265_) );
NAND2X1 NAND2X1_58 ( .A(_265_), .B(_269_), .Y(_0__26_) );
OAI21X1 OAI21X1_53 ( .A(_266_), .B(_263_), .C(_268_), .Y(_17__3_) );
INVX1 INVX1_50 ( .A(i_add_term1[24]), .Y(_270_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[24]), .B(_270_), .Y(_271_) );
INVX1 INVX1_51 ( .A(i_add_term2[24]), .Y(_272_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term1[24]), .B(_272_), .Y(_273_) );
INVX1 INVX1_52 ( .A(i_add_term1[25]), .Y(_274_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[25]), .B(_274_), .Y(_275_) );
INVX1 INVX1_53 ( .A(i_add_term2[25]), .Y(_276_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term1[25]), .B(_276_), .Y(_277_) );
OAI22X1 OAI22X1_6 ( .A(_271_), .B(_273_), .C(_275_), .D(_277_), .Y(_278_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_279_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_280_) );
NOR2X1 NOR2X1_65 ( .A(_279_), .B(_280_), .Y(_281_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_282_) );
NAND2X1 NAND2X1_59 ( .A(_281_), .B(_282_), .Y(_283_) );
NOR2X1 NOR2X1_66 ( .A(_278_), .B(_283_), .Y(_18_) );
INVX1 INVX1_54 ( .A(_16_), .Y(_284_) );
NAND2X1 NAND2X1_60 ( .A(gnd), .B(_18_), .Y(_285_) );
OAI21X1 OAI21X1_54 ( .A(_18_), .B(_284_), .C(_285_), .Y(w_cout_6_) );
INVX1 INVX1_55 ( .A(w_cout_6_), .Y(_289_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_290_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_291_) );
NAND3X1 NAND3X1_25 ( .A(_289_), .B(_291_), .C(_290_), .Y(_292_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_286_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_287_) );
OAI21X1 OAI21X1_55 ( .A(_286_), .B(_287_), .C(w_cout_6_), .Y(_288_) );
NAND2X1 NAND2X1_62 ( .A(_288_), .B(_292_), .Y(_0__28_) );
OAI21X1 OAI21X1_56 ( .A(_289_), .B(_286_), .C(_291_), .Y(_20__1_) );
INVX1 INVX1_56 ( .A(_20__3_), .Y(_296_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_297_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_298_) );
NAND3X1 NAND3X1_26 ( .A(_296_), .B(_298_), .C(_297_), .Y(_299_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_293_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_294_) );
OAI21X1 OAI21X1_57 ( .A(_293_), .B(_294_), .C(_20__3_), .Y(_295_) );
NAND2X1 NAND2X1_64 ( .A(_295_), .B(_299_), .Y(_0__31_) );
OAI21X1 OAI21X1_58 ( .A(_296_), .B(_293_), .C(_298_), .Y(_19_) );
INVX1 INVX1_57 ( .A(_20__1_), .Y(_303_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_304_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_305_) );
NAND3X1 NAND3X1_27 ( .A(_303_), .B(_305_), .C(_304_), .Y(_306_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_300_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_301_) );
OAI21X1 OAI21X1_59 ( .A(_300_), .B(_301_), .C(_20__1_), .Y(_302_) );
NAND2X1 NAND2X1_66 ( .A(_302_), .B(_306_), .Y(_0__29_) );
OAI21X1 OAI21X1_60 ( .A(_303_), .B(_300_), .C(_305_), .Y(_20__2_) );
INVX1 INVX1_58 ( .A(_20__2_), .Y(_310_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_311_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_312_) );
NAND3X1 NAND3X1_28 ( .A(_310_), .B(_312_), .C(_311_), .Y(_313_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_307_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_308_) );
OAI21X1 OAI21X1_61 ( .A(_307_), .B(_308_), .C(_20__2_), .Y(_309_) );
NAND2X1 NAND2X1_68 ( .A(_309_), .B(_313_), .Y(_0__30_) );
OAI21X1 OAI21X1_62 ( .A(_310_), .B(_307_), .C(_312_), .Y(_20__3_) );
INVX1 INVX1_59 ( .A(i_add_term1[28]), .Y(_314_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[28]), .B(_314_), .Y(_315_) );
INVX1 INVX1_60 ( .A(i_add_term2[28]), .Y(_316_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term1[28]), .B(_316_), .Y(_317_) );
INVX1 INVX1_61 ( .A(i_add_term1[29]), .Y(_318_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[29]), .B(_318_), .Y(_319_) );
INVX1 INVX1_62 ( .A(i_add_term2[29]), .Y(_320_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term1[29]), .B(_320_), .Y(_321_) );
OAI22X1 OAI22X1_7 ( .A(_315_), .B(_317_), .C(_319_), .D(_321_), .Y(_322_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_323_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_324_) );
NOR2X1 NOR2X1_76 ( .A(_323_), .B(_324_), .Y(_325_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_326_) );
NAND2X1 NAND2X1_69 ( .A(_325_), .B(_326_), .Y(_327_) );
NOR2X1 NOR2X1_77 ( .A(_322_), .B(_327_), .Y(_21_) );
INVX1 INVX1_63 ( .A(_19_), .Y(_328_) );
NAND2X1 NAND2X1_70 ( .A(gnd), .B(_21_), .Y(_329_) );
OAI21X1 OAI21X1_63 ( .A(_21_), .B(_328_), .C(_329_), .Y(w_cout_7_) );
INVX1 INVX1_64 ( .A(gnd), .Y(_333_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_334_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_335_) );
NAND3X1 NAND3X1_29 ( .A(_333_), .B(_335_), .C(_334_), .Y(_336_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_330_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_331_) );
OAI21X1 OAI21X1_64 ( .A(_330_), .B(_331_), .C(gnd), .Y(_332_) );
NAND2X1 NAND2X1_72 ( .A(_332_), .B(_336_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_65 ( .A(_333_), .B(_330_), .C(_335_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_65 ( .A(rca_inst_fa3_i_carry), .Y(_340_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_341_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_342_) );
NAND3X1 NAND3X1_30 ( .A(_340_), .B(_342_), .C(_341_), .Y(_343_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_337_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_338_) );
OAI21X1 OAI21X1_66 ( .A(_337_), .B(_338_), .C(rca_inst_fa3_i_carry), .Y(_339_) );
NAND2X1 NAND2X1_74 ( .A(_339_), .B(_343_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_67 ( .A(_340_), .B(_337_), .C(_342_), .Y(cout0) );
INVX1 INVX1_66 ( .A(rca_inst_fa0_o_carry), .Y(_347_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_348_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_349_) );
NAND3X1 NAND3X1_31 ( .A(_347_), .B(_349_), .C(_348_), .Y(_350_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_344_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_345_) );
OAI21X1 OAI21X1_68 ( .A(_344_), .B(_345_), .C(rca_inst_fa0_o_carry), .Y(_346_) );
NAND2X1 NAND2X1_76 ( .A(_346_), .B(_350_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_69 ( .A(_347_), .B(_344_), .C(_349_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_67 ( .A(rca_inst_fa_1__o_carry), .Y(_354_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_355_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_356_) );
NAND3X1 NAND3X1_32 ( .A(_354_), .B(_356_), .C(_355_), .Y(_357_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_351_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_352_) );
OAI21X1 OAI21X1_70 ( .A(_351_), .B(_352_), .C(rca_inst_fa_1__o_carry), .Y(_353_) );
NAND2X1 NAND2X1_78 ( .A(_353_), .B(_357_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_71 ( .A(_354_), .B(_351_), .C(_356_), .Y(rca_inst_fa3_i_carry) );
INVX1 INVX1_68 ( .A(i_add_term1[0]), .Y(_358_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[0]), .B(_358_), .Y(_359_) );
INVX1 INVX1_69 ( .A(i_add_term2[0]), .Y(_360_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term1[0]), .B(_360_), .Y(_361_) );
INVX1 INVX1_70 ( .A(i_add_term1[1]), .Y(_362_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[1]), .B(_362_), .Y(_363_) );
INVX1 INVX1_71 ( .A(i_add_term2[1]), .Y(_364_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term1[1]), .B(_364_), .Y(_365_) );
OAI22X1 OAI22X1_8 ( .A(_359_), .B(_361_), .C(_363_), .D(_365_), .Y(_366_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_367_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_368_) );
NOR2X1 NOR2X1_87 ( .A(_367_), .B(_368_), .Y(_369_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_370_) );
NAND2X1 NAND2X1_79 ( .A(_369_), .B(_370_), .Y(_371_) );
NOR2X1 NOR2X1_88 ( .A(_366_), .B(_371_), .Y(skip0_P) );
INVX1 INVX1_72 ( .A(cout0), .Y(_372_) );
NAND2X1 NAND2X1_80 ( .A(gnd), .B(skip0_P), .Y(_373_) );
OAI21X1 OAI21X1_72 ( .A(skip0_P), .B(_372_), .C(_373_), .Y(skip0_cin_next) );
BUFX2 BUFX2_34 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_35 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_36 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_37 ( .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_38 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
