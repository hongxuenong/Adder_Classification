module cla_33bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [32:0] i_add1;
input [32:0] i_add2;
output [33:0] o_result;

NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_7_), .Y(w_C_3_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .Y(_8_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add1[3]), .Y(_9_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_9_), .Y(_10_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_11_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_11_), .C(_7_), .Y(_12_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_10_), .Y(w_C_4_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_14_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_14_), .C(_12_), .Y(_15_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_15_), .Y(w_C_5_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_16_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_17_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_18_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_18_), .C(_15_), .Y(_19_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_17_), .Y(w_C_6_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .Y(_20_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add1[6]), .Y(_21_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_23_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_23_), .C(_19_), .Y(_24_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .C(_24_), .Y(w_C_7_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .Y(_25_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(_26_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_27_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(_28_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_28_), .C(_24_), .Y(_29_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .C(_29_), .Y(_30_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(w_C_8_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .Y(_31_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add1[8]), .Y(_32_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_33_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_33_), .Y(_34_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_35_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_35_), .Y(_36_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_36_), .C(_29_), .Y(_37_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_32_), .C(_37_), .Y(w_C_9_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_32_), .Y(_38_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_38_), .Y(_39_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_40_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_40_), .Y(_41_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_41_), .C(_37_), .Y(_42_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .C(_42_), .Y(_43_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(w_C_10_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .Y(_44_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add1[10]), .Y(_45_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_46_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_46_), .Y(_47_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_48_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_48_), .Y(_49_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_49_), .C(_42_), .Y(_50_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_45_), .C(_50_), .Y(w_C_11_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_45_), .Y(_51_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_51_), .Y(_52_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_53_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_53_), .Y(_54_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_54_), .C(_50_), .Y(_55_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .C(_55_), .Y(_56_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_56_), .Y(w_C_12_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .Y(_57_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add1[12]), .Y(_58_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_59_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_59_), .Y(_60_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_61_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_61_), .Y(_62_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_62_), .C(_55_), .Y(_63_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_58_), .C(_63_), .Y(w_C_13_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_58_), .Y(_64_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_64_), .Y(_65_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_66_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_66_), .Y(_67_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_67_), .C(_63_), .Y(_68_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .C(_68_), .Y(_69_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(w_C_14_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .Y(_70_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add1[14]), .Y(_71_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_72_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_72_), .Y(_73_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_74_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_74_), .Y(_75_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_75_), .C(_68_), .Y(_76_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_71_), .C(_76_), .Y(w_C_15_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_71_), .Y(_77_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(_78_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_79_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_79_), .Y(_80_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_80_), .C(_76_), .Y(_81_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .C(_81_), .Y(_82_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_82_), .Y(w_C_16_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .Y(_83_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add1[16]), .Y(_84_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_84_), .Y(_85_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_85_), .Y(_86_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_87_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_87_), .Y(_88_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_89_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_89_), .Y(_90_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_90_), .C(_81_), .Y(_91_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_86_), .Y(_92_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_92_), .Y(w_C_17_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_93_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_93_), .Y(_94_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_94_), .C(_91_), .Y(_95_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .C(_95_), .Y(_96_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_96_), .Y(w_C_18_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .Y(_97_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add1[18]), .Y(_98_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_98_), .Y(_99_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_99_), .Y(_100_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_101_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_101_), .Y(_102_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_103_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_103_), .Y(_104_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_104_), .C(_95_), .Y(_105_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_100_), .Y(_106_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_106_), .Y(w_C_19_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_107_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_107_), .Y(_108_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_108_), .C(_105_), .Y(_109_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .C(_109_), .Y(_110_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_110_), .Y(w_C_20_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .Y(_111_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add1[20]), .Y(_112_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_112_), .Y(_113_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_113_), .Y(_114_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_115_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_115_), .Y(_116_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_117_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_117_), .Y(_118_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_118_), .C(_109_), .Y(_119_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_114_), .Y(_120_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_120_), .Y(w_C_21_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_121_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_121_), .Y(_122_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_122_), .C(_119_), .Y(_123_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .C(_123_), .Y(_124_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_124_), .Y(w_C_22_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .Y(_125_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add1[22]), .Y(_126_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_126_), .Y(_127_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_127_), .Y(_128_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_129_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_129_), .Y(_130_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_131_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_131_), .Y(_132_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_132_), .C(_123_), .Y(_133_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_128_), .Y(_134_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_134_), .Y(w_C_23_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_135_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_135_), .Y(_136_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_136_), .C(_133_), .Y(_137_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .C(_137_), .Y(_138_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(_138_), .Y(w_C_24_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .Y(_139_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add1[24]), .Y(_140_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_140_), .Y(_141_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_141_), .Y(_142_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_143_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_143_), .Y(_144_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_145_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_145_), .Y(_146_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_146_), .C(_137_), .Y(_147_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_142_), .Y(_148_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_148_), .Y(w_C_25_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_149_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_149_), .Y(_150_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_150_), .C(_147_), .Y(_151_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .C(_151_), .Y(_152_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(_152_), .Y(w_C_26_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_153_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_154_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_152_), .C(_153_), .Y(w_C_27_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_155_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_156_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_157_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_154_), .Y(_158_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_158_), .C(_151_), .Y(_159_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_160_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_160_), .C(_159_), .Y(_161_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_155_), .Y(w_C_28_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .Y(_162_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add1[28]), .Y(_163_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_163_), .Y(_164_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_164_), .C(_161_), .Y(_165_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_163_), .C(_165_), .Y(w_C_29_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .Y(_166_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add1[29]), .Y(_167_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_167_), .Y(_168_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_169_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_170_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_170_), .C(_165_), .Y(_171_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_168_), .Y(w_C_30_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .Y(_172_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add1[30]), .Y(_173_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_173_), .Y(_174_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_174_), .C(_171_), .Y(_175_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_173_), .C(_175_), .Y(w_C_31_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_176_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_177_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_178_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_178_), .C(_175_), .Y(_179_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_176_), .Y(w_C_32_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_180_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_181_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_181_), .C(_179_), .Y(_182_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_182_), .Y(w_C_33_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_183__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_183__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_183__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_183__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_183__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_183__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_183__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_183__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_183__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_183__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_183__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_183__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_183__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_183__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_183__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_183__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_183__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_183__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_183__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_183__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_183__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_183__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_183__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_183__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_183__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_183__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_183__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_183__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_183__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_183__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_183__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_183__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_183__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(w_C_33_), .Y(o_result[33]) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_187_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_188_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_189_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(_189_), .C(_188_), .Y(_190_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_184_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_185_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_185_), .C(w_C_4_), .Y(_186_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_190_), .Y(_183__4_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_194_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_195_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_196_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_196_), .C(_195_), .Y(_197_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_191_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_192_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_192_), .C(w_C_5_), .Y(_193_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_197_), .Y(_183__5_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_201_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_202_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_203_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_203_), .C(_202_), .Y(_204_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_198_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_199_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_199_), .C(w_C_6_), .Y(_200_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_204_), .Y(_183__6_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_208_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_209_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_210_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_210_), .C(_209_), .Y(_211_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_205_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_206_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_206_), .C(w_C_7_), .Y(_207_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_211_), .Y(_183__7_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_215_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_216_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_217_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_217_), .C(_216_), .Y(_218_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_212_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_213_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_213_), .C(w_C_8_), .Y(_214_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_218_), .Y(_183__8_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_222_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_223_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_224_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_224_), .C(_223_), .Y(_225_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_219_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_220_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_220_), .C(w_C_9_), .Y(_221_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_225_), .Y(_183__9_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_229_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_230_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_231_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_231_), .C(_230_), .Y(_232_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_226_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_227_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_227_), .C(w_C_10_), .Y(_228_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_232_), .Y(_183__10_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_236_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_237_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_238_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_238_), .C(_237_), .Y(_239_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_233_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_234_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_234_), .C(w_C_11_), .Y(_235_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_239_), .Y(_183__11_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(w_C_12_), .Y(_243_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_244_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_245_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_245_), .C(_244_), .Y(_246_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_240_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_241_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_241_), .C(w_C_12_), .Y(_242_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_246_), .Y(_183__12_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(w_C_13_), .Y(_250_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_251_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_252_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_252_), .C(_251_), .Y(_253_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_247_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_248_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_248_), .C(w_C_13_), .Y(_249_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_253_), .Y(_183__13_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(w_C_14_), .Y(_257_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_258_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_259_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_259_), .C(_258_), .Y(_260_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_254_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_255_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_255_), .C(w_C_14_), .Y(_256_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_260_), .Y(_183__14_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(_264_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_265_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_266_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_266_), .C(_265_), .Y(_267_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_261_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_262_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_262_), .C(w_C_15_), .Y(_263_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_267_), .Y(_183__15_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(w_C_16_), .Y(_271_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_272_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_273_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_273_), .C(_272_), .Y(_274_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_268_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_269_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_269_), .C(w_C_16_), .Y(_270_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_274_), .Y(_183__16_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(w_C_17_), .Y(_278_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_279_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_280_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_280_), .C(_279_), .Y(_281_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_275_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_276_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_276_), .C(w_C_17_), .Y(_277_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_281_), .Y(_183__17_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(w_C_18_), .Y(_285_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_286_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_287_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_287_), .C(_286_), .Y(_288_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_282_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_283_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_283_), .C(w_C_18_), .Y(_284_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_288_), .Y(_183__18_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(w_C_19_), .Y(_292_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_293_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_294_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_292_), .B(_294_), .C(_293_), .Y(_295_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_289_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_290_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_290_), .C(w_C_19_), .Y(_291_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_295_), .Y(_183__19_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(w_C_20_), .Y(_299_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_300_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_301_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_301_), .C(_300_), .Y(_302_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_296_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_297_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_297_), .C(w_C_20_), .Y(_298_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_302_), .Y(_183__20_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(w_C_21_), .Y(_306_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_307_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_308_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_308_), .C(_307_), .Y(_309_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_303_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_304_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_304_), .C(w_C_21_), .Y(_305_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_309_), .Y(_183__21_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(w_C_22_), .Y(_313_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_314_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_315_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_315_), .C(_314_), .Y(_316_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_310_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_311_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_311_), .C(w_C_22_), .Y(_312_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_316_), .Y(_183__22_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(w_C_23_), .Y(_320_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_321_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_322_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_322_), .C(_321_), .Y(_323_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_317_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_318_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_318_), .C(w_C_23_), .Y(_319_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_323_), .Y(_183__23_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(w_C_24_), .Y(_327_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_328_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_329_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_329_), .C(_328_), .Y(_330_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_324_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_325_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_325_), .C(w_C_24_), .Y(_326_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_330_), .Y(_183__24_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(w_C_25_), .Y(_334_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_335_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_336_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_336_), .C(_335_), .Y(_337_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_331_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_332_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_332_), .C(w_C_25_), .Y(_333_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_337_), .Y(_183__25_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(w_C_26_), .Y(_341_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_342_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_343_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_343_), .C(_342_), .Y(_344_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_338_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_339_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_339_), .C(w_C_26_), .Y(_340_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_344_), .Y(_183__26_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(w_C_27_), .Y(_348_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_349_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_350_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_350_), .C(_349_), .Y(_351_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_345_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_346_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_346_), .C(w_C_27_), .Y(_347_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_351_), .Y(_183__27_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(w_C_28_), .Y(_355_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_356_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_357_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_357_), .C(_356_), .Y(_358_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_352_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_353_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_353_), .C(w_C_28_), .Y(_354_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_358_), .Y(_183__28_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(w_C_29_), .Y(_362_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_363_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_364_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_364_), .C(_363_), .Y(_365_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_359_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_360_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_360_), .C(w_C_29_), .Y(_361_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_365_), .Y(_183__29_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(w_C_30_), .Y(_369_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_370_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_371_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_371_), .C(_370_), .Y(_372_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_366_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_367_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_367_), .C(w_C_30_), .Y(_368_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_372_), .Y(_183__30_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(w_C_31_), .Y(_376_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_377_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_378_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_378_), .C(_377_), .Y(_379_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_373_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_374_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_373_), .B(_374_), .C(w_C_31_), .Y(_375_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_379_), .Y(_183__31_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(w_C_32_), .Y(_383_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_384_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_385_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_385_), .C(_384_), .Y(_386_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_380_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_381_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_381_), .C(w_C_32_), .Y(_382_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_382_), .B(_386_), .Y(_183__32_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_390_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_391_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_392_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_392_), .C(_391_), .Y(_393_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_387_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_388_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_388_), .C(gnd), .Y(_389_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_393_), .Y(_183__0_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_397_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_398_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_399_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_399_), .C(_398_), .Y(_400_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_394_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_395_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_395_), .C(w_C_1_), .Y(_396_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_400_), .Y(_183__1_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_404_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_405_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_406_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_406_), .C(_405_), .Y(_407_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_401_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_402_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_402_), .C(w_C_2_), .Y(_403_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_407_), .Y(_183__2_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_411_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_412_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_413_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_413_), .C(_412_), .Y(_414_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_408_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_409_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_409_), .C(w_C_3_), .Y(_410_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(_414_), .Y(_183__3_) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(w_C_33_), .Y(_183__33_) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
