module cla_63bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [62:0] i_add1;
input [62:0] i_add2;
output [63:0] o_result;

NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_175_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_175_), .Y(_176_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_176_), .C(_167_), .Y(_177_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_172_), .Y(_178_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_178_), .Y(w_C_29_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_179_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_179_), .Y(_180_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_180_), .C(_177_), .Y(_181_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .C(_181_), .Y(_182_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_182_), .Y(w_C_30_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .Y(_183_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add1[30]), .Y(_184_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_184_), .Y(_185_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_185_), .Y(_186_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_187_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_187_), .Y(_188_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_189_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_189_), .Y(_190_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_190_), .C(_181_), .Y(_191_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_186_), .Y(_192_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_192_), .Y(w_C_31_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_193_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_193_), .Y(_194_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_194_), .C(_191_), .Y(_195_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .C(_195_), .Y(_196_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_196_), .Y(w_C_32_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .Y(_197_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add1[32]), .Y(_198_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_198_), .Y(_199_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_199_), .Y(_200_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_201_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_201_), .Y(_202_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_203_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_203_), .Y(_204_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_204_), .C(_195_), .Y(_205_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_200_), .Y(_206_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_206_), .Y(w_C_33_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_207_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_207_), .Y(_208_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_208_), .C(_205_), .Y(_209_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .C(_209_), .Y(_210_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_210_), .Y(w_C_34_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .Y(_211_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add1[34]), .Y(_212_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_212_), .Y(_213_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_213_), .Y(_214_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_215_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_215_), .Y(_216_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_217_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_217_), .Y(_218_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_218_), .C(_209_), .Y(_219_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_214_), .Y(_220_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_220_), .Y(w_C_35_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_221_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_221_), .Y(_222_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_222_), .C(_219_), .Y(_223_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .C(_223_), .Y(_224_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_224_), .Y(w_C_36_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .Y(_225_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add1[36]), .Y(_226_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_226_), .Y(_227_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_227_), .Y(_228_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_229_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_229_), .Y(_230_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_231_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_231_), .Y(_232_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_232_), .C(_223_), .Y(_233_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_228_), .Y(_234_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_234_), .Y(w_C_37_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_235_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_235_), .Y(_236_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_236_), .C(_233_), .Y(_237_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .C(_237_), .Y(_238_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_238_), .Y(w_C_38_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .Y(_239_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add1[38]), .Y(_240_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_240_), .Y(_241_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_241_), .Y(_242_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_243_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_243_), .Y(_244_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_245_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_245_), .Y(_246_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_246_), .C(_237_), .Y(_247_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_242_), .Y(_248_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_248_), .Y(w_C_39_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_249_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_249_), .Y(_250_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_250_), .C(_247_), .Y(_251_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .C(_251_), .Y(_252_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_252_), .Y(w_C_40_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .Y(_253_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add1[40]), .Y(_254_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_253_), .B(_254_), .Y(_255_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_255_), .Y(_256_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_257_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_257_), .Y(_258_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_259_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_259_), .Y(_260_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_260_), .C(_251_), .Y(_261_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_256_), .Y(_262_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_262_), .Y(w_C_41_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_263_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_263_), .Y(_264_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_264_), .C(_261_), .Y(_265_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .C(_265_), .Y(_266_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_266_), .Y(w_C_42_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .Y(_267_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add1[42]), .Y(_268_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_268_), .Y(_269_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_269_), .Y(_270_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_271_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_271_), .Y(_272_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_273_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_273_), .Y(_274_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_274_), .C(_265_), .Y(_275_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_270_), .Y(_276_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_276_), .Y(w_C_43_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_277_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_277_), .Y(_278_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_278_), .C(_275_), .Y(_279_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .C(_279_), .Y(_280_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_280_), .Y(w_C_44_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .Y(_281_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add1[44]), .Y(_282_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_282_), .Y(_283_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_283_), .Y(_284_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_285_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_285_), .Y(_286_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_287_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_287_), .Y(_288_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_288_), .C(_279_), .Y(_289_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_284_), .Y(_290_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_290_), .Y(w_C_45_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_291_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_291_), .Y(_292_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_292_), .C(_289_), .Y(_293_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .C(_293_), .Y(_294_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_294_), .Y(w_C_46_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .Y(_295_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add1[46]), .Y(_296_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_296_), .Y(_297_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(_297_), .Y(_298_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_299_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_299_), .Y(_300_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_301_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(_301_), .Y(_302_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_302_), .C(_293_), .Y(_303_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_298_), .Y(_304_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_304_), .Y(w_C_47_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_305_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_305_), .Y(_306_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_306_), .C(_303_), .Y(_307_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .C(_307_), .Y(_308_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_308_), .Y(w_C_48_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .Y(_309_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add1[48]), .Y(_310_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_310_), .Y(_311_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(_311_), .Y(_312_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_313_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_313_), .Y(_314_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_315_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_315_), .Y(_316_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_316_), .C(_307_), .Y(_317_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_312_), .Y(_318_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_318_), .Y(w_C_49_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_319_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_319_), .Y(_320_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_320_), .C(_317_), .Y(_321_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .C(_321_), .Y(_322_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(_322_), .Y(w_C_50_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_323_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_324_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_322_), .C(_323_), .Y(w_C_51_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_325_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_326_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_326_), .Y(_327_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_324_), .Y(_328_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_328_), .C(_321_), .Y(_329_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_330_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_330_), .C(_329_), .Y(_331_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_325_), .Y(w_C_52_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .Y(_332_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add1[52]), .Y(_333_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_333_), .Y(_334_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_334_), .C(_331_), .Y(_335_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_333_), .C(_335_), .Y(w_C_53_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .Y(_336_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add1[53]), .Y(_337_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_337_), .Y(_338_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_339_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_340_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_340_), .C(_335_), .Y(_341_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_338_), .Y(w_C_54_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .Y(_342_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add1[54]), .Y(_343_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_343_), .Y(_344_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_344_), .C(_341_), .Y(_345_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_343_), .C(_345_), .Y(w_C_55_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_346_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(_346_), .Y(_347_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_343_), .Y(_348_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_348_), .Y(_349_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .Y(_350_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add1[55]), .Y(_351_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_351_), .Y(_352_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(_352_), .Y(_353_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_353_), .C(_345_), .Y(_354_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_347_), .Y(w_C_56_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .Y(_355_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add1[56]), .Y(_356_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_357_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(_357_), .Y(_358_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_358_), .C(_354_), .Y(_359_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_356_), .C(_359_), .Y(w_C_57_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .Y(_360_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add1[57]), .Y(_361_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .C(w_C_57_), .Y(_362_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_361_), .C(_362_), .Y(w_C_58_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_361_), .Y(_363_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_363_), .Y(_364_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_365_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(_365_), .Y(_366_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_366_), .C(_362_), .Y(_367_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .C(_367_), .Y(_368_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_368_), .Y(w_C_59_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_369_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_370_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_368_), .C(_369_), .Y(w_C_60_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[60]), .B(i_add1[60]), .Y(_371_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_370_), .Y(_372_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_373_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_373_), .Y(_374_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_356_), .Y(_375_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_375_), .Y(_376_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_364_), .C(_359_), .Y(_377_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_378_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_378_), .Y(_379_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_379_), .C(_377_), .Y(_380_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_369_), .C(_380_), .Y(_381_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[60]), .B(i_add1[60]), .Y(_382_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_382_), .C(_381_), .Y(_383_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_383_), .Y(w_C_61_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[61]), .B(i_add1[61]), .Y(_384_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[61]), .B(i_add1[61]), .Y(_385_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_385_), .C(_383_), .Y(_386_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_384_), .Y(w_C_62_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[62]), .B(i_add1[62]), .Y(_387_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[62]), .B(i_add1[62]), .Y(_388_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_388_), .C(_386_), .Y(_389_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_389_), .Y(w_C_63_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_7_), .Y(w_C_3_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_8_), .C(_7_), .Y(_9_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .C(_9_), .Y(_10_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(w_C_4_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_12_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_13_), .C(_9_), .Y(_14_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_14_), .Y(w_C_5_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_15_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_15_), .C(_14_), .Y(_16_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .C(_16_), .Y(_17_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(_17_), .Y(w_C_6_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .Y(_18_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add1[6]), .Y(_19_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_20_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(_20_), .Y(_21_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_23_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_23_), .C(_16_), .Y(_24_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_19_), .C(_24_), .Y(w_C_7_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_19_), .Y(_25_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(_26_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_27_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_390__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_390__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_390__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_390__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_390__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_390__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_390__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_390__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_390__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_390__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_390__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_390__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_390__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_390__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_390__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_390__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_390__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_390__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_390__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_390__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_390__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_390__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_390__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_390__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_390__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_390__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_390__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_390__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_390__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_390__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_390__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_390__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_390__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_390__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_390__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_390__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_390__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_390__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_390__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_390__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_390__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_390__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_390__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_390__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_390__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_390__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_390__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_390__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_390__48_), .Y(o_result[48]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_390__49_), .Y(o_result[49]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_390__50_), .Y(o_result[50]) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_390__51_), .Y(o_result[51]) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(_390__52_), .Y(o_result[52]) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(_390__53_), .Y(o_result[53]) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(_390__54_), .Y(o_result[54]) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_390__55_), .Y(o_result[55]) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_390__56_), .Y(o_result[56]) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_390__57_), .Y(o_result[57]) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_390__58_), .Y(o_result[58]) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(_390__59_), .Y(o_result[59]) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(_390__60_), .Y(o_result[60]) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(_390__61_), .Y(o_result[61]) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(_390__62_), .Y(o_result[62]) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(w_C_63_), .Y(o_result[63]) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_394_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_395_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_396_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_396_), .C(_395_), .Y(_397_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_391_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_392_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_392_), .C(w_C_4_), .Y(_393_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_397_), .Y(_390__4_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_401_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_402_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_403_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_403_), .C(_402_), .Y(_404_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_398_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_399_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_399_), .C(w_C_5_), .Y(_400_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_400_), .B(_404_), .Y(_390__5_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_408_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_409_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_410_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_410_), .C(_409_), .Y(_411_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_405_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_406_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_406_), .C(w_C_6_), .Y(_407_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_411_), .Y(_390__6_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_415_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_416_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_417_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_415_), .B(_417_), .C(_416_), .Y(_418_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_412_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_413_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_413_), .C(w_C_7_), .Y(_414_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_414_), .B(_418_), .Y(_390__7_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_422_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_423_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_424_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_422_), .B(_424_), .C(_423_), .Y(_425_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_419_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_420_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_420_), .C(w_C_8_), .Y(_421_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_425_), .Y(_390__8_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_429_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_430_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_431_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(_431_), .C(_430_), .Y(_432_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_426_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_427_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_427_), .C(w_C_9_), .Y(_428_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_432_), .Y(_390__9_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_436_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_437_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_438_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_438_), .C(_437_), .Y(_439_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_433_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_434_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_434_), .C(w_C_10_), .Y(_435_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_439_), .Y(_390__10_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_443_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_444_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_445_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_445_), .C(_444_), .Y(_446_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_440_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_441_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_441_), .C(w_C_11_), .Y(_442_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_446_), .Y(_390__11_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(w_C_12_), .Y(_450_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_451_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_452_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_452_), .C(_451_), .Y(_453_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_447_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_448_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_448_), .C(w_C_12_), .Y(_449_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_453_), .Y(_390__12_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(w_C_13_), .Y(_457_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_458_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_459_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_459_), .C(_458_), .Y(_460_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_454_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_455_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_454_), .B(_455_), .C(w_C_13_), .Y(_456_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_456_), .B(_460_), .Y(_390__13_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(w_C_14_), .Y(_464_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_465_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_466_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_466_), .C(_465_), .Y(_467_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_461_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_462_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_462_), .C(w_C_14_), .Y(_463_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_467_), .Y(_390__14_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(_471_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_472_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_473_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_473_), .C(_472_), .Y(_474_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_468_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_469_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_468_), .B(_469_), .C(w_C_15_), .Y(_470_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_470_), .B(_474_), .Y(_390__15_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(w_C_16_), .Y(_478_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_479_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_480_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_480_), .C(_479_), .Y(_481_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_475_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_476_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_476_), .C(w_C_16_), .Y(_477_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_477_), .B(_481_), .Y(_390__16_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(w_C_17_), .Y(_485_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_486_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_487_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_487_), .C(_486_), .Y(_488_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_482_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_483_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_482_), .B(_483_), .C(w_C_17_), .Y(_484_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_484_), .B(_488_), .Y(_390__17_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(w_C_18_), .Y(_492_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_493_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_494_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_492_), .B(_494_), .C(_493_), .Y(_495_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_489_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_490_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_490_), .C(w_C_18_), .Y(_491_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_495_), .Y(_390__18_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(w_C_19_), .Y(_499_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_500_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_501_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_501_), .C(_500_), .Y(_502_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_496_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_497_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_497_), .C(w_C_19_), .Y(_498_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_502_), .Y(_390__19_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(w_C_20_), .Y(_506_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_507_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_508_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_508_), .C(_507_), .Y(_509_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_503_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_504_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_504_), .C(w_C_20_), .Y(_505_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(_509_), .Y(_390__20_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(w_C_21_), .Y(_513_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_514_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_515_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_515_), .C(_514_), .Y(_516_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_510_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_511_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_511_), .C(w_C_21_), .Y(_512_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_516_), .Y(_390__21_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(w_C_22_), .Y(_520_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_521_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_522_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_522_), .C(_521_), .Y(_523_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_517_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_518_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_517_), .B(_518_), .C(w_C_22_), .Y(_519_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_523_), .Y(_390__22_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(w_C_23_), .Y(_527_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_528_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_529_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_529_), .C(_528_), .Y(_530_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_524_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_525_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_525_), .C(w_C_23_), .Y(_526_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_530_), .Y(_390__23_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(w_C_24_), .Y(_534_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_535_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_536_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_536_), .C(_535_), .Y(_537_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_531_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_532_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_532_), .C(w_C_24_), .Y(_533_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_537_), .Y(_390__24_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(w_C_25_), .Y(_541_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_542_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_543_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_541_), .B(_543_), .C(_542_), .Y(_544_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_538_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_539_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_539_), .C(w_C_25_), .Y(_540_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_544_), .Y(_390__25_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(w_C_26_), .Y(_548_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_549_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_550_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_550_), .C(_549_), .Y(_551_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_545_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_546_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_546_), .C(w_C_26_), .Y(_547_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_547_), .B(_551_), .Y(_390__26_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(w_C_27_), .Y(_555_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_556_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_557_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_555_), .B(_557_), .C(_556_), .Y(_558_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_552_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_553_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_552_), .B(_553_), .C(w_C_27_), .Y(_554_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_558_), .Y(_390__27_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(w_C_28_), .Y(_562_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_563_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_564_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_562_), .B(_564_), .C(_563_), .Y(_565_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_559_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_560_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_560_), .C(w_C_28_), .Y(_561_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_565_), .Y(_390__28_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(w_C_29_), .Y(_569_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_570_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_571_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_569_), .B(_571_), .C(_570_), .Y(_572_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_566_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_567_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_567_), .C(w_C_29_), .Y(_568_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_572_), .Y(_390__29_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(w_C_30_), .Y(_576_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_577_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_578_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_576_), .B(_578_), .C(_577_), .Y(_579_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_573_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_574_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_574_), .C(w_C_30_), .Y(_575_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_579_), .Y(_390__30_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(w_C_31_), .Y(_583_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_584_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_585_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_583_), .B(_585_), .C(_584_), .Y(_586_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_580_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_581_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(_581_), .C(w_C_31_), .Y(_582_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_586_), .Y(_390__31_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(w_C_32_), .Y(_590_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_591_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_592_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_590_), .B(_592_), .C(_591_), .Y(_593_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_587_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_588_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(_588_), .C(w_C_32_), .Y(_589_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_589_), .B(_593_), .Y(_390__32_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(w_C_33_), .Y(_597_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_598_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_599_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_597_), .B(_599_), .C(_598_), .Y(_600_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_594_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_595_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_594_), .B(_595_), .C(w_C_33_), .Y(_596_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_600_), .Y(_390__33_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(w_C_34_), .Y(_604_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_605_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_606_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(_606_), .C(_605_), .Y(_607_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_601_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_602_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_601_), .B(_602_), .C(w_C_34_), .Y(_603_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_603_), .B(_607_), .Y(_390__34_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(w_C_35_), .Y(_611_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_612_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_613_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_613_), .C(_612_), .Y(_614_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_608_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_609_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_608_), .B(_609_), .C(w_C_35_), .Y(_610_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_614_), .Y(_390__35_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(w_C_36_), .Y(_618_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_619_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_620_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_618_), .B(_620_), .C(_619_), .Y(_621_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_615_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_616_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(_616_), .C(w_C_36_), .Y(_617_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_617_), .B(_621_), .Y(_390__36_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(w_C_37_), .Y(_625_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_626_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_627_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_625_), .B(_627_), .C(_626_), .Y(_628_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_622_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_623_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_622_), .B(_623_), .C(w_C_37_), .Y(_624_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_624_), .B(_628_), .Y(_390__37_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(w_C_38_), .Y(_632_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_633_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_634_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_632_), .B(_634_), .C(_633_), .Y(_635_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_629_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_630_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_629_), .B(_630_), .C(w_C_38_), .Y(_631_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_631_), .B(_635_), .Y(_390__38_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(w_C_39_), .Y(_639_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_640_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_641_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_641_), .C(_640_), .Y(_642_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_636_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_637_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_636_), .B(_637_), .C(w_C_39_), .Y(_638_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_642_), .Y(_390__39_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(w_C_40_), .Y(_646_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_647_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_648_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_646_), .B(_648_), .C(_647_), .Y(_649_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_643_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_644_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_644_), .C(w_C_40_), .Y(_645_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_645_), .B(_649_), .Y(_390__40_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(w_C_41_), .Y(_653_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_654_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_655_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_653_), .B(_655_), .C(_654_), .Y(_656_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_650_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_651_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(_651_), .C(w_C_41_), .Y(_652_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_656_), .Y(_390__41_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(w_C_42_), .Y(_660_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_661_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_662_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_660_), .B(_662_), .C(_661_), .Y(_663_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_657_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_658_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_657_), .B(_658_), .C(w_C_42_), .Y(_659_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(_663_), .Y(_390__42_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(w_C_43_), .Y(_667_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_668_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_669_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_667_), .B(_669_), .C(_668_), .Y(_670_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_664_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_665_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_665_), .C(w_C_43_), .Y(_666_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_666_), .B(_670_), .Y(_390__43_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(w_C_44_), .Y(_674_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_675_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_676_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_676_), .C(_675_), .Y(_677_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_671_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_672_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_671_), .B(_672_), .C(w_C_44_), .Y(_673_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_673_), .B(_677_), .Y(_390__44_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(w_C_45_), .Y(_681_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_682_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_683_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_681_), .B(_683_), .C(_682_), .Y(_684_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_678_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_679_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_679_), .C(w_C_45_), .Y(_680_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_680_), .B(_684_), .Y(_390__45_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(w_C_46_), .Y(_688_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_689_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_690_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_688_), .B(_690_), .C(_689_), .Y(_691_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_685_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_686_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_686_), .C(w_C_46_), .Y(_687_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_687_), .B(_691_), .Y(_390__46_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(w_C_47_), .Y(_695_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_696_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_697_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_695_), .B(_697_), .C(_696_), .Y(_698_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_692_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_693_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_692_), .B(_693_), .C(w_C_47_), .Y(_694_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_698_), .Y(_390__47_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(w_C_48_), .Y(_702_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_703_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_704_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(_704_), .C(_703_), .Y(_705_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_699_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_700_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_700_), .C(w_C_48_), .Y(_701_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_701_), .B(_705_), .Y(_390__48_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(w_C_49_), .Y(_709_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_710_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_711_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_711_), .C(_710_), .Y(_712_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_706_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_707_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_707_), .C(w_C_49_), .Y(_708_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_708_), .B(_712_), .Y(_390__49_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(w_C_50_), .Y(_716_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_717_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_718_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_716_), .B(_718_), .C(_717_), .Y(_719_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_713_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_714_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_714_), .C(w_C_50_), .Y(_715_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(_719_), .Y(_390__50_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(w_C_51_), .Y(_723_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_724_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_725_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_723_), .B(_725_), .C(_724_), .Y(_726_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_720_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_721_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_720_), .B(_721_), .C(w_C_51_), .Y(_722_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_722_), .B(_726_), .Y(_390__51_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(w_C_52_), .Y(_730_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_731_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_732_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_730_), .B(_732_), .C(_731_), .Y(_733_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_727_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_728_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_727_), .B(_728_), .C(w_C_52_), .Y(_729_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_733_), .Y(_390__52_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(w_C_53_), .Y(_737_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_738_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_739_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_737_), .B(_739_), .C(_738_), .Y(_740_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_734_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_735_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_734_), .B(_735_), .C(w_C_53_), .Y(_736_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_736_), .B(_740_), .Y(_390__53_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(w_C_54_), .Y(_744_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_745_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_746_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_744_), .B(_746_), .C(_745_), .Y(_747_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_741_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_742_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_741_), .B(_742_), .C(w_C_54_), .Y(_743_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_743_), .B(_747_), .Y(_390__54_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(w_C_55_), .Y(_751_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_752_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_753_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_751_), .B(_753_), .C(_752_), .Y(_754_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_748_) );
AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_749_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_748_), .B(_749_), .C(w_C_55_), .Y(_750_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_750_), .B(_754_), .Y(_390__55_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(w_C_56_), .Y(_758_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_759_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_760_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_758_), .B(_760_), .C(_759_), .Y(_761_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_755_) );
AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_756_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_756_), .C(w_C_56_), .Y(_757_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_757_), .B(_761_), .Y(_390__56_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(w_C_57_), .Y(_765_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_766_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_767_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_765_), .B(_767_), .C(_766_), .Y(_768_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_762_) );
AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_763_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_762_), .B(_763_), .C(w_C_57_), .Y(_764_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_764_), .B(_768_), .Y(_390__57_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(w_C_58_), .Y(_772_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_773_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_774_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_772_), .B(_774_), .C(_773_), .Y(_775_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_769_) );
AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_770_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_769_), .B(_770_), .C(w_C_58_), .Y(_771_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_771_), .B(_775_), .Y(_390__58_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(w_C_59_), .Y(_779_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_780_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_781_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_779_), .B(_781_), .C(_780_), .Y(_782_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_776_) );
AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[59]), .B(i_add1[59]), .Y(_777_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_776_), .B(_777_), .C(w_C_59_), .Y(_778_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_778_), .B(_782_), .Y(_390__59_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(w_C_60_), .Y(_786_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[60]), .B(i_add1[60]), .Y(_787_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(i_add2[60]), .B(i_add1[60]), .Y(_788_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(_788_), .C(_787_), .Y(_789_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add2[60]), .B(i_add1[60]), .Y(_783_) );
AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[60]), .B(i_add1[60]), .Y(_784_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(_784_), .C(w_C_60_), .Y(_785_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_789_), .Y(_390__60_) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(w_C_61_), .Y(_793_) );
OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[61]), .B(i_add1[61]), .Y(_794_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(i_add2[61]), .B(i_add1[61]), .Y(_795_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(_795_), .C(_794_), .Y(_796_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add2[61]), .B(i_add1[61]), .Y(_790_) );
AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[61]), .B(i_add1[61]), .Y(_791_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(_791_), .C(w_C_61_), .Y(_792_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_792_), .B(_796_), .Y(_390__61_) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(w_C_62_), .Y(_800_) );
OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[62]), .B(i_add1[62]), .Y(_801_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(i_add2[62]), .B(i_add1[62]), .Y(_802_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_800_), .B(_802_), .C(_801_), .Y(_803_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add2[62]), .B(i_add1[62]), .Y(_797_) );
AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[62]), .B(i_add1[62]), .Y(_798_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_797_), .B(_798_), .C(w_C_62_), .Y(_799_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_799_), .B(_803_), .Y(_390__62_) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_807_) );
OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_808_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_809_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_807_), .B(_809_), .C(_808_), .Y(_810_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_804_) );
AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_805_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_804_), .B(_805_), .C(gnd), .Y(_806_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_806_), .B(_810_), .Y(_390__0_) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_814_) );
OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_815_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_816_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_814_), .B(_816_), .C(_815_), .Y(_817_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_811_) );
AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_812_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_811_), .B(_812_), .C(w_C_1_), .Y(_813_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_813_), .B(_817_), .Y(_390__1_) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_821_) );
OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_822_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_823_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_821_), .B(_823_), .C(_822_), .Y(_824_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_818_) );
AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_819_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_819_), .C(w_C_2_), .Y(_820_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_820_), .B(_824_), .Y(_390__2_) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_828_) );
OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_829_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_830_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_828_), .B(_830_), .C(_829_), .Y(_831_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_825_) );
AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_826_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_825_), .B(_826_), .C(w_C_3_), .Y(_827_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_827_), .B(_831_), .Y(_390__3_) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(_28_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_28_), .C(_24_), .Y(_29_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .C(_29_), .Y(_30_) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(w_C_8_) );
INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .Y(_31_) );
INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(i_add1[8]), .Y(_32_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_33_) );
INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(_33_), .Y(_34_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_35_) );
INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(_35_), .Y(_36_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_36_), .C(_29_), .Y(_37_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_32_), .C(_37_), .Y(w_C_9_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_32_), .Y(_38_) );
INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(_38_), .Y(_39_) );
AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_40_) );
INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(_40_), .Y(_41_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_41_), .C(_37_), .Y(_42_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .C(_42_), .Y(_43_) );
INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(w_C_10_) );
INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .Y(_44_) );
INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(i_add1[10]), .Y(_45_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_46_) );
INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(_46_), .Y(_47_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_48_) );
INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(_48_), .Y(_49_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_49_), .C(_42_), .Y(_50_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_45_), .C(_50_), .Y(w_C_11_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_45_), .Y(_51_) );
INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(_51_), .Y(_52_) );
AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_53_) );
INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(_53_), .Y(_54_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_54_), .C(_50_), .Y(_55_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .C(_55_), .Y(_56_) );
INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(_56_), .Y(w_C_12_) );
INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .Y(_57_) );
INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(i_add1[12]), .Y(_58_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_58_), .Y(_59_) );
INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(_59_), .Y(_60_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_61_) );
INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(_61_), .Y(_62_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_63_) );
INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(_63_), .Y(_64_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_64_), .C(_55_), .Y(_65_) );
AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_60_), .Y(_66_) );
INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(_66_), .Y(w_C_13_) );
AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_67_) );
INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(_67_), .Y(_68_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_68_), .C(_65_), .Y(_69_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .C(_69_), .Y(_70_) );
INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(_70_), .Y(w_C_14_) );
INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .Y(_71_) );
INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(i_add1[14]), .Y(_72_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_72_), .Y(_73_) );
INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(_73_), .Y(_74_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_75_) );
INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(_75_), .Y(_76_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_77_) );
INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(_78_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_78_), .C(_69_), .Y(_79_) );
AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_74_), .Y(_80_) );
INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(_80_), .Y(w_C_15_) );
AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_81_) );
INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(_81_), .Y(_82_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_82_), .C(_79_), .Y(_83_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .C(_83_), .Y(_84_) );
INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(_84_), .Y(w_C_16_) );
INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .Y(_85_) );
INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(i_add1[16]), .Y(_86_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_86_), .Y(_87_) );
INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(_87_), .Y(_88_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_89_) );
INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(_89_), .Y(_90_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_91_) );
INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(_91_), .Y(_92_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_92_), .C(_83_), .Y(_93_) );
AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_88_), .Y(_94_) );
INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(_94_), .Y(w_C_17_) );
AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_95_) );
INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(_95_), .Y(_96_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_96_), .C(_93_), .Y(_97_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .C(_97_), .Y(_98_) );
INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(_98_), .Y(w_C_18_) );
INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .Y(_99_) );
INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(i_add1[18]), .Y(_100_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_100_), .Y(_101_) );
INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(_101_), .Y(_102_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_103_) );
INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(_103_), .Y(_104_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_105_) );
INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(_105_), .Y(_106_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_106_), .C(_97_), .Y(_107_) );
AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_102_), .Y(_108_) );
INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(_108_), .Y(w_C_19_) );
AND2X2 AND2X2_101 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_109_) );
INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(_109_), .Y(_110_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_110_), .C(_107_), .Y(_111_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .C(_111_), .Y(_112_) );
INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(_112_), .Y(w_C_20_) );
INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .Y(_113_) );
INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(i_add1[20]), .Y(_114_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_114_), .Y(_115_) );
INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(_115_), .Y(_116_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_117_) );
INVX1 INVX1_233 ( .gnd(gnd), .vdd(vdd), .A(_117_), .Y(_118_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_119_) );
INVX1 INVX1_234 ( .gnd(gnd), .vdd(vdd), .A(_119_), .Y(_120_) );
NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_120_), .C(_111_), .Y(_121_) );
AND2X2 AND2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_116_), .Y(_122_) );
INVX1 INVX1_235 ( .gnd(gnd), .vdd(vdd), .A(_122_), .Y(w_C_21_) );
AND2X2 AND2X2_103 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_123_) );
INVX1 INVX1_236 ( .gnd(gnd), .vdd(vdd), .A(_123_), .Y(_124_) );
NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_124_), .C(_121_), .Y(_125_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .C(_125_), .Y(_126_) );
INVX1 INVX1_237 ( .gnd(gnd), .vdd(vdd), .A(_126_), .Y(w_C_22_) );
INVX1 INVX1_238 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .Y(_127_) );
INVX1 INVX1_239 ( .gnd(gnd), .vdd(vdd), .A(i_add1[22]), .Y(_128_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_128_), .Y(_129_) );
INVX1 INVX1_240 ( .gnd(gnd), .vdd(vdd), .A(_129_), .Y(_130_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_131_) );
INVX1 INVX1_241 ( .gnd(gnd), .vdd(vdd), .A(_131_), .Y(_132_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_133_) );
INVX1 INVX1_242 ( .gnd(gnd), .vdd(vdd), .A(_133_), .Y(_134_) );
NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_134_), .C(_125_), .Y(_135_) );
AND2X2 AND2X2_104 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_130_), .Y(_136_) );
INVX1 INVX1_243 ( .gnd(gnd), .vdd(vdd), .A(_136_), .Y(w_C_23_) );
AND2X2 AND2X2_105 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_137_) );
INVX1 INVX1_244 ( .gnd(gnd), .vdd(vdd), .A(_137_), .Y(_138_) );
NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_138_), .C(_135_), .Y(_139_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .C(_139_), .Y(_140_) );
INVX1 INVX1_245 ( .gnd(gnd), .vdd(vdd), .A(_140_), .Y(w_C_24_) );
INVX1 INVX1_246 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .Y(_141_) );
INVX1 INVX1_247 ( .gnd(gnd), .vdd(vdd), .A(i_add1[24]), .Y(_142_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_142_), .Y(_143_) );
INVX1 INVX1_248 ( .gnd(gnd), .vdd(vdd), .A(_143_), .Y(_144_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_145_) );
INVX1 INVX1_249 ( .gnd(gnd), .vdd(vdd), .A(_145_), .Y(_146_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_147_) );
INVX1 INVX1_250 ( .gnd(gnd), .vdd(vdd), .A(_147_), .Y(_148_) );
NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_148_), .C(_139_), .Y(_149_) );
AND2X2 AND2X2_106 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_144_), .Y(_150_) );
INVX1 INVX1_251 ( .gnd(gnd), .vdd(vdd), .A(_150_), .Y(w_C_25_) );
AND2X2 AND2X2_107 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_151_) );
INVX1 INVX1_252 ( .gnd(gnd), .vdd(vdd), .A(_151_), .Y(_152_) );
NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_152_), .C(_149_), .Y(_153_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .C(_153_), .Y(_154_) );
INVX1 INVX1_253 ( .gnd(gnd), .vdd(vdd), .A(_154_), .Y(w_C_26_) );
INVX1 INVX1_254 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .Y(_155_) );
INVX1 INVX1_255 ( .gnd(gnd), .vdd(vdd), .A(i_add1[26]), .Y(_156_) );
NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_156_), .Y(_157_) );
INVX1 INVX1_256 ( .gnd(gnd), .vdd(vdd), .A(_157_), .Y(_158_) );
NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_159_) );
INVX1 INVX1_257 ( .gnd(gnd), .vdd(vdd), .A(_159_), .Y(_160_) );
NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_161_) );
INVX1 INVX1_258 ( .gnd(gnd), .vdd(vdd), .A(_161_), .Y(_162_) );
NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_162_), .C(_153_), .Y(_163_) );
AND2X2 AND2X2_108 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_158_), .Y(_164_) );
INVX1 INVX1_259 ( .gnd(gnd), .vdd(vdd), .A(_164_), .Y(w_C_27_) );
AND2X2 AND2X2_109 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_165_) );
INVX1 INVX1_260 ( .gnd(gnd), .vdd(vdd), .A(_165_), .Y(_166_) );
NAND3X1 NAND3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_166_), .C(_163_), .Y(_167_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .C(_167_), .Y(_168_) );
INVX1 INVX1_261 ( .gnd(gnd), .vdd(vdd), .A(_168_), .Y(w_C_28_) );
INVX1 INVX1_262 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .Y(_169_) );
INVX1 INVX1_263 ( .gnd(gnd), .vdd(vdd), .A(i_add1[28]), .Y(_170_) );
NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_170_), .Y(_171_) );
INVX1 INVX1_264 ( .gnd(gnd), .vdd(vdd), .A(_171_), .Y(_172_) );
NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_173_) );
INVX1 INVX1_265 ( .gnd(gnd), .vdd(vdd), .A(_173_), .Y(_174_) );
BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(w_C_63_), .Y(_390__63_) );
BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
