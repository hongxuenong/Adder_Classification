module CSkipA_28bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [27:0] i_add_term1;
input [27:0] i_add_term2;
output [27:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX2 BUFX2_1 ( .A(w_cout_6_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
INVX1 INVX1_1 ( .A(skip0_cin_next), .Y(_22_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_23_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_24_) );
NAND3X1 NAND3X1_1 ( .A(_22_), .B(_24_), .C(_23_), .Y(_25_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_19_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_20_) );
OAI21X1 OAI21X1_1 ( .A(_19_), .B(_20_), .C(skip0_cin_next), .Y(_21_) );
NAND2X1 NAND2X1_2 ( .A(_21_), .B(_25_), .Y(_0__4_) );
OAI21X1 OAI21X1_2 ( .A(_22_), .B(_19_), .C(_24_), .Y(_2__1_) );
INVX1 INVX1_2 ( .A(_2__3_), .Y(_29_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_30_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_31_) );
NAND3X1 NAND3X1_2 ( .A(_29_), .B(_31_), .C(_30_), .Y(_32_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_26_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_27_) );
OAI21X1 OAI21X1_3 ( .A(_26_), .B(_27_), .C(_2__3_), .Y(_28_) );
NAND2X1 NAND2X1_4 ( .A(_28_), .B(_32_), .Y(_0__7_) );
OAI21X1 OAI21X1_4 ( .A(_29_), .B(_26_), .C(_31_), .Y(_1_) );
INVX1 INVX1_3 ( .A(_2__1_), .Y(_36_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_37_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_38_) );
NAND3X1 NAND3X1_3 ( .A(_36_), .B(_38_), .C(_37_), .Y(_39_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_33_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_34_) );
OAI21X1 OAI21X1_5 ( .A(_33_), .B(_34_), .C(_2__1_), .Y(_35_) );
NAND2X1 NAND2X1_6 ( .A(_35_), .B(_39_), .Y(_0__5_) );
OAI21X1 OAI21X1_6 ( .A(_36_), .B(_33_), .C(_38_), .Y(_2__2_) );
INVX1 INVX1_4 ( .A(_2__2_), .Y(_43_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_44_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_45_) );
NAND3X1 NAND3X1_4 ( .A(_43_), .B(_45_), .C(_44_), .Y(_46_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_40_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_41_) );
OAI21X1 OAI21X1_7 ( .A(_40_), .B(_41_), .C(_2__2_), .Y(_42_) );
NAND2X1 NAND2X1_8 ( .A(_42_), .B(_46_), .Y(_0__6_) );
OAI21X1 OAI21X1_8 ( .A(_43_), .B(_40_), .C(_45_), .Y(_2__3_) );
INVX1 INVX1_5 ( .A(i_add_term1[4]), .Y(_47_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[4]), .B(_47_), .Y(_48_) );
INVX1 INVX1_6 ( .A(i_add_term2[4]), .Y(_49_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term1[4]), .B(_49_), .Y(_50_) );
INVX1 INVX1_7 ( .A(i_add_term1[5]), .Y(_51_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[5]), .B(_51_), .Y(_52_) );
INVX1 INVX1_8 ( .A(i_add_term2[5]), .Y(_53_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term1[5]), .B(_53_), .Y(_54_) );
OAI22X1 OAI22X1_1 ( .A(_48_), .B(_50_), .C(_52_), .D(_54_), .Y(_55_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_56_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_57_) );
NOR2X1 NOR2X1_10 ( .A(_56_), .B(_57_), .Y(_58_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_59_) );
NAND2X1 NAND2X1_9 ( .A(_58_), .B(_59_), .Y(_60_) );
NOR2X1 NOR2X1_11 ( .A(_55_), .B(_60_), .Y(_3_) );
INVX1 INVX1_9 ( .A(_1_), .Y(_61_) );
NAND2X1 NAND2X1_10 ( .A(gnd), .B(_3_), .Y(_62_) );
OAI21X1 OAI21X1_9 ( .A(_3_), .B(_61_), .C(_62_), .Y(w_cout_1_) );
INVX1 INVX1_10 ( .A(w_cout_1_), .Y(_66_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_67_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_68_) );
NAND3X1 NAND3X1_5 ( .A(_66_), .B(_68_), .C(_67_), .Y(_69_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_63_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_64_) );
OAI21X1 OAI21X1_10 ( .A(_63_), .B(_64_), .C(w_cout_1_), .Y(_65_) );
NAND2X1 NAND2X1_12 ( .A(_65_), .B(_69_), .Y(_0__8_) );
OAI21X1 OAI21X1_11 ( .A(_66_), .B(_63_), .C(_68_), .Y(_5__1_) );
INVX1 INVX1_11 ( .A(_5__3_), .Y(_73_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_74_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_75_) );
NAND3X1 NAND3X1_6 ( .A(_73_), .B(_75_), .C(_74_), .Y(_76_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_70_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_71_) );
OAI21X1 OAI21X1_12 ( .A(_70_), .B(_71_), .C(_5__3_), .Y(_72_) );
NAND2X1 NAND2X1_14 ( .A(_72_), .B(_76_), .Y(_0__11_) );
OAI21X1 OAI21X1_13 ( .A(_73_), .B(_70_), .C(_75_), .Y(_4_) );
INVX1 INVX1_12 ( .A(_5__1_), .Y(_80_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_81_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_82_) );
NAND3X1 NAND3X1_7 ( .A(_80_), .B(_82_), .C(_81_), .Y(_83_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_77_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_78_) );
OAI21X1 OAI21X1_14 ( .A(_77_), .B(_78_), .C(_5__1_), .Y(_79_) );
NAND2X1 NAND2X1_16 ( .A(_79_), .B(_83_), .Y(_0__9_) );
OAI21X1 OAI21X1_15 ( .A(_80_), .B(_77_), .C(_82_), .Y(_5__2_) );
INVX1 INVX1_13 ( .A(_5__2_), .Y(_87_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_88_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_89_) );
NAND3X1 NAND3X1_8 ( .A(_87_), .B(_89_), .C(_88_), .Y(_90_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_84_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_85_) );
OAI21X1 OAI21X1_16 ( .A(_84_), .B(_85_), .C(_5__2_), .Y(_86_) );
NAND2X1 NAND2X1_18 ( .A(_86_), .B(_90_), .Y(_0__10_) );
OAI21X1 OAI21X1_17 ( .A(_87_), .B(_84_), .C(_89_), .Y(_5__3_) );
INVX1 INVX1_14 ( .A(i_add_term1[8]), .Y(_91_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[8]), .B(_91_), .Y(_92_) );
INVX1 INVX1_15 ( .A(i_add_term2[8]), .Y(_93_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term1[8]), .B(_93_), .Y(_94_) );
INVX1 INVX1_16 ( .A(i_add_term1[9]), .Y(_95_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[9]), .B(_95_), .Y(_96_) );
INVX1 INVX1_17 ( .A(i_add_term2[9]), .Y(_97_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term1[9]), .B(_97_), .Y(_98_) );
OAI22X1 OAI22X1_2 ( .A(_92_), .B(_94_), .C(_96_), .D(_98_), .Y(_99_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_100_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_101_) );
NOR2X1 NOR2X1_21 ( .A(_100_), .B(_101_), .Y(_102_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_103_) );
NAND2X1 NAND2X1_19 ( .A(_102_), .B(_103_), .Y(_104_) );
NOR2X1 NOR2X1_22 ( .A(_99_), .B(_104_), .Y(_6_) );
INVX1 INVX1_18 ( .A(_4_), .Y(_105_) );
NAND2X1 NAND2X1_20 ( .A(gnd), .B(_6_), .Y(_106_) );
OAI21X1 OAI21X1_18 ( .A(_6_), .B(_105_), .C(_106_), .Y(w_cout_2_) );
INVX1 INVX1_19 ( .A(w_cout_2_), .Y(_110_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_111_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_112_) );
NAND3X1 NAND3X1_9 ( .A(_110_), .B(_112_), .C(_111_), .Y(_113_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_107_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_108_) );
OAI21X1 OAI21X1_19 ( .A(_107_), .B(_108_), .C(w_cout_2_), .Y(_109_) );
NAND2X1 NAND2X1_22 ( .A(_109_), .B(_113_), .Y(_0__12_) );
OAI21X1 OAI21X1_20 ( .A(_110_), .B(_107_), .C(_112_), .Y(_8__1_) );
INVX1 INVX1_20 ( .A(_8__3_), .Y(_117_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_118_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_119_) );
NAND3X1 NAND3X1_10 ( .A(_117_), .B(_119_), .C(_118_), .Y(_120_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_114_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_115_) );
OAI21X1 OAI21X1_21 ( .A(_114_), .B(_115_), .C(_8__3_), .Y(_116_) );
NAND2X1 NAND2X1_24 ( .A(_116_), .B(_120_), .Y(_0__15_) );
OAI21X1 OAI21X1_22 ( .A(_117_), .B(_114_), .C(_119_), .Y(_7_) );
INVX1 INVX1_21 ( .A(_8__1_), .Y(_124_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_125_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_126_) );
NAND3X1 NAND3X1_11 ( .A(_124_), .B(_126_), .C(_125_), .Y(_127_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_121_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_122_) );
OAI21X1 OAI21X1_23 ( .A(_121_), .B(_122_), .C(_8__1_), .Y(_123_) );
NAND2X1 NAND2X1_26 ( .A(_123_), .B(_127_), .Y(_0__13_) );
OAI21X1 OAI21X1_24 ( .A(_124_), .B(_121_), .C(_126_), .Y(_8__2_) );
INVX1 INVX1_22 ( .A(_8__2_), .Y(_131_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_132_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_133_) );
NAND3X1 NAND3X1_12 ( .A(_131_), .B(_133_), .C(_132_), .Y(_134_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_128_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_129_) );
OAI21X1 OAI21X1_25 ( .A(_128_), .B(_129_), .C(_8__2_), .Y(_130_) );
NAND2X1 NAND2X1_28 ( .A(_130_), .B(_134_), .Y(_0__14_) );
OAI21X1 OAI21X1_26 ( .A(_131_), .B(_128_), .C(_133_), .Y(_8__3_) );
INVX1 INVX1_23 ( .A(i_add_term1[12]), .Y(_135_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[12]), .B(_135_), .Y(_136_) );
INVX1 INVX1_24 ( .A(i_add_term2[12]), .Y(_137_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term1[12]), .B(_137_), .Y(_138_) );
INVX1 INVX1_25 ( .A(i_add_term1[13]), .Y(_139_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[13]), .B(_139_), .Y(_140_) );
INVX1 INVX1_26 ( .A(i_add_term2[13]), .Y(_141_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term1[13]), .B(_141_), .Y(_142_) );
OAI22X1 OAI22X1_3 ( .A(_136_), .B(_138_), .C(_140_), .D(_142_), .Y(_143_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_144_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_145_) );
NOR2X1 NOR2X1_32 ( .A(_144_), .B(_145_), .Y(_146_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_147_) );
NAND2X1 NAND2X1_29 ( .A(_146_), .B(_147_), .Y(_148_) );
NOR2X1 NOR2X1_33 ( .A(_143_), .B(_148_), .Y(_9_) );
INVX1 INVX1_27 ( .A(_7_), .Y(_149_) );
NAND2X1 NAND2X1_30 ( .A(gnd), .B(_9_), .Y(_150_) );
OAI21X1 OAI21X1_27 ( .A(_9_), .B(_149_), .C(_150_), .Y(w_cout_3_) );
INVX1 INVX1_28 ( .A(w_cout_3_), .Y(_154_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_155_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_156_) );
NAND3X1 NAND3X1_13 ( .A(_154_), .B(_156_), .C(_155_), .Y(_157_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_151_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_152_) );
OAI21X1 OAI21X1_28 ( .A(_151_), .B(_152_), .C(w_cout_3_), .Y(_153_) );
NAND2X1 NAND2X1_32 ( .A(_153_), .B(_157_), .Y(_0__16_) );
OAI21X1 OAI21X1_29 ( .A(_154_), .B(_151_), .C(_156_), .Y(_11__1_) );
INVX1 INVX1_29 ( .A(_11__3_), .Y(_161_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_162_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_163_) );
NAND3X1 NAND3X1_14 ( .A(_161_), .B(_163_), .C(_162_), .Y(_164_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_158_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_159_) );
OAI21X1 OAI21X1_30 ( .A(_158_), .B(_159_), .C(_11__3_), .Y(_160_) );
NAND2X1 NAND2X1_34 ( .A(_160_), .B(_164_), .Y(_0__19_) );
OAI21X1 OAI21X1_31 ( .A(_161_), .B(_158_), .C(_163_), .Y(_10_) );
INVX1 INVX1_30 ( .A(_11__1_), .Y(_168_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_169_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_170_) );
NAND3X1 NAND3X1_15 ( .A(_168_), .B(_170_), .C(_169_), .Y(_171_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_165_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_166_) );
OAI21X1 OAI21X1_32 ( .A(_165_), .B(_166_), .C(_11__1_), .Y(_167_) );
NAND2X1 NAND2X1_36 ( .A(_167_), .B(_171_), .Y(_0__17_) );
OAI21X1 OAI21X1_33 ( .A(_168_), .B(_165_), .C(_170_), .Y(_11__2_) );
INVX1 INVX1_31 ( .A(_11__2_), .Y(_175_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_176_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_177_) );
NAND3X1 NAND3X1_16 ( .A(_175_), .B(_177_), .C(_176_), .Y(_178_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_172_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_173_) );
OAI21X1 OAI21X1_34 ( .A(_172_), .B(_173_), .C(_11__2_), .Y(_174_) );
NAND2X1 NAND2X1_38 ( .A(_174_), .B(_178_), .Y(_0__18_) );
OAI21X1 OAI21X1_35 ( .A(_175_), .B(_172_), .C(_177_), .Y(_11__3_) );
INVX1 INVX1_32 ( .A(i_add_term1[16]), .Y(_179_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[16]), .B(_179_), .Y(_180_) );
INVX1 INVX1_33 ( .A(i_add_term2[16]), .Y(_181_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term1[16]), .B(_181_), .Y(_182_) );
INVX1 INVX1_34 ( .A(i_add_term1[17]), .Y(_183_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[17]), .B(_183_), .Y(_184_) );
INVX1 INVX1_35 ( .A(i_add_term2[17]), .Y(_185_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term1[17]), .B(_185_), .Y(_186_) );
OAI22X1 OAI22X1_4 ( .A(_180_), .B(_182_), .C(_184_), .D(_186_), .Y(_187_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_188_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_189_) );
NOR2X1 NOR2X1_43 ( .A(_188_), .B(_189_), .Y(_190_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_191_) );
NAND2X1 NAND2X1_39 ( .A(_190_), .B(_191_), .Y(_192_) );
NOR2X1 NOR2X1_44 ( .A(_187_), .B(_192_), .Y(_12_) );
INVX1 INVX1_36 ( .A(_10_), .Y(_193_) );
NAND2X1 NAND2X1_40 ( .A(gnd), .B(_12_), .Y(_194_) );
OAI21X1 OAI21X1_36 ( .A(_12_), .B(_193_), .C(_194_), .Y(w_cout_4_) );
INVX1 INVX1_37 ( .A(w_cout_4_), .Y(_198_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_199_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_200_) );
NAND3X1 NAND3X1_17 ( .A(_198_), .B(_200_), .C(_199_), .Y(_201_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_195_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_196_) );
OAI21X1 OAI21X1_37 ( .A(_195_), .B(_196_), .C(w_cout_4_), .Y(_197_) );
NAND2X1 NAND2X1_42 ( .A(_197_), .B(_201_), .Y(_0__20_) );
OAI21X1 OAI21X1_38 ( .A(_198_), .B(_195_), .C(_200_), .Y(_14__1_) );
INVX1 INVX1_38 ( .A(_14__3_), .Y(_205_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_206_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_207_) );
NAND3X1 NAND3X1_18 ( .A(_205_), .B(_207_), .C(_206_), .Y(_208_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_202_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_203_) );
OAI21X1 OAI21X1_39 ( .A(_202_), .B(_203_), .C(_14__3_), .Y(_204_) );
NAND2X1 NAND2X1_44 ( .A(_204_), .B(_208_), .Y(_0__23_) );
OAI21X1 OAI21X1_40 ( .A(_205_), .B(_202_), .C(_207_), .Y(_13_) );
INVX1 INVX1_39 ( .A(_14__1_), .Y(_212_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_213_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_214_) );
NAND3X1 NAND3X1_19 ( .A(_212_), .B(_214_), .C(_213_), .Y(_215_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_209_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_210_) );
OAI21X1 OAI21X1_41 ( .A(_209_), .B(_210_), .C(_14__1_), .Y(_211_) );
NAND2X1 NAND2X1_46 ( .A(_211_), .B(_215_), .Y(_0__21_) );
OAI21X1 OAI21X1_42 ( .A(_212_), .B(_209_), .C(_214_), .Y(_14__2_) );
INVX1 INVX1_40 ( .A(_14__2_), .Y(_219_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_220_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_221_) );
NAND3X1 NAND3X1_20 ( .A(_219_), .B(_221_), .C(_220_), .Y(_222_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_216_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_217_) );
OAI21X1 OAI21X1_43 ( .A(_216_), .B(_217_), .C(_14__2_), .Y(_218_) );
NAND2X1 NAND2X1_48 ( .A(_218_), .B(_222_), .Y(_0__22_) );
OAI21X1 OAI21X1_44 ( .A(_219_), .B(_216_), .C(_221_), .Y(_14__3_) );
INVX1 INVX1_41 ( .A(i_add_term1[20]), .Y(_223_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[20]), .B(_223_), .Y(_224_) );
INVX1 INVX1_42 ( .A(i_add_term2[20]), .Y(_225_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term1[20]), .B(_225_), .Y(_226_) );
INVX1 INVX1_43 ( .A(i_add_term1[21]), .Y(_227_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[21]), .B(_227_), .Y(_228_) );
INVX1 INVX1_44 ( .A(i_add_term2[21]), .Y(_229_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term1[21]), .B(_229_), .Y(_230_) );
OAI22X1 OAI22X1_5 ( .A(_224_), .B(_226_), .C(_228_), .D(_230_), .Y(_231_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_232_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_233_) );
NOR2X1 NOR2X1_54 ( .A(_232_), .B(_233_), .Y(_234_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_235_) );
NAND2X1 NAND2X1_49 ( .A(_234_), .B(_235_), .Y(_236_) );
NOR2X1 NOR2X1_55 ( .A(_231_), .B(_236_), .Y(_15_) );
INVX1 INVX1_45 ( .A(_13_), .Y(_237_) );
NAND2X1 NAND2X1_50 ( .A(gnd), .B(_15_), .Y(_238_) );
OAI21X1 OAI21X1_45 ( .A(_15_), .B(_237_), .C(_238_), .Y(w_cout_5_) );
INVX1 INVX1_46 ( .A(w_cout_5_), .Y(_242_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_243_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_244_) );
NAND3X1 NAND3X1_21 ( .A(_242_), .B(_244_), .C(_243_), .Y(_245_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_239_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_240_) );
OAI21X1 OAI21X1_46 ( .A(_239_), .B(_240_), .C(w_cout_5_), .Y(_241_) );
NAND2X1 NAND2X1_52 ( .A(_241_), .B(_245_), .Y(_0__24_) );
OAI21X1 OAI21X1_47 ( .A(_242_), .B(_239_), .C(_244_), .Y(_17__1_) );
INVX1 INVX1_47 ( .A(_17__3_), .Y(_249_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_250_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_251_) );
NAND3X1 NAND3X1_22 ( .A(_249_), .B(_251_), .C(_250_), .Y(_252_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_246_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_247_) );
OAI21X1 OAI21X1_48 ( .A(_246_), .B(_247_), .C(_17__3_), .Y(_248_) );
NAND2X1 NAND2X1_54 ( .A(_248_), .B(_252_), .Y(_0__27_) );
OAI21X1 OAI21X1_49 ( .A(_249_), .B(_246_), .C(_251_), .Y(_16_) );
INVX1 INVX1_48 ( .A(_17__1_), .Y(_256_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_257_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_258_) );
NAND3X1 NAND3X1_23 ( .A(_256_), .B(_258_), .C(_257_), .Y(_259_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_253_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_254_) );
OAI21X1 OAI21X1_50 ( .A(_253_), .B(_254_), .C(_17__1_), .Y(_255_) );
NAND2X1 NAND2X1_56 ( .A(_255_), .B(_259_), .Y(_0__25_) );
OAI21X1 OAI21X1_51 ( .A(_256_), .B(_253_), .C(_258_), .Y(_17__2_) );
INVX1 INVX1_49 ( .A(_17__2_), .Y(_263_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_264_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_265_) );
NAND3X1 NAND3X1_24 ( .A(_263_), .B(_265_), .C(_264_), .Y(_266_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_260_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_261_) );
OAI21X1 OAI21X1_52 ( .A(_260_), .B(_261_), .C(_17__2_), .Y(_262_) );
NAND2X1 NAND2X1_58 ( .A(_262_), .B(_266_), .Y(_0__26_) );
OAI21X1 OAI21X1_53 ( .A(_263_), .B(_260_), .C(_265_), .Y(_17__3_) );
INVX1 INVX1_50 ( .A(i_add_term1[24]), .Y(_267_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[24]), .B(_267_), .Y(_268_) );
INVX1 INVX1_51 ( .A(i_add_term2[24]), .Y(_269_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term1[24]), .B(_269_), .Y(_270_) );
INVX1 INVX1_52 ( .A(i_add_term1[25]), .Y(_271_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[25]), .B(_271_), .Y(_272_) );
INVX1 INVX1_53 ( .A(i_add_term2[25]), .Y(_273_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term1[25]), .B(_273_), .Y(_274_) );
OAI22X1 OAI22X1_6 ( .A(_268_), .B(_270_), .C(_272_), .D(_274_), .Y(_275_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_276_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_277_) );
NOR2X1 NOR2X1_65 ( .A(_276_), .B(_277_), .Y(_278_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_279_) );
NAND2X1 NAND2X1_59 ( .A(_278_), .B(_279_), .Y(_280_) );
NOR2X1 NOR2X1_66 ( .A(_275_), .B(_280_), .Y(_18_) );
INVX1 INVX1_54 ( .A(_16_), .Y(_281_) );
NAND2X1 NAND2X1_60 ( .A(gnd), .B(_18_), .Y(_282_) );
OAI21X1 OAI21X1_54 ( .A(_18_), .B(_281_), .C(_282_), .Y(w_cout_6_) );
INVX1 INVX1_55 ( .A(gnd), .Y(_286_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_287_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_288_) );
NAND3X1 NAND3X1_25 ( .A(_286_), .B(_288_), .C(_287_), .Y(_289_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_283_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_284_) );
OAI21X1 OAI21X1_55 ( .A(_283_), .B(_284_), .C(gnd), .Y(_285_) );
NAND2X1 NAND2X1_62 ( .A(_285_), .B(_289_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_56 ( .A(_286_), .B(_283_), .C(_288_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_56 ( .A(rca_inst_fa3_i_carry), .Y(_293_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_294_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_295_) );
NAND3X1 NAND3X1_26 ( .A(_293_), .B(_295_), .C(_294_), .Y(_296_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_290_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_291_) );
OAI21X1 OAI21X1_57 ( .A(_290_), .B(_291_), .C(rca_inst_fa3_i_carry), .Y(_292_) );
NAND2X1 NAND2X1_64 ( .A(_292_), .B(_296_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_58 ( .A(_293_), .B(_290_), .C(_295_), .Y(cout0) );
INVX1 INVX1_57 ( .A(rca_inst_fa0_o_carry), .Y(_300_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_301_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_302_) );
NAND3X1 NAND3X1_27 ( .A(_300_), .B(_302_), .C(_301_), .Y(_303_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_297_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_298_) );
OAI21X1 OAI21X1_59 ( .A(_297_), .B(_298_), .C(rca_inst_fa0_o_carry), .Y(_299_) );
NAND2X1 NAND2X1_66 ( .A(_299_), .B(_303_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_60 ( .A(_300_), .B(_297_), .C(_302_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_58 ( .A(rca_inst_fa_1__o_carry), .Y(_307_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_308_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_309_) );
NAND3X1 NAND3X1_28 ( .A(_307_), .B(_309_), .C(_308_), .Y(_310_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_304_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_305_) );
OAI21X1 OAI21X1_61 ( .A(_304_), .B(_305_), .C(rca_inst_fa_1__o_carry), .Y(_306_) );
NAND2X1 NAND2X1_68 ( .A(_306_), .B(_310_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_62 ( .A(_307_), .B(_304_), .C(_309_), .Y(rca_inst_fa3_i_carry) );
INVX1 INVX1_59 ( .A(i_add_term1[0]), .Y(_311_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[0]), .B(_311_), .Y(_312_) );
INVX1 INVX1_60 ( .A(i_add_term2[0]), .Y(_313_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term1[0]), .B(_313_), .Y(_314_) );
INVX1 INVX1_61 ( .A(i_add_term1[1]), .Y(_315_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[1]), .B(_315_), .Y(_316_) );
INVX1 INVX1_62 ( .A(i_add_term2[1]), .Y(_317_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term1[1]), .B(_317_), .Y(_318_) );
OAI22X1 OAI22X1_7 ( .A(_312_), .B(_314_), .C(_316_), .D(_318_), .Y(_319_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_320_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_321_) );
NOR2X1 NOR2X1_76 ( .A(_320_), .B(_321_), .Y(_322_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_323_) );
NAND2X1 NAND2X1_69 ( .A(_322_), .B(_323_), .Y(_324_) );
NOR2X1 NOR2X1_77 ( .A(_319_), .B(_324_), .Y(skip0_P) );
INVX1 INVX1_63 ( .A(cout0), .Y(_325_) );
NAND2X1 NAND2X1_70 ( .A(gnd), .B(skip0_P), .Y(_326_) );
OAI21X1 OAI21X1_63 ( .A(skip0_P), .B(_325_), .C(_326_), .Y(skip0_cin_next) );
BUFX2 BUFX2_30 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_31 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_32 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_33 ( .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_34 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
