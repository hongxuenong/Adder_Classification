module csa_60bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term1[45], i_add_term1[46], i_add_term1[47], i_add_term1[48], i_add_term1[49], i_add_term1[50], i_add_term1[51], i_add_term1[52], i_add_term1[53], i_add_term1[54], i_add_term1[55], i_add_term1[56], i_add_term1[57], i_add_term1[58], i_add_term1[59], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], i_add_term2[45], i_add_term2[46], i_add_term2[47], i_add_term2[48], i_add_term2[49], i_add_term2[50], i_add_term2[51], i_add_term2[52], i_add_term2[53], i_add_term2[54], i_add_term2[55], i_add_term2[56], i_add_term2[57], i_add_term2[58], i_add_term2[59], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], sum[45], sum[46], sum[47], sum[48], sum[49], sum[50], sum[51], sum[52], sum[53], sum[54], sum[55], sum[56], sum[57], sum[58], sum[59], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term1[45];
input i_add_term1[46];
input i_add_term1[47];
input i_add_term1[48];
input i_add_term1[49];
input i_add_term1[50];
input i_add_term1[51];
input i_add_term1[52];
input i_add_term1[53];
input i_add_term1[54];
input i_add_term1[55];
input i_add_term1[56];
input i_add_term1[57];
input i_add_term1[58];
input i_add_term1[59];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
input i_add_term2[45];
input i_add_term2[46];
input i_add_term2[47];
input i_add_term2[48];
input i_add_term2[49];
input i_add_term2[50];
input i_add_term2[51];
input i_add_term2[52];
input i_add_term2[53];
input i_add_term2[54];
input i_add_term2[55];
input i_add_term2[56];
input i_add_term2[57];
input i_add_term2[58];
input i_add_term2[59];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output sum[45];
output sum[46];
output sum[47];
output sum[48];
output sum[49];
output sum[50];
output sum[51];
output sum[52];
output sum[53];
output sum[54];
output sum[55];
output sum[56];
output sum[57];
output sum[58];
output sum[59];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_14_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .A(_0__54_), .Y(sum[54]) );
BUFX2 BUFX2_57 ( .A(_0__55_), .Y(sum[55]) );
BUFX2 BUFX2_58 ( .A(_0__56_), .Y(sum[56]) );
BUFX2 BUFX2_59 ( .A(_0__57_), .Y(sum[57]) );
BUFX2 BUFX2_60 ( .A(_0__58_), .Y(sum[58]) );
BUFX2 BUFX2_61 ( .A(_0__59_), .Y(sum[59]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_85_) );
NAND2X1 NAND2X1_1 ( .A(_2_), .B(rca_inst_cout), .Y(_86_) );
OAI21X1 OAI21X1_1 ( .A(rca_inst_cout), .B(_85_), .C(_86_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3__0_), .Y(_87_) );
NAND2X1 NAND2X1_2 ( .A(_4__0_), .B(rca_inst_cout), .Y(_88_) );
OAI21X1 OAI21X1_2 ( .A(rca_inst_cout), .B(_87_), .C(_88_), .Y(_0__4_) );
INVX1 INVX1_3 ( .A(_3__1_), .Y(_89_) );
NAND2X1 NAND2X1_3 ( .A(rca_inst_cout), .B(_4__1_), .Y(_90_) );
OAI21X1 OAI21X1_3 ( .A(rca_inst_cout), .B(_89_), .C(_90_), .Y(_0__5_) );
INVX1 INVX1_4 ( .A(_3__2_), .Y(_91_) );
NAND2X1 NAND2X1_4 ( .A(rca_inst_cout), .B(_4__2_), .Y(_92_) );
OAI21X1 OAI21X1_4 ( .A(rca_inst_cout), .B(_91_), .C(_92_), .Y(_0__6_) );
INVX1 INVX1_5 ( .A(_3__3_), .Y(_93_) );
NAND2X1 NAND2X1_5 ( .A(rca_inst_cout), .B(_4__3_), .Y(_94_) );
OAI21X1 OAI21X1_5 ( .A(rca_inst_cout), .B(_93_), .C(_94_), .Y(_0__7_) );
INVX1 INVX1_6 ( .A(_7_), .Y(_95_) );
NAND2X1 NAND2X1_6 ( .A(_8_), .B(w_cout_1_), .Y(_96_) );
OAI21X1 OAI21X1_6 ( .A(w_cout_1_), .B(_95_), .C(_96_), .Y(w_cout_2_) );
INVX1 INVX1_7 ( .A(_9__0_), .Y(_97_) );
NAND2X1 NAND2X1_7 ( .A(_10__0_), .B(w_cout_1_), .Y(_98_) );
OAI21X1 OAI21X1_7 ( .A(w_cout_1_), .B(_97_), .C(_98_), .Y(_0__8_) );
INVX1 INVX1_8 ( .A(_9__1_), .Y(_99_) );
NAND2X1 NAND2X1_8 ( .A(w_cout_1_), .B(_10__1_), .Y(_100_) );
OAI21X1 OAI21X1_8 ( .A(w_cout_1_), .B(_99_), .C(_100_), .Y(_0__9_) );
INVX1 INVX1_9 ( .A(_9__2_), .Y(_101_) );
NAND2X1 NAND2X1_9 ( .A(w_cout_1_), .B(_10__2_), .Y(_102_) );
OAI21X1 OAI21X1_9 ( .A(w_cout_1_), .B(_101_), .C(_102_), .Y(_0__10_) );
INVX1 INVX1_10 ( .A(_9__3_), .Y(_103_) );
NAND2X1 NAND2X1_10 ( .A(w_cout_1_), .B(_10__3_), .Y(_104_) );
OAI21X1 OAI21X1_10 ( .A(w_cout_1_), .B(_103_), .C(_104_), .Y(_0__11_) );
INVX1 INVX1_11 ( .A(_13_), .Y(_105_) );
NAND2X1 NAND2X1_11 ( .A(_14_), .B(w_cout_2_), .Y(_106_) );
OAI21X1 OAI21X1_11 ( .A(w_cout_2_), .B(_105_), .C(_106_), .Y(w_cout_3_) );
INVX1 INVX1_12 ( .A(_15__0_), .Y(_107_) );
NAND2X1 NAND2X1_12 ( .A(_16__0_), .B(w_cout_2_), .Y(_108_) );
OAI21X1 OAI21X1_12 ( .A(w_cout_2_), .B(_107_), .C(_108_), .Y(_0__12_) );
INVX1 INVX1_13 ( .A(_15__1_), .Y(_109_) );
NAND2X1 NAND2X1_13 ( .A(w_cout_2_), .B(_16__1_), .Y(_110_) );
OAI21X1 OAI21X1_13 ( .A(w_cout_2_), .B(_109_), .C(_110_), .Y(_0__13_) );
INVX1 INVX1_14 ( .A(_15__2_), .Y(_111_) );
NAND2X1 NAND2X1_14 ( .A(w_cout_2_), .B(_16__2_), .Y(_112_) );
OAI21X1 OAI21X1_14 ( .A(w_cout_2_), .B(_111_), .C(_112_), .Y(_0__14_) );
INVX1 INVX1_15 ( .A(_15__3_), .Y(_113_) );
NAND2X1 NAND2X1_15 ( .A(w_cout_2_), .B(_16__3_), .Y(_114_) );
OAI21X1 OAI21X1_15 ( .A(w_cout_2_), .B(_113_), .C(_114_), .Y(_0__15_) );
INVX1 INVX1_16 ( .A(_19_), .Y(_115_) );
NAND2X1 NAND2X1_16 ( .A(_20_), .B(w_cout_3_), .Y(_116_) );
OAI21X1 OAI21X1_16 ( .A(w_cout_3_), .B(_115_), .C(_116_), .Y(w_cout_4_) );
INVX1 INVX1_17 ( .A(_21__0_), .Y(_117_) );
NAND2X1 NAND2X1_17 ( .A(_22__0_), .B(w_cout_3_), .Y(_118_) );
OAI21X1 OAI21X1_17 ( .A(w_cout_3_), .B(_117_), .C(_118_), .Y(_0__16_) );
INVX1 INVX1_18 ( .A(_21__1_), .Y(_119_) );
NAND2X1 NAND2X1_18 ( .A(w_cout_3_), .B(_22__1_), .Y(_120_) );
OAI21X1 OAI21X1_18 ( .A(w_cout_3_), .B(_119_), .C(_120_), .Y(_0__17_) );
INVX1 INVX1_19 ( .A(_21__2_), .Y(_121_) );
NAND2X1 NAND2X1_19 ( .A(w_cout_3_), .B(_22__2_), .Y(_122_) );
OAI21X1 OAI21X1_19 ( .A(w_cout_3_), .B(_121_), .C(_122_), .Y(_0__18_) );
INVX1 INVX1_20 ( .A(_21__3_), .Y(_123_) );
NAND2X1 NAND2X1_20 ( .A(w_cout_3_), .B(_22__3_), .Y(_124_) );
OAI21X1 OAI21X1_20 ( .A(w_cout_3_), .B(_123_), .C(_124_), .Y(_0__19_) );
INVX1 INVX1_21 ( .A(_25_), .Y(_125_) );
NAND2X1 NAND2X1_21 ( .A(_26_), .B(w_cout_4_), .Y(_126_) );
OAI21X1 OAI21X1_21 ( .A(w_cout_4_), .B(_125_), .C(_126_), .Y(w_cout_5_) );
INVX1 INVX1_22 ( .A(_27__0_), .Y(_127_) );
NAND2X1 NAND2X1_22 ( .A(_28__0_), .B(w_cout_4_), .Y(_128_) );
OAI21X1 OAI21X1_22 ( .A(w_cout_4_), .B(_127_), .C(_128_), .Y(_0__20_) );
INVX1 INVX1_23 ( .A(_27__1_), .Y(_129_) );
NAND2X1 NAND2X1_23 ( .A(w_cout_4_), .B(_28__1_), .Y(_130_) );
OAI21X1 OAI21X1_23 ( .A(w_cout_4_), .B(_129_), .C(_130_), .Y(_0__21_) );
INVX1 INVX1_24 ( .A(_27__2_), .Y(_131_) );
NAND2X1 NAND2X1_24 ( .A(w_cout_4_), .B(_28__2_), .Y(_132_) );
OAI21X1 OAI21X1_24 ( .A(w_cout_4_), .B(_131_), .C(_132_), .Y(_0__22_) );
INVX1 INVX1_25 ( .A(_27__3_), .Y(_133_) );
NAND2X1 NAND2X1_25 ( .A(w_cout_4_), .B(_28__3_), .Y(_134_) );
OAI21X1 OAI21X1_25 ( .A(w_cout_4_), .B(_133_), .C(_134_), .Y(_0__23_) );
INVX1 INVX1_26 ( .A(_31_), .Y(_135_) );
NAND2X1 NAND2X1_26 ( .A(_32_), .B(w_cout_5_), .Y(_136_) );
OAI21X1 OAI21X1_26 ( .A(w_cout_5_), .B(_135_), .C(_136_), .Y(w_cout_6_) );
INVX1 INVX1_27 ( .A(_33__0_), .Y(_137_) );
NAND2X1 NAND2X1_27 ( .A(_34__0_), .B(w_cout_5_), .Y(_138_) );
OAI21X1 OAI21X1_27 ( .A(w_cout_5_), .B(_137_), .C(_138_), .Y(_0__24_) );
INVX1 INVX1_28 ( .A(_33__1_), .Y(_139_) );
NAND2X1 NAND2X1_28 ( .A(w_cout_5_), .B(_34__1_), .Y(_140_) );
OAI21X1 OAI21X1_28 ( .A(w_cout_5_), .B(_139_), .C(_140_), .Y(_0__25_) );
INVX1 INVX1_29 ( .A(_33__2_), .Y(_141_) );
NAND2X1 NAND2X1_29 ( .A(w_cout_5_), .B(_34__2_), .Y(_142_) );
OAI21X1 OAI21X1_29 ( .A(w_cout_5_), .B(_141_), .C(_142_), .Y(_0__26_) );
INVX1 INVX1_30 ( .A(_33__3_), .Y(_143_) );
NAND2X1 NAND2X1_30 ( .A(w_cout_5_), .B(_34__3_), .Y(_144_) );
OAI21X1 OAI21X1_30 ( .A(w_cout_5_), .B(_143_), .C(_144_), .Y(_0__27_) );
INVX1 INVX1_31 ( .A(_37_), .Y(_145_) );
NAND2X1 NAND2X1_31 ( .A(_38_), .B(w_cout_6_), .Y(_146_) );
OAI21X1 OAI21X1_31 ( .A(w_cout_6_), .B(_145_), .C(_146_), .Y(w_cout_7_) );
INVX1 INVX1_32 ( .A(_39__0_), .Y(_147_) );
NAND2X1 NAND2X1_32 ( .A(_40__0_), .B(w_cout_6_), .Y(_148_) );
OAI21X1 OAI21X1_32 ( .A(w_cout_6_), .B(_147_), .C(_148_), .Y(_0__28_) );
INVX1 INVX1_33 ( .A(_39__1_), .Y(_149_) );
NAND2X1 NAND2X1_33 ( .A(w_cout_6_), .B(_40__1_), .Y(_150_) );
OAI21X1 OAI21X1_33 ( .A(w_cout_6_), .B(_149_), .C(_150_), .Y(_0__29_) );
INVX1 INVX1_34 ( .A(_39__2_), .Y(_151_) );
NAND2X1 NAND2X1_34 ( .A(w_cout_6_), .B(_40__2_), .Y(_152_) );
OAI21X1 OAI21X1_34 ( .A(w_cout_6_), .B(_151_), .C(_152_), .Y(_0__30_) );
INVX1 INVX1_35 ( .A(_39__3_), .Y(_153_) );
NAND2X1 NAND2X1_35 ( .A(w_cout_6_), .B(_40__3_), .Y(_154_) );
OAI21X1 OAI21X1_35 ( .A(w_cout_6_), .B(_153_), .C(_154_), .Y(_0__31_) );
INVX1 INVX1_36 ( .A(_43_), .Y(_155_) );
NAND2X1 NAND2X1_36 ( .A(_44_), .B(w_cout_7_), .Y(_156_) );
OAI21X1 OAI21X1_36 ( .A(w_cout_7_), .B(_155_), .C(_156_), .Y(w_cout_8_) );
INVX1 INVX1_37 ( .A(_45__0_), .Y(_157_) );
NAND2X1 NAND2X1_37 ( .A(_46__0_), .B(w_cout_7_), .Y(_158_) );
OAI21X1 OAI21X1_37 ( .A(w_cout_7_), .B(_157_), .C(_158_), .Y(_0__32_) );
INVX1 INVX1_38 ( .A(_45__1_), .Y(_159_) );
NAND2X1 NAND2X1_38 ( .A(w_cout_7_), .B(_46__1_), .Y(_160_) );
OAI21X1 OAI21X1_38 ( .A(w_cout_7_), .B(_159_), .C(_160_), .Y(_0__33_) );
INVX1 INVX1_39 ( .A(_45__2_), .Y(_161_) );
NAND2X1 NAND2X1_39 ( .A(w_cout_7_), .B(_46__2_), .Y(_162_) );
OAI21X1 OAI21X1_39 ( .A(w_cout_7_), .B(_161_), .C(_162_), .Y(_0__34_) );
INVX1 INVX1_40 ( .A(_45__3_), .Y(_163_) );
NAND2X1 NAND2X1_40 ( .A(w_cout_7_), .B(_46__3_), .Y(_164_) );
OAI21X1 OAI21X1_40 ( .A(w_cout_7_), .B(_163_), .C(_164_), .Y(_0__35_) );
INVX1 INVX1_41 ( .A(_49_), .Y(_165_) );
NAND2X1 NAND2X1_41 ( .A(_50_), .B(w_cout_8_), .Y(_166_) );
OAI21X1 OAI21X1_41 ( .A(w_cout_8_), .B(_165_), .C(_166_), .Y(w_cout_9_) );
INVX1 INVX1_42 ( .A(_51__0_), .Y(_167_) );
NAND2X1 NAND2X1_42 ( .A(_52__0_), .B(w_cout_8_), .Y(_168_) );
OAI21X1 OAI21X1_42 ( .A(w_cout_8_), .B(_167_), .C(_168_), .Y(_0__36_) );
INVX1 INVX1_43 ( .A(_51__1_), .Y(_169_) );
NAND2X1 NAND2X1_43 ( .A(w_cout_8_), .B(_52__1_), .Y(_170_) );
OAI21X1 OAI21X1_43 ( .A(w_cout_8_), .B(_169_), .C(_170_), .Y(_0__37_) );
INVX1 INVX1_44 ( .A(_51__2_), .Y(_171_) );
NAND2X1 NAND2X1_44 ( .A(w_cout_8_), .B(_52__2_), .Y(_172_) );
OAI21X1 OAI21X1_44 ( .A(w_cout_8_), .B(_171_), .C(_172_), .Y(_0__38_) );
INVX1 INVX1_45 ( .A(_51__3_), .Y(_173_) );
NAND2X1 NAND2X1_45 ( .A(w_cout_8_), .B(_52__3_), .Y(_174_) );
OAI21X1 OAI21X1_45 ( .A(w_cout_8_), .B(_173_), .C(_174_), .Y(_0__39_) );
INVX1 INVX1_46 ( .A(_55_), .Y(_175_) );
NAND2X1 NAND2X1_46 ( .A(_56_), .B(w_cout_9_), .Y(_176_) );
OAI21X1 OAI21X1_46 ( .A(w_cout_9_), .B(_175_), .C(_176_), .Y(w_cout_10_) );
INVX1 INVX1_47 ( .A(_57__0_), .Y(_177_) );
NAND2X1 NAND2X1_47 ( .A(_58__0_), .B(w_cout_9_), .Y(_178_) );
OAI21X1 OAI21X1_47 ( .A(w_cout_9_), .B(_177_), .C(_178_), .Y(_0__40_) );
INVX1 INVX1_48 ( .A(_57__1_), .Y(_179_) );
NAND2X1 NAND2X1_48 ( .A(w_cout_9_), .B(_58__1_), .Y(_180_) );
OAI21X1 OAI21X1_48 ( .A(w_cout_9_), .B(_179_), .C(_180_), .Y(_0__41_) );
INVX1 INVX1_49 ( .A(_57__2_), .Y(_181_) );
NAND2X1 NAND2X1_49 ( .A(w_cout_9_), .B(_58__2_), .Y(_182_) );
OAI21X1 OAI21X1_49 ( .A(w_cout_9_), .B(_181_), .C(_182_), .Y(_0__42_) );
INVX1 INVX1_50 ( .A(_57__3_), .Y(_183_) );
NAND2X1 NAND2X1_50 ( .A(w_cout_9_), .B(_58__3_), .Y(_184_) );
OAI21X1 OAI21X1_50 ( .A(w_cout_9_), .B(_183_), .C(_184_), .Y(_0__43_) );
INVX1 INVX1_51 ( .A(_61_), .Y(_185_) );
NAND2X1 NAND2X1_51 ( .A(_62_), .B(w_cout_10_), .Y(_186_) );
OAI21X1 OAI21X1_51 ( .A(w_cout_10_), .B(_185_), .C(_186_), .Y(w_cout_11_) );
INVX1 INVX1_52 ( .A(_63__0_), .Y(_187_) );
NAND2X1 NAND2X1_52 ( .A(_64__0_), .B(w_cout_10_), .Y(_188_) );
OAI21X1 OAI21X1_52 ( .A(w_cout_10_), .B(_187_), .C(_188_), .Y(_0__44_) );
INVX1 INVX1_53 ( .A(_63__1_), .Y(_189_) );
NAND2X1 NAND2X1_53 ( .A(w_cout_10_), .B(_64__1_), .Y(_190_) );
OAI21X1 OAI21X1_53 ( .A(w_cout_10_), .B(_189_), .C(_190_), .Y(_0__45_) );
INVX1 INVX1_54 ( .A(_63__2_), .Y(_191_) );
NAND2X1 NAND2X1_54 ( .A(w_cout_10_), .B(_64__2_), .Y(_192_) );
OAI21X1 OAI21X1_54 ( .A(w_cout_10_), .B(_191_), .C(_192_), .Y(_0__46_) );
INVX1 INVX1_55 ( .A(_63__3_), .Y(_193_) );
NAND2X1 NAND2X1_55 ( .A(w_cout_10_), .B(_64__3_), .Y(_194_) );
OAI21X1 OAI21X1_55 ( .A(w_cout_10_), .B(_193_), .C(_194_), .Y(_0__47_) );
INVX1 INVX1_56 ( .A(_67_), .Y(_195_) );
NAND2X1 NAND2X1_56 ( .A(_68_), .B(w_cout_11_), .Y(_196_) );
OAI21X1 OAI21X1_56 ( .A(w_cout_11_), .B(_195_), .C(_196_), .Y(w_cout_12_) );
INVX1 INVX1_57 ( .A(_69__0_), .Y(_197_) );
NAND2X1 NAND2X1_57 ( .A(_70__0_), .B(w_cout_11_), .Y(_198_) );
OAI21X1 OAI21X1_57 ( .A(w_cout_11_), .B(_197_), .C(_198_), .Y(_0__48_) );
INVX1 INVX1_58 ( .A(_69__1_), .Y(_199_) );
NAND2X1 NAND2X1_58 ( .A(w_cout_11_), .B(_70__1_), .Y(_200_) );
OAI21X1 OAI21X1_58 ( .A(w_cout_11_), .B(_199_), .C(_200_), .Y(_0__49_) );
INVX1 INVX1_59 ( .A(_69__2_), .Y(_201_) );
NAND2X1 NAND2X1_59 ( .A(w_cout_11_), .B(_70__2_), .Y(_202_) );
OAI21X1 OAI21X1_59 ( .A(w_cout_11_), .B(_201_), .C(_202_), .Y(_0__50_) );
INVX1 INVX1_60 ( .A(_69__3_), .Y(_203_) );
NAND2X1 NAND2X1_60 ( .A(w_cout_11_), .B(_70__3_), .Y(_204_) );
OAI21X1 OAI21X1_60 ( .A(w_cout_11_), .B(_203_), .C(_204_), .Y(_0__51_) );
INVX1 INVX1_61 ( .A(_73_), .Y(_205_) );
NAND2X1 NAND2X1_61 ( .A(_74_), .B(w_cout_12_), .Y(_206_) );
OAI21X1 OAI21X1_61 ( .A(w_cout_12_), .B(_205_), .C(_206_), .Y(w_cout_13_) );
INVX1 INVX1_62 ( .A(_75__0_), .Y(_207_) );
NAND2X1 NAND2X1_62 ( .A(_76__0_), .B(w_cout_12_), .Y(_208_) );
OAI21X1 OAI21X1_62 ( .A(w_cout_12_), .B(_207_), .C(_208_), .Y(_0__52_) );
INVX1 INVX1_63 ( .A(_75__1_), .Y(_209_) );
NAND2X1 NAND2X1_63 ( .A(w_cout_12_), .B(_76__1_), .Y(_210_) );
OAI21X1 OAI21X1_63 ( .A(w_cout_12_), .B(_209_), .C(_210_), .Y(_0__53_) );
INVX1 INVX1_64 ( .A(_75__2_), .Y(_211_) );
NAND2X1 NAND2X1_64 ( .A(w_cout_12_), .B(_76__2_), .Y(_212_) );
OAI21X1 OAI21X1_64 ( .A(w_cout_12_), .B(_211_), .C(_212_), .Y(_0__54_) );
INVX1 INVX1_65 ( .A(_75__3_), .Y(_213_) );
NAND2X1 NAND2X1_65 ( .A(w_cout_12_), .B(_76__3_), .Y(_214_) );
OAI21X1 OAI21X1_65 ( .A(w_cout_12_), .B(_213_), .C(_214_), .Y(_0__55_) );
INVX1 INVX1_66 ( .A(_79_), .Y(_215_) );
NAND2X1 NAND2X1_66 ( .A(_80_), .B(w_cout_13_), .Y(_216_) );
OAI21X1 OAI21X1_66 ( .A(w_cout_13_), .B(_215_), .C(_216_), .Y(w_cout_14_) );
INVX1 INVX1_67 ( .A(_81__0_), .Y(_217_) );
NAND2X1 NAND2X1_67 ( .A(_82__0_), .B(w_cout_13_), .Y(_218_) );
OAI21X1 OAI21X1_67 ( .A(w_cout_13_), .B(_217_), .C(_218_), .Y(_0__56_) );
INVX1 INVX1_68 ( .A(_81__1_), .Y(_219_) );
NAND2X1 NAND2X1_68 ( .A(w_cout_13_), .B(_82__1_), .Y(_220_) );
OAI21X1 OAI21X1_68 ( .A(w_cout_13_), .B(_219_), .C(_220_), .Y(_0__57_) );
INVX1 INVX1_69 ( .A(_81__2_), .Y(_221_) );
NAND2X1 NAND2X1_69 ( .A(w_cout_13_), .B(_82__2_), .Y(_222_) );
OAI21X1 OAI21X1_69 ( .A(w_cout_13_), .B(_221_), .C(_222_), .Y(_0__58_) );
INVX1 INVX1_70 ( .A(_81__3_), .Y(_223_) );
NAND2X1 NAND2X1_70 ( .A(w_cout_13_), .B(_82__3_), .Y(_224_) );
OAI21X1 OAI21X1_70 ( .A(w_cout_13_), .B(_223_), .C(_224_), .Y(_0__59_) );
INVX1 INVX1_71 ( .A(1'b0), .Y(_228_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_229_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_230_) );
NAND3X1 NAND3X1_1 ( .A(_228_), .B(_230_), .C(_229_), .Y(_231_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_225_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_226_) );
OAI21X1 OAI21X1_71 ( .A(_225_), .B(_226_), .C(1'b0), .Y(_227_) );
NAND2X1 NAND2X1_72 ( .A(_227_), .B(_231_), .Y(_3__0_) );
OAI21X1 OAI21X1_72 ( .A(_228_), .B(_225_), .C(_230_), .Y(_5__1_) );
INVX1 INVX1_72 ( .A(_5__1_), .Y(_235_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_236_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_237_) );
NAND3X1 NAND3X1_2 ( .A(_235_), .B(_237_), .C(_236_), .Y(_238_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_232_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_233_) );
OAI21X1 OAI21X1_73 ( .A(_232_), .B(_233_), .C(_5__1_), .Y(_234_) );
NAND2X1 NAND2X1_74 ( .A(_234_), .B(_238_), .Y(_3__1_) );
OAI21X1 OAI21X1_74 ( .A(_235_), .B(_232_), .C(_237_), .Y(_5__2_) );
INVX1 INVX1_73 ( .A(_5__2_), .Y(_242_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_243_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_244_) );
NAND3X1 NAND3X1_3 ( .A(_242_), .B(_244_), .C(_243_), .Y(_245_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_239_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_240_) );
OAI21X1 OAI21X1_75 ( .A(_239_), .B(_240_), .C(_5__2_), .Y(_241_) );
NAND2X1 NAND2X1_76 ( .A(_241_), .B(_245_), .Y(_3__2_) );
OAI21X1 OAI21X1_76 ( .A(_242_), .B(_239_), .C(_244_), .Y(_5__3_) );
INVX1 INVX1_74 ( .A(_5__3_), .Y(_249_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_250_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_251_) );
NAND3X1 NAND3X1_4 ( .A(_249_), .B(_251_), .C(_250_), .Y(_252_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_246_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_247_) );
OAI21X1 OAI21X1_77 ( .A(_246_), .B(_247_), .C(_5__3_), .Y(_248_) );
NAND2X1 NAND2X1_78 ( .A(_248_), .B(_252_), .Y(_3__3_) );
OAI21X1 OAI21X1_78 ( .A(_249_), .B(_246_), .C(_251_), .Y(_1_) );
INVX1 INVX1_75 ( .A(1'b1), .Y(_256_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_257_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_258_) );
NAND3X1 NAND3X1_5 ( .A(_256_), .B(_258_), .C(_257_), .Y(_259_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_253_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_254_) );
OAI21X1 OAI21X1_79 ( .A(_253_), .B(_254_), .C(1'b1), .Y(_255_) );
NAND2X1 NAND2X1_80 ( .A(_255_), .B(_259_), .Y(_4__0_) );
OAI21X1 OAI21X1_80 ( .A(_256_), .B(_253_), .C(_258_), .Y(_6__1_) );
INVX1 INVX1_76 ( .A(_6__1_), .Y(_263_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_264_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_265_) );
NAND3X1 NAND3X1_6 ( .A(_263_), .B(_265_), .C(_264_), .Y(_266_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_260_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_261_) );
OAI21X1 OAI21X1_81 ( .A(_260_), .B(_261_), .C(_6__1_), .Y(_262_) );
NAND2X1 NAND2X1_82 ( .A(_262_), .B(_266_), .Y(_4__1_) );
OAI21X1 OAI21X1_82 ( .A(_263_), .B(_260_), .C(_265_), .Y(_6__2_) );
INVX1 INVX1_77 ( .A(_6__2_), .Y(_270_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_271_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_272_) );
NAND3X1 NAND3X1_7 ( .A(_270_), .B(_272_), .C(_271_), .Y(_273_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_267_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_268_) );
OAI21X1 OAI21X1_83 ( .A(_267_), .B(_268_), .C(_6__2_), .Y(_269_) );
NAND2X1 NAND2X1_84 ( .A(_269_), .B(_273_), .Y(_4__2_) );
OAI21X1 OAI21X1_84 ( .A(_270_), .B(_267_), .C(_272_), .Y(_6__3_) );
INVX1 INVX1_78 ( .A(_6__3_), .Y(_277_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_278_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_279_) );
NAND3X1 NAND3X1_8 ( .A(_277_), .B(_279_), .C(_278_), .Y(_280_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_274_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_275_) );
OAI21X1 OAI21X1_85 ( .A(_274_), .B(_275_), .C(_6__3_), .Y(_276_) );
NAND2X1 NAND2X1_86 ( .A(_276_), .B(_280_), .Y(_4__3_) );
OAI21X1 OAI21X1_86 ( .A(_277_), .B(_274_), .C(_279_), .Y(_2_) );
INVX1 INVX1_79 ( .A(1'b0), .Y(_284_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_285_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_286_) );
NAND3X1 NAND3X1_9 ( .A(_284_), .B(_286_), .C(_285_), .Y(_287_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_281_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_282_) );
OAI21X1 OAI21X1_87 ( .A(_281_), .B(_282_), .C(1'b0), .Y(_283_) );
NAND2X1 NAND2X1_88 ( .A(_283_), .B(_287_), .Y(_9__0_) );
OAI21X1 OAI21X1_88 ( .A(_284_), .B(_281_), .C(_286_), .Y(_11__1_) );
INVX1 INVX1_80 ( .A(_11__1_), .Y(_291_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_292_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_293_) );
NAND3X1 NAND3X1_10 ( .A(_291_), .B(_293_), .C(_292_), .Y(_294_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_288_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_289_) );
OAI21X1 OAI21X1_89 ( .A(_288_), .B(_289_), .C(_11__1_), .Y(_290_) );
NAND2X1 NAND2X1_90 ( .A(_290_), .B(_294_), .Y(_9__1_) );
OAI21X1 OAI21X1_90 ( .A(_291_), .B(_288_), .C(_293_), .Y(_11__2_) );
INVX1 INVX1_81 ( .A(_11__2_), .Y(_298_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_299_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_300_) );
NAND3X1 NAND3X1_11 ( .A(_298_), .B(_300_), .C(_299_), .Y(_301_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_295_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_296_) );
OAI21X1 OAI21X1_91 ( .A(_295_), .B(_296_), .C(_11__2_), .Y(_297_) );
NAND2X1 NAND2X1_92 ( .A(_297_), .B(_301_), .Y(_9__2_) );
OAI21X1 OAI21X1_92 ( .A(_298_), .B(_295_), .C(_300_), .Y(_11__3_) );
INVX1 INVX1_82 ( .A(_11__3_), .Y(_305_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_306_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_307_) );
NAND3X1 NAND3X1_12 ( .A(_305_), .B(_307_), .C(_306_), .Y(_308_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_302_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_303_) );
OAI21X1 OAI21X1_93 ( .A(_302_), .B(_303_), .C(_11__3_), .Y(_304_) );
NAND2X1 NAND2X1_94 ( .A(_304_), .B(_308_), .Y(_9__3_) );
OAI21X1 OAI21X1_94 ( .A(_305_), .B(_302_), .C(_307_), .Y(_7_) );
INVX1 INVX1_83 ( .A(1'b1), .Y(_312_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_313_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_314_) );
NAND3X1 NAND3X1_13 ( .A(_312_), .B(_314_), .C(_313_), .Y(_315_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_309_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_310_) );
OAI21X1 OAI21X1_95 ( .A(_309_), .B(_310_), .C(1'b1), .Y(_311_) );
NAND2X1 NAND2X1_96 ( .A(_311_), .B(_315_), .Y(_10__0_) );
OAI21X1 OAI21X1_96 ( .A(_312_), .B(_309_), .C(_314_), .Y(_12__1_) );
INVX1 INVX1_84 ( .A(_12__1_), .Y(_319_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_320_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_321_) );
NAND3X1 NAND3X1_14 ( .A(_319_), .B(_321_), .C(_320_), .Y(_322_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_316_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_317_) );
OAI21X1 OAI21X1_97 ( .A(_316_), .B(_317_), .C(_12__1_), .Y(_318_) );
NAND2X1 NAND2X1_98 ( .A(_318_), .B(_322_), .Y(_10__1_) );
OAI21X1 OAI21X1_98 ( .A(_319_), .B(_316_), .C(_321_), .Y(_12__2_) );
INVX1 INVX1_85 ( .A(_12__2_), .Y(_326_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_327_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_328_) );
NAND3X1 NAND3X1_15 ( .A(_326_), .B(_328_), .C(_327_), .Y(_329_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_323_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_324_) );
OAI21X1 OAI21X1_99 ( .A(_323_), .B(_324_), .C(_12__2_), .Y(_325_) );
NAND2X1 NAND2X1_100 ( .A(_325_), .B(_329_), .Y(_10__2_) );
OAI21X1 OAI21X1_100 ( .A(_326_), .B(_323_), .C(_328_), .Y(_12__3_) );
INVX1 INVX1_86 ( .A(_12__3_), .Y(_333_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_334_) );
NAND2X1 NAND2X1_101 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_335_) );
NAND3X1 NAND3X1_16 ( .A(_333_), .B(_335_), .C(_334_), .Y(_336_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_330_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_331_) );
OAI21X1 OAI21X1_101 ( .A(_330_), .B(_331_), .C(_12__3_), .Y(_332_) );
NAND2X1 NAND2X1_102 ( .A(_332_), .B(_336_), .Y(_10__3_) );
OAI21X1 OAI21X1_102 ( .A(_333_), .B(_330_), .C(_335_), .Y(_8_) );
INVX1 INVX1_87 ( .A(1'b0), .Y(_340_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_341_) );
NAND2X1 NAND2X1_103 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_342_) );
NAND3X1 NAND3X1_17 ( .A(_340_), .B(_342_), .C(_341_), .Y(_343_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_337_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_338_) );
OAI21X1 OAI21X1_103 ( .A(_337_), .B(_338_), .C(1'b0), .Y(_339_) );
NAND2X1 NAND2X1_104 ( .A(_339_), .B(_343_), .Y(_15__0_) );
OAI21X1 OAI21X1_104 ( .A(_340_), .B(_337_), .C(_342_), .Y(_17__1_) );
INVX1 INVX1_88 ( .A(_17__1_), .Y(_347_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_348_) );
NAND2X1 NAND2X1_105 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_349_) );
NAND3X1 NAND3X1_18 ( .A(_347_), .B(_349_), .C(_348_), .Y(_350_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_344_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_345_) );
OAI21X1 OAI21X1_105 ( .A(_344_), .B(_345_), .C(_17__1_), .Y(_346_) );
NAND2X1 NAND2X1_106 ( .A(_346_), .B(_350_), .Y(_15__1_) );
OAI21X1 OAI21X1_106 ( .A(_347_), .B(_344_), .C(_349_), .Y(_17__2_) );
INVX1 INVX1_89 ( .A(_17__2_), .Y(_354_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_355_) );
NAND2X1 NAND2X1_107 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_356_) );
NAND3X1 NAND3X1_19 ( .A(_354_), .B(_356_), .C(_355_), .Y(_357_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_351_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_352_) );
OAI21X1 OAI21X1_107 ( .A(_351_), .B(_352_), .C(_17__2_), .Y(_353_) );
NAND2X1 NAND2X1_108 ( .A(_353_), .B(_357_), .Y(_15__2_) );
OAI21X1 OAI21X1_108 ( .A(_354_), .B(_351_), .C(_356_), .Y(_17__3_) );
INVX1 INVX1_90 ( .A(_17__3_), .Y(_361_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_362_) );
NAND2X1 NAND2X1_109 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_363_) );
NAND3X1 NAND3X1_20 ( .A(_361_), .B(_363_), .C(_362_), .Y(_364_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_358_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_359_) );
OAI21X1 OAI21X1_109 ( .A(_358_), .B(_359_), .C(_17__3_), .Y(_360_) );
NAND2X1 NAND2X1_110 ( .A(_360_), .B(_364_), .Y(_15__3_) );
OAI21X1 OAI21X1_110 ( .A(_361_), .B(_358_), .C(_363_), .Y(_13_) );
INVX1 INVX1_91 ( .A(1'b1), .Y(_368_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_369_) );
NAND2X1 NAND2X1_111 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_370_) );
NAND3X1 NAND3X1_21 ( .A(_368_), .B(_370_), .C(_369_), .Y(_371_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_365_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_366_) );
OAI21X1 OAI21X1_111 ( .A(_365_), .B(_366_), .C(1'b1), .Y(_367_) );
NAND2X1 NAND2X1_112 ( .A(_367_), .B(_371_), .Y(_16__0_) );
OAI21X1 OAI21X1_112 ( .A(_368_), .B(_365_), .C(_370_), .Y(_18__1_) );
INVX1 INVX1_92 ( .A(_18__1_), .Y(_375_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_376_) );
NAND2X1 NAND2X1_113 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_377_) );
NAND3X1 NAND3X1_22 ( .A(_375_), .B(_377_), .C(_376_), .Y(_378_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_372_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_373_) );
OAI21X1 OAI21X1_113 ( .A(_372_), .B(_373_), .C(_18__1_), .Y(_374_) );
NAND2X1 NAND2X1_114 ( .A(_374_), .B(_378_), .Y(_16__1_) );
OAI21X1 OAI21X1_114 ( .A(_375_), .B(_372_), .C(_377_), .Y(_18__2_) );
INVX1 INVX1_93 ( .A(_18__2_), .Y(_382_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_383_) );
NAND2X1 NAND2X1_115 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_384_) );
NAND3X1 NAND3X1_23 ( .A(_382_), .B(_384_), .C(_383_), .Y(_385_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_379_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_380_) );
OAI21X1 OAI21X1_115 ( .A(_379_), .B(_380_), .C(_18__2_), .Y(_381_) );
NAND2X1 NAND2X1_116 ( .A(_381_), .B(_385_), .Y(_16__2_) );
OAI21X1 OAI21X1_116 ( .A(_382_), .B(_379_), .C(_384_), .Y(_18__3_) );
INVX1 INVX1_94 ( .A(_18__3_), .Y(_389_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_390_) );
NAND2X1 NAND2X1_117 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_391_) );
NAND3X1 NAND3X1_24 ( .A(_389_), .B(_391_), .C(_390_), .Y(_392_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_386_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_387_) );
OAI21X1 OAI21X1_117 ( .A(_386_), .B(_387_), .C(_18__3_), .Y(_388_) );
NAND2X1 NAND2X1_118 ( .A(_388_), .B(_392_), .Y(_16__3_) );
OAI21X1 OAI21X1_118 ( .A(_389_), .B(_386_), .C(_391_), .Y(_14_) );
INVX1 INVX1_95 ( .A(1'b0), .Y(_396_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_397_) );
NAND2X1 NAND2X1_119 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_398_) );
NAND3X1 NAND3X1_25 ( .A(_396_), .B(_398_), .C(_397_), .Y(_399_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_393_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_394_) );
OAI21X1 OAI21X1_119 ( .A(_393_), .B(_394_), .C(1'b0), .Y(_395_) );
NAND2X1 NAND2X1_120 ( .A(_395_), .B(_399_), .Y(_21__0_) );
OAI21X1 OAI21X1_120 ( .A(_396_), .B(_393_), .C(_398_), .Y(_23__1_) );
INVX1 INVX1_96 ( .A(_23__1_), .Y(_403_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_404_) );
NAND2X1 NAND2X1_121 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_405_) );
NAND3X1 NAND3X1_26 ( .A(_403_), .B(_405_), .C(_404_), .Y(_406_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_400_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_401_) );
OAI21X1 OAI21X1_121 ( .A(_400_), .B(_401_), .C(_23__1_), .Y(_402_) );
NAND2X1 NAND2X1_122 ( .A(_402_), .B(_406_), .Y(_21__1_) );
OAI21X1 OAI21X1_122 ( .A(_403_), .B(_400_), .C(_405_), .Y(_23__2_) );
INVX1 INVX1_97 ( .A(_23__2_), .Y(_410_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_411_) );
NAND2X1 NAND2X1_123 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_412_) );
NAND3X1 NAND3X1_27 ( .A(_410_), .B(_412_), .C(_411_), .Y(_413_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_407_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_408_) );
OAI21X1 OAI21X1_123 ( .A(_407_), .B(_408_), .C(_23__2_), .Y(_409_) );
NAND2X1 NAND2X1_124 ( .A(_409_), .B(_413_), .Y(_21__2_) );
OAI21X1 OAI21X1_124 ( .A(_410_), .B(_407_), .C(_412_), .Y(_23__3_) );
INVX1 INVX1_98 ( .A(_23__3_), .Y(_417_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_418_) );
NAND2X1 NAND2X1_125 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_419_) );
NAND3X1 NAND3X1_28 ( .A(_417_), .B(_419_), .C(_418_), .Y(_420_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_414_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_415_) );
OAI21X1 OAI21X1_125 ( .A(_414_), .B(_415_), .C(_23__3_), .Y(_416_) );
NAND2X1 NAND2X1_126 ( .A(_416_), .B(_420_), .Y(_21__3_) );
OAI21X1 OAI21X1_126 ( .A(_417_), .B(_414_), .C(_419_), .Y(_19_) );
INVX1 INVX1_99 ( .A(1'b1), .Y(_424_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_425_) );
NAND2X1 NAND2X1_127 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_426_) );
NAND3X1 NAND3X1_29 ( .A(_424_), .B(_426_), .C(_425_), .Y(_427_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_421_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_422_) );
OAI21X1 OAI21X1_127 ( .A(_421_), .B(_422_), .C(1'b1), .Y(_423_) );
NAND2X1 NAND2X1_128 ( .A(_423_), .B(_427_), .Y(_22__0_) );
OAI21X1 OAI21X1_128 ( .A(_424_), .B(_421_), .C(_426_), .Y(_24__1_) );
INVX1 INVX1_100 ( .A(_24__1_), .Y(_431_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_432_) );
NAND2X1 NAND2X1_129 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_433_) );
NAND3X1 NAND3X1_30 ( .A(_431_), .B(_433_), .C(_432_), .Y(_434_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_428_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_429_) );
OAI21X1 OAI21X1_129 ( .A(_428_), .B(_429_), .C(_24__1_), .Y(_430_) );
NAND2X1 NAND2X1_130 ( .A(_430_), .B(_434_), .Y(_22__1_) );
OAI21X1 OAI21X1_130 ( .A(_431_), .B(_428_), .C(_433_), .Y(_24__2_) );
INVX1 INVX1_101 ( .A(_24__2_), .Y(_438_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_439_) );
NAND2X1 NAND2X1_131 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_440_) );
NAND3X1 NAND3X1_31 ( .A(_438_), .B(_440_), .C(_439_), .Y(_441_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_435_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_436_) );
OAI21X1 OAI21X1_131 ( .A(_435_), .B(_436_), .C(_24__2_), .Y(_437_) );
NAND2X1 NAND2X1_132 ( .A(_437_), .B(_441_), .Y(_22__2_) );
OAI21X1 OAI21X1_132 ( .A(_438_), .B(_435_), .C(_440_), .Y(_24__3_) );
INVX1 INVX1_102 ( .A(_24__3_), .Y(_445_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_446_) );
NAND2X1 NAND2X1_133 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_447_) );
NAND3X1 NAND3X1_32 ( .A(_445_), .B(_447_), .C(_446_), .Y(_448_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_442_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_443_) );
OAI21X1 OAI21X1_133 ( .A(_442_), .B(_443_), .C(_24__3_), .Y(_444_) );
NAND2X1 NAND2X1_134 ( .A(_444_), .B(_448_), .Y(_22__3_) );
OAI21X1 OAI21X1_134 ( .A(_445_), .B(_442_), .C(_447_), .Y(_20_) );
INVX1 INVX1_103 ( .A(1'b0), .Y(_452_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_453_) );
NAND2X1 NAND2X1_135 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_454_) );
NAND3X1 NAND3X1_33 ( .A(_452_), .B(_454_), .C(_453_), .Y(_455_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_449_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_450_) );
OAI21X1 OAI21X1_135 ( .A(_449_), .B(_450_), .C(1'b0), .Y(_451_) );
NAND2X1 NAND2X1_136 ( .A(_451_), .B(_455_), .Y(_27__0_) );
OAI21X1 OAI21X1_136 ( .A(_452_), .B(_449_), .C(_454_), .Y(_29__1_) );
INVX1 INVX1_104 ( .A(_29__1_), .Y(_459_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_460_) );
NAND2X1 NAND2X1_137 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_461_) );
NAND3X1 NAND3X1_34 ( .A(_459_), .B(_461_), .C(_460_), .Y(_462_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_456_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_457_) );
OAI21X1 OAI21X1_137 ( .A(_456_), .B(_457_), .C(_29__1_), .Y(_458_) );
NAND2X1 NAND2X1_138 ( .A(_458_), .B(_462_), .Y(_27__1_) );
OAI21X1 OAI21X1_138 ( .A(_459_), .B(_456_), .C(_461_), .Y(_29__2_) );
INVX1 INVX1_105 ( .A(_29__2_), .Y(_466_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_467_) );
NAND2X1 NAND2X1_139 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_468_) );
NAND3X1 NAND3X1_35 ( .A(_466_), .B(_468_), .C(_467_), .Y(_469_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_463_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_464_) );
OAI21X1 OAI21X1_139 ( .A(_463_), .B(_464_), .C(_29__2_), .Y(_465_) );
NAND2X1 NAND2X1_140 ( .A(_465_), .B(_469_), .Y(_27__2_) );
OAI21X1 OAI21X1_140 ( .A(_466_), .B(_463_), .C(_468_), .Y(_29__3_) );
INVX1 INVX1_106 ( .A(_29__3_), .Y(_473_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_474_) );
NAND2X1 NAND2X1_141 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_475_) );
NAND3X1 NAND3X1_36 ( .A(_473_), .B(_475_), .C(_474_), .Y(_476_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_470_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_471_) );
OAI21X1 OAI21X1_141 ( .A(_470_), .B(_471_), .C(_29__3_), .Y(_472_) );
NAND2X1 NAND2X1_142 ( .A(_472_), .B(_476_), .Y(_27__3_) );
OAI21X1 OAI21X1_142 ( .A(_473_), .B(_470_), .C(_475_), .Y(_25_) );
INVX1 INVX1_107 ( .A(1'b1), .Y(_480_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_481_) );
NAND2X1 NAND2X1_143 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_482_) );
NAND3X1 NAND3X1_37 ( .A(_480_), .B(_482_), .C(_481_), .Y(_483_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_477_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_478_) );
OAI21X1 OAI21X1_143 ( .A(_477_), .B(_478_), .C(1'b1), .Y(_479_) );
NAND2X1 NAND2X1_144 ( .A(_479_), .B(_483_), .Y(_28__0_) );
OAI21X1 OAI21X1_144 ( .A(_480_), .B(_477_), .C(_482_), .Y(_30__1_) );
INVX1 INVX1_108 ( .A(_30__1_), .Y(_487_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_488_) );
NAND2X1 NAND2X1_145 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_489_) );
NAND3X1 NAND3X1_38 ( .A(_487_), .B(_489_), .C(_488_), .Y(_490_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_484_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_485_) );
OAI21X1 OAI21X1_145 ( .A(_484_), .B(_485_), .C(_30__1_), .Y(_486_) );
NAND2X1 NAND2X1_146 ( .A(_486_), .B(_490_), .Y(_28__1_) );
OAI21X1 OAI21X1_146 ( .A(_487_), .B(_484_), .C(_489_), .Y(_30__2_) );
INVX1 INVX1_109 ( .A(_30__2_), .Y(_494_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_495_) );
NAND2X1 NAND2X1_147 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_496_) );
NAND3X1 NAND3X1_39 ( .A(_494_), .B(_496_), .C(_495_), .Y(_497_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_491_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_492_) );
OAI21X1 OAI21X1_147 ( .A(_491_), .B(_492_), .C(_30__2_), .Y(_493_) );
NAND2X1 NAND2X1_148 ( .A(_493_), .B(_497_), .Y(_28__2_) );
OAI21X1 OAI21X1_148 ( .A(_494_), .B(_491_), .C(_496_), .Y(_30__3_) );
INVX1 INVX1_110 ( .A(_30__3_), .Y(_501_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_502_) );
NAND2X1 NAND2X1_149 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_503_) );
NAND3X1 NAND3X1_40 ( .A(_501_), .B(_503_), .C(_502_), .Y(_504_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_498_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_499_) );
OAI21X1 OAI21X1_149 ( .A(_498_), .B(_499_), .C(_30__3_), .Y(_500_) );
NAND2X1 NAND2X1_150 ( .A(_500_), .B(_504_), .Y(_28__3_) );
OAI21X1 OAI21X1_150 ( .A(_501_), .B(_498_), .C(_503_), .Y(_26_) );
INVX1 INVX1_111 ( .A(1'b0), .Y(_508_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_509_) );
NAND2X1 NAND2X1_151 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_510_) );
NAND3X1 NAND3X1_41 ( .A(_508_), .B(_510_), .C(_509_), .Y(_511_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_505_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_506_) );
OAI21X1 OAI21X1_151 ( .A(_505_), .B(_506_), .C(1'b0), .Y(_507_) );
NAND2X1 NAND2X1_152 ( .A(_507_), .B(_511_), .Y(_33__0_) );
OAI21X1 OAI21X1_152 ( .A(_508_), .B(_505_), .C(_510_), .Y(_35__1_) );
INVX1 INVX1_112 ( .A(_35__1_), .Y(_515_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_516_) );
NAND2X1 NAND2X1_153 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_517_) );
NAND3X1 NAND3X1_42 ( .A(_515_), .B(_517_), .C(_516_), .Y(_518_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_512_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_513_) );
OAI21X1 OAI21X1_153 ( .A(_512_), .B(_513_), .C(_35__1_), .Y(_514_) );
NAND2X1 NAND2X1_154 ( .A(_514_), .B(_518_), .Y(_33__1_) );
OAI21X1 OAI21X1_154 ( .A(_515_), .B(_512_), .C(_517_), .Y(_35__2_) );
INVX1 INVX1_113 ( .A(_35__2_), .Y(_522_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_523_) );
NAND2X1 NAND2X1_155 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_524_) );
NAND3X1 NAND3X1_43 ( .A(_522_), .B(_524_), .C(_523_), .Y(_525_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_519_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_520_) );
OAI21X1 OAI21X1_155 ( .A(_519_), .B(_520_), .C(_35__2_), .Y(_521_) );
NAND2X1 NAND2X1_156 ( .A(_521_), .B(_525_), .Y(_33__2_) );
OAI21X1 OAI21X1_156 ( .A(_522_), .B(_519_), .C(_524_), .Y(_35__3_) );
INVX1 INVX1_114 ( .A(_35__3_), .Y(_529_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_530_) );
NAND2X1 NAND2X1_157 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_531_) );
NAND3X1 NAND3X1_44 ( .A(_529_), .B(_531_), .C(_530_), .Y(_532_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_526_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_527_) );
OAI21X1 OAI21X1_157 ( .A(_526_), .B(_527_), .C(_35__3_), .Y(_528_) );
NAND2X1 NAND2X1_158 ( .A(_528_), .B(_532_), .Y(_33__3_) );
OAI21X1 OAI21X1_158 ( .A(_529_), .B(_526_), .C(_531_), .Y(_31_) );
INVX1 INVX1_115 ( .A(1'b1), .Y(_536_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_537_) );
NAND2X1 NAND2X1_159 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_538_) );
NAND3X1 NAND3X1_45 ( .A(_536_), .B(_538_), .C(_537_), .Y(_539_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_533_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_534_) );
OAI21X1 OAI21X1_159 ( .A(_533_), .B(_534_), .C(1'b1), .Y(_535_) );
NAND2X1 NAND2X1_160 ( .A(_535_), .B(_539_), .Y(_34__0_) );
OAI21X1 OAI21X1_160 ( .A(_536_), .B(_533_), .C(_538_), .Y(_36__1_) );
INVX1 INVX1_116 ( .A(_36__1_), .Y(_543_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_544_) );
NAND2X1 NAND2X1_161 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_545_) );
NAND3X1 NAND3X1_46 ( .A(_543_), .B(_545_), .C(_544_), .Y(_546_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_540_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_541_) );
OAI21X1 OAI21X1_161 ( .A(_540_), .B(_541_), .C(_36__1_), .Y(_542_) );
NAND2X1 NAND2X1_162 ( .A(_542_), .B(_546_), .Y(_34__1_) );
OAI21X1 OAI21X1_162 ( .A(_543_), .B(_540_), .C(_545_), .Y(_36__2_) );
INVX1 INVX1_117 ( .A(_36__2_), .Y(_550_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_551_) );
NAND2X1 NAND2X1_163 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_552_) );
NAND3X1 NAND3X1_47 ( .A(_550_), .B(_552_), .C(_551_), .Y(_553_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_547_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_548_) );
OAI21X1 OAI21X1_163 ( .A(_547_), .B(_548_), .C(_36__2_), .Y(_549_) );
NAND2X1 NAND2X1_164 ( .A(_549_), .B(_553_), .Y(_34__2_) );
OAI21X1 OAI21X1_164 ( .A(_550_), .B(_547_), .C(_552_), .Y(_36__3_) );
INVX1 INVX1_118 ( .A(_36__3_), .Y(_557_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_558_) );
NAND2X1 NAND2X1_165 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_559_) );
NAND3X1 NAND3X1_48 ( .A(_557_), .B(_559_), .C(_558_), .Y(_560_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_554_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_555_) );
OAI21X1 OAI21X1_165 ( .A(_554_), .B(_555_), .C(_36__3_), .Y(_556_) );
NAND2X1 NAND2X1_166 ( .A(_556_), .B(_560_), .Y(_34__3_) );
OAI21X1 OAI21X1_166 ( .A(_557_), .B(_554_), .C(_559_), .Y(_32_) );
INVX1 INVX1_119 ( .A(1'b0), .Y(_564_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_565_) );
NAND2X1 NAND2X1_167 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_566_) );
NAND3X1 NAND3X1_49 ( .A(_564_), .B(_566_), .C(_565_), .Y(_567_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_561_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_562_) );
OAI21X1 OAI21X1_167 ( .A(_561_), .B(_562_), .C(1'b0), .Y(_563_) );
NAND2X1 NAND2X1_168 ( .A(_563_), .B(_567_), .Y(_39__0_) );
OAI21X1 OAI21X1_168 ( .A(_564_), .B(_561_), .C(_566_), .Y(_41__1_) );
INVX1 INVX1_120 ( .A(_41__1_), .Y(_571_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_572_) );
NAND2X1 NAND2X1_169 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_573_) );
NAND3X1 NAND3X1_50 ( .A(_571_), .B(_573_), .C(_572_), .Y(_574_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_568_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_569_) );
OAI21X1 OAI21X1_169 ( .A(_568_), .B(_569_), .C(_41__1_), .Y(_570_) );
NAND2X1 NAND2X1_170 ( .A(_570_), .B(_574_), .Y(_39__1_) );
OAI21X1 OAI21X1_170 ( .A(_571_), .B(_568_), .C(_573_), .Y(_41__2_) );
INVX1 INVX1_121 ( .A(_41__2_), .Y(_578_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_579_) );
NAND2X1 NAND2X1_171 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_580_) );
NAND3X1 NAND3X1_51 ( .A(_578_), .B(_580_), .C(_579_), .Y(_581_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_575_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_576_) );
OAI21X1 OAI21X1_171 ( .A(_575_), .B(_576_), .C(_41__2_), .Y(_577_) );
NAND2X1 NAND2X1_172 ( .A(_577_), .B(_581_), .Y(_39__2_) );
OAI21X1 OAI21X1_172 ( .A(_578_), .B(_575_), .C(_580_), .Y(_41__3_) );
INVX1 INVX1_122 ( .A(_41__3_), .Y(_585_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_586_) );
NAND2X1 NAND2X1_173 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_587_) );
NAND3X1 NAND3X1_52 ( .A(_585_), .B(_587_), .C(_586_), .Y(_588_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_582_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_583_) );
OAI21X1 OAI21X1_173 ( .A(_582_), .B(_583_), .C(_41__3_), .Y(_584_) );
NAND2X1 NAND2X1_174 ( .A(_584_), .B(_588_), .Y(_39__3_) );
OAI21X1 OAI21X1_174 ( .A(_585_), .B(_582_), .C(_587_), .Y(_37_) );
INVX1 INVX1_123 ( .A(1'b1), .Y(_592_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_593_) );
NAND2X1 NAND2X1_175 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_594_) );
NAND3X1 NAND3X1_53 ( .A(_592_), .B(_594_), .C(_593_), .Y(_595_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_589_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_590_) );
OAI21X1 OAI21X1_175 ( .A(_589_), .B(_590_), .C(1'b1), .Y(_591_) );
NAND2X1 NAND2X1_176 ( .A(_591_), .B(_595_), .Y(_40__0_) );
OAI21X1 OAI21X1_176 ( .A(_592_), .B(_589_), .C(_594_), .Y(_42__1_) );
INVX1 INVX1_124 ( .A(_42__1_), .Y(_599_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_600_) );
NAND2X1 NAND2X1_177 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_601_) );
NAND3X1 NAND3X1_54 ( .A(_599_), .B(_601_), .C(_600_), .Y(_602_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_596_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_597_) );
OAI21X1 OAI21X1_177 ( .A(_596_), .B(_597_), .C(_42__1_), .Y(_598_) );
NAND2X1 NAND2X1_178 ( .A(_598_), .B(_602_), .Y(_40__1_) );
OAI21X1 OAI21X1_178 ( .A(_599_), .B(_596_), .C(_601_), .Y(_42__2_) );
INVX1 INVX1_125 ( .A(_42__2_), .Y(_606_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_607_) );
NAND2X1 NAND2X1_179 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_608_) );
NAND3X1 NAND3X1_55 ( .A(_606_), .B(_608_), .C(_607_), .Y(_609_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_603_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_604_) );
OAI21X1 OAI21X1_179 ( .A(_603_), .B(_604_), .C(_42__2_), .Y(_605_) );
NAND2X1 NAND2X1_180 ( .A(_605_), .B(_609_), .Y(_40__2_) );
OAI21X1 OAI21X1_180 ( .A(_606_), .B(_603_), .C(_608_), .Y(_42__3_) );
INVX1 INVX1_126 ( .A(_42__3_), .Y(_613_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_614_) );
NAND2X1 NAND2X1_181 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_615_) );
NAND3X1 NAND3X1_56 ( .A(_613_), .B(_615_), .C(_614_), .Y(_616_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_610_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_611_) );
OAI21X1 OAI21X1_181 ( .A(_610_), .B(_611_), .C(_42__3_), .Y(_612_) );
NAND2X1 NAND2X1_182 ( .A(_612_), .B(_616_), .Y(_40__3_) );
OAI21X1 OAI21X1_182 ( .A(_613_), .B(_610_), .C(_615_), .Y(_38_) );
INVX1 INVX1_127 ( .A(1'b0), .Y(_620_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_621_) );
NAND2X1 NAND2X1_183 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_622_) );
NAND3X1 NAND3X1_57 ( .A(_620_), .B(_622_), .C(_621_), .Y(_623_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_617_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_618_) );
OAI21X1 OAI21X1_183 ( .A(_617_), .B(_618_), .C(1'b0), .Y(_619_) );
NAND2X1 NAND2X1_184 ( .A(_619_), .B(_623_), .Y(_45__0_) );
OAI21X1 OAI21X1_184 ( .A(_620_), .B(_617_), .C(_622_), .Y(_47__1_) );
INVX1 INVX1_128 ( .A(_47__1_), .Y(_627_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_628_) );
NAND2X1 NAND2X1_185 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_629_) );
NAND3X1 NAND3X1_58 ( .A(_627_), .B(_629_), .C(_628_), .Y(_630_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_624_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_625_) );
OAI21X1 OAI21X1_185 ( .A(_624_), .B(_625_), .C(_47__1_), .Y(_626_) );
NAND2X1 NAND2X1_186 ( .A(_626_), .B(_630_), .Y(_45__1_) );
OAI21X1 OAI21X1_186 ( .A(_627_), .B(_624_), .C(_629_), .Y(_47__2_) );
INVX1 INVX1_129 ( .A(_47__2_), .Y(_634_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_635_) );
NAND2X1 NAND2X1_187 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_636_) );
NAND3X1 NAND3X1_59 ( .A(_634_), .B(_636_), .C(_635_), .Y(_637_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_631_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_632_) );
OAI21X1 OAI21X1_187 ( .A(_631_), .B(_632_), .C(_47__2_), .Y(_633_) );
NAND2X1 NAND2X1_188 ( .A(_633_), .B(_637_), .Y(_45__2_) );
OAI21X1 OAI21X1_188 ( .A(_634_), .B(_631_), .C(_636_), .Y(_47__3_) );
INVX1 INVX1_130 ( .A(_47__3_), .Y(_641_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_642_) );
NAND2X1 NAND2X1_189 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_643_) );
NAND3X1 NAND3X1_60 ( .A(_641_), .B(_643_), .C(_642_), .Y(_644_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_638_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_639_) );
OAI21X1 OAI21X1_189 ( .A(_638_), .B(_639_), .C(_47__3_), .Y(_640_) );
NAND2X1 NAND2X1_190 ( .A(_640_), .B(_644_), .Y(_45__3_) );
OAI21X1 OAI21X1_190 ( .A(_641_), .B(_638_), .C(_643_), .Y(_43_) );
INVX1 INVX1_131 ( .A(1'b1), .Y(_648_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_649_) );
NAND2X1 NAND2X1_191 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_650_) );
NAND3X1 NAND3X1_61 ( .A(_648_), .B(_650_), .C(_649_), .Y(_651_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_645_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_646_) );
OAI21X1 OAI21X1_191 ( .A(_645_), .B(_646_), .C(1'b1), .Y(_647_) );
NAND2X1 NAND2X1_192 ( .A(_647_), .B(_651_), .Y(_46__0_) );
OAI21X1 OAI21X1_192 ( .A(_648_), .B(_645_), .C(_650_), .Y(_48__1_) );
INVX1 INVX1_132 ( .A(_48__1_), .Y(_655_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_656_) );
NAND2X1 NAND2X1_193 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_657_) );
NAND3X1 NAND3X1_62 ( .A(_655_), .B(_657_), .C(_656_), .Y(_658_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_652_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_653_) );
OAI21X1 OAI21X1_193 ( .A(_652_), .B(_653_), .C(_48__1_), .Y(_654_) );
NAND2X1 NAND2X1_194 ( .A(_654_), .B(_658_), .Y(_46__1_) );
OAI21X1 OAI21X1_194 ( .A(_655_), .B(_652_), .C(_657_), .Y(_48__2_) );
INVX1 INVX1_133 ( .A(_48__2_), .Y(_662_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_663_) );
NAND2X1 NAND2X1_195 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_664_) );
NAND3X1 NAND3X1_63 ( .A(_662_), .B(_664_), .C(_663_), .Y(_665_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_659_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_660_) );
OAI21X1 OAI21X1_195 ( .A(_659_), .B(_660_), .C(_48__2_), .Y(_661_) );
NAND2X1 NAND2X1_196 ( .A(_661_), .B(_665_), .Y(_46__2_) );
OAI21X1 OAI21X1_196 ( .A(_662_), .B(_659_), .C(_664_), .Y(_48__3_) );
INVX1 INVX1_134 ( .A(_48__3_), .Y(_669_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_670_) );
NAND2X1 NAND2X1_197 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_671_) );
NAND3X1 NAND3X1_64 ( .A(_669_), .B(_671_), .C(_670_), .Y(_672_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_666_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_667_) );
OAI21X1 OAI21X1_197 ( .A(_666_), .B(_667_), .C(_48__3_), .Y(_668_) );
NAND2X1 NAND2X1_198 ( .A(_668_), .B(_672_), .Y(_46__3_) );
OAI21X1 OAI21X1_198 ( .A(_669_), .B(_666_), .C(_671_), .Y(_44_) );
INVX1 INVX1_135 ( .A(1'b0), .Y(_676_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_677_) );
NAND2X1 NAND2X1_199 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_678_) );
NAND3X1 NAND3X1_65 ( .A(_676_), .B(_678_), .C(_677_), .Y(_679_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_673_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_674_) );
OAI21X1 OAI21X1_199 ( .A(_673_), .B(_674_), .C(1'b0), .Y(_675_) );
NAND2X1 NAND2X1_200 ( .A(_675_), .B(_679_), .Y(_51__0_) );
OAI21X1 OAI21X1_200 ( .A(_676_), .B(_673_), .C(_678_), .Y(_53__1_) );
INVX1 INVX1_136 ( .A(_53__1_), .Y(_683_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_684_) );
NAND2X1 NAND2X1_201 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_685_) );
NAND3X1 NAND3X1_66 ( .A(_683_), .B(_685_), .C(_684_), .Y(_686_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_680_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_681_) );
OAI21X1 OAI21X1_201 ( .A(_680_), .B(_681_), .C(_53__1_), .Y(_682_) );
NAND2X1 NAND2X1_202 ( .A(_682_), .B(_686_), .Y(_51__1_) );
OAI21X1 OAI21X1_202 ( .A(_683_), .B(_680_), .C(_685_), .Y(_53__2_) );
INVX1 INVX1_137 ( .A(_53__2_), .Y(_690_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_691_) );
NAND2X1 NAND2X1_203 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_692_) );
NAND3X1 NAND3X1_67 ( .A(_690_), .B(_692_), .C(_691_), .Y(_693_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_687_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_688_) );
OAI21X1 OAI21X1_203 ( .A(_687_), .B(_688_), .C(_53__2_), .Y(_689_) );
NAND2X1 NAND2X1_204 ( .A(_689_), .B(_693_), .Y(_51__2_) );
OAI21X1 OAI21X1_204 ( .A(_690_), .B(_687_), .C(_692_), .Y(_53__3_) );
INVX1 INVX1_138 ( .A(_53__3_), .Y(_697_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_698_) );
NAND2X1 NAND2X1_205 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_699_) );
NAND3X1 NAND3X1_68 ( .A(_697_), .B(_699_), .C(_698_), .Y(_700_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_694_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_695_) );
OAI21X1 OAI21X1_205 ( .A(_694_), .B(_695_), .C(_53__3_), .Y(_696_) );
NAND2X1 NAND2X1_206 ( .A(_696_), .B(_700_), .Y(_51__3_) );
OAI21X1 OAI21X1_206 ( .A(_697_), .B(_694_), .C(_699_), .Y(_49_) );
INVX1 INVX1_139 ( .A(1'b1), .Y(_704_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_705_) );
NAND2X1 NAND2X1_207 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_706_) );
NAND3X1 NAND3X1_69 ( .A(_704_), .B(_706_), .C(_705_), .Y(_707_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_701_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_702_) );
OAI21X1 OAI21X1_207 ( .A(_701_), .B(_702_), .C(1'b1), .Y(_703_) );
NAND2X1 NAND2X1_208 ( .A(_703_), .B(_707_), .Y(_52__0_) );
OAI21X1 OAI21X1_208 ( .A(_704_), .B(_701_), .C(_706_), .Y(_54__1_) );
INVX1 INVX1_140 ( .A(_54__1_), .Y(_711_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_712_) );
NAND2X1 NAND2X1_209 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_713_) );
NAND3X1 NAND3X1_70 ( .A(_711_), .B(_713_), .C(_712_), .Y(_714_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_708_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_709_) );
OAI21X1 OAI21X1_209 ( .A(_708_), .B(_709_), .C(_54__1_), .Y(_710_) );
NAND2X1 NAND2X1_210 ( .A(_710_), .B(_714_), .Y(_52__1_) );
OAI21X1 OAI21X1_210 ( .A(_711_), .B(_708_), .C(_713_), .Y(_54__2_) );
INVX1 INVX1_141 ( .A(_54__2_), .Y(_718_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_719_) );
NAND2X1 NAND2X1_211 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_720_) );
NAND3X1 NAND3X1_71 ( .A(_718_), .B(_720_), .C(_719_), .Y(_721_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_715_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_716_) );
OAI21X1 OAI21X1_211 ( .A(_715_), .B(_716_), .C(_54__2_), .Y(_717_) );
NAND2X1 NAND2X1_212 ( .A(_717_), .B(_721_), .Y(_52__2_) );
OAI21X1 OAI21X1_212 ( .A(_718_), .B(_715_), .C(_720_), .Y(_54__3_) );
INVX1 INVX1_142 ( .A(_54__3_), .Y(_725_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_726_) );
NAND2X1 NAND2X1_213 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_727_) );
NAND3X1 NAND3X1_72 ( .A(_725_), .B(_727_), .C(_726_), .Y(_728_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_722_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_723_) );
OAI21X1 OAI21X1_213 ( .A(_722_), .B(_723_), .C(_54__3_), .Y(_724_) );
NAND2X1 NAND2X1_214 ( .A(_724_), .B(_728_), .Y(_52__3_) );
OAI21X1 OAI21X1_214 ( .A(_725_), .B(_722_), .C(_727_), .Y(_50_) );
INVX1 INVX1_143 ( .A(1'b0), .Y(_732_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_733_) );
NAND2X1 NAND2X1_215 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_734_) );
NAND3X1 NAND3X1_73 ( .A(_732_), .B(_734_), .C(_733_), .Y(_735_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_729_) );
AND2X2 AND2X2_73 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_730_) );
OAI21X1 OAI21X1_215 ( .A(_729_), .B(_730_), .C(1'b0), .Y(_731_) );
NAND2X1 NAND2X1_216 ( .A(_731_), .B(_735_), .Y(_57__0_) );
OAI21X1 OAI21X1_216 ( .A(_732_), .B(_729_), .C(_734_), .Y(_59__1_) );
INVX1 INVX1_144 ( .A(_59__1_), .Y(_739_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_740_) );
NAND2X1 NAND2X1_217 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_741_) );
NAND3X1 NAND3X1_74 ( .A(_739_), .B(_741_), .C(_740_), .Y(_742_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_736_) );
AND2X2 AND2X2_74 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_737_) );
OAI21X1 OAI21X1_217 ( .A(_736_), .B(_737_), .C(_59__1_), .Y(_738_) );
NAND2X1 NAND2X1_218 ( .A(_738_), .B(_742_), .Y(_57__1_) );
OAI21X1 OAI21X1_218 ( .A(_739_), .B(_736_), .C(_741_), .Y(_59__2_) );
INVX1 INVX1_145 ( .A(_59__2_), .Y(_746_) );
OR2X2 OR2X2_75 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_747_) );
NAND2X1 NAND2X1_219 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_748_) );
NAND3X1 NAND3X1_75 ( .A(_746_), .B(_748_), .C(_747_), .Y(_749_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_743_) );
AND2X2 AND2X2_75 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_744_) );
OAI21X1 OAI21X1_219 ( .A(_743_), .B(_744_), .C(_59__2_), .Y(_745_) );
NAND2X1 NAND2X1_220 ( .A(_745_), .B(_749_), .Y(_57__2_) );
OAI21X1 OAI21X1_220 ( .A(_746_), .B(_743_), .C(_748_), .Y(_59__3_) );
INVX1 INVX1_146 ( .A(_59__3_), .Y(_753_) );
OR2X2 OR2X2_76 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_754_) );
NAND2X1 NAND2X1_221 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_755_) );
NAND3X1 NAND3X1_76 ( .A(_753_), .B(_755_), .C(_754_), .Y(_756_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_750_) );
AND2X2 AND2X2_76 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_751_) );
OAI21X1 OAI21X1_221 ( .A(_750_), .B(_751_), .C(_59__3_), .Y(_752_) );
NAND2X1 NAND2X1_222 ( .A(_752_), .B(_756_), .Y(_57__3_) );
OAI21X1 OAI21X1_222 ( .A(_753_), .B(_750_), .C(_755_), .Y(_55_) );
INVX1 INVX1_147 ( .A(1'b1), .Y(_760_) );
OR2X2 OR2X2_77 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_761_) );
NAND2X1 NAND2X1_223 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_762_) );
NAND3X1 NAND3X1_77 ( .A(_760_), .B(_762_), .C(_761_), .Y(_763_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_757_) );
AND2X2 AND2X2_77 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_758_) );
OAI21X1 OAI21X1_223 ( .A(_757_), .B(_758_), .C(1'b1), .Y(_759_) );
NAND2X1 NAND2X1_224 ( .A(_759_), .B(_763_), .Y(_58__0_) );
OAI21X1 OAI21X1_224 ( .A(_760_), .B(_757_), .C(_762_), .Y(_60__1_) );
INVX1 INVX1_148 ( .A(_60__1_), .Y(_767_) );
OR2X2 OR2X2_78 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_768_) );
NAND2X1 NAND2X1_225 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_769_) );
NAND3X1 NAND3X1_78 ( .A(_767_), .B(_769_), .C(_768_), .Y(_770_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_764_) );
AND2X2 AND2X2_78 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_765_) );
OAI21X1 OAI21X1_225 ( .A(_764_), .B(_765_), .C(_60__1_), .Y(_766_) );
NAND2X1 NAND2X1_226 ( .A(_766_), .B(_770_), .Y(_58__1_) );
OAI21X1 OAI21X1_226 ( .A(_767_), .B(_764_), .C(_769_), .Y(_60__2_) );
INVX1 INVX1_149 ( .A(_60__2_), .Y(_774_) );
OR2X2 OR2X2_79 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_775_) );
NAND2X1 NAND2X1_227 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_776_) );
NAND3X1 NAND3X1_79 ( .A(_774_), .B(_776_), .C(_775_), .Y(_777_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_771_) );
AND2X2 AND2X2_79 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_772_) );
OAI21X1 OAI21X1_227 ( .A(_771_), .B(_772_), .C(_60__2_), .Y(_773_) );
NAND2X1 NAND2X1_228 ( .A(_773_), .B(_777_), .Y(_58__2_) );
OAI21X1 OAI21X1_228 ( .A(_774_), .B(_771_), .C(_776_), .Y(_60__3_) );
INVX1 INVX1_150 ( .A(_60__3_), .Y(_781_) );
OR2X2 OR2X2_80 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_782_) );
NAND2X1 NAND2X1_229 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_783_) );
NAND3X1 NAND3X1_80 ( .A(_781_), .B(_783_), .C(_782_), .Y(_784_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_778_) );
AND2X2 AND2X2_80 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_779_) );
OAI21X1 OAI21X1_229 ( .A(_778_), .B(_779_), .C(_60__3_), .Y(_780_) );
NAND2X1 NAND2X1_230 ( .A(_780_), .B(_784_), .Y(_58__3_) );
OAI21X1 OAI21X1_230 ( .A(_781_), .B(_778_), .C(_783_), .Y(_56_) );
INVX1 INVX1_151 ( .A(1'b0), .Y(_788_) );
OR2X2 OR2X2_81 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_789_) );
NAND2X1 NAND2X1_231 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_790_) );
NAND3X1 NAND3X1_81 ( .A(_788_), .B(_790_), .C(_789_), .Y(_791_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_785_) );
AND2X2 AND2X2_81 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_786_) );
OAI21X1 OAI21X1_231 ( .A(_785_), .B(_786_), .C(1'b0), .Y(_787_) );
NAND2X1 NAND2X1_232 ( .A(_787_), .B(_791_), .Y(_63__0_) );
OAI21X1 OAI21X1_232 ( .A(_788_), .B(_785_), .C(_790_), .Y(_65__1_) );
INVX1 INVX1_152 ( .A(_65__1_), .Y(_795_) );
OR2X2 OR2X2_82 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_796_) );
NAND2X1 NAND2X1_233 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_797_) );
NAND3X1 NAND3X1_82 ( .A(_795_), .B(_797_), .C(_796_), .Y(_798_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_792_) );
AND2X2 AND2X2_82 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_793_) );
OAI21X1 OAI21X1_233 ( .A(_792_), .B(_793_), .C(_65__1_), .Y(_794_) );
NAND2X1 NAND2X1_234 ( .A(_794_), .B(_798_), .Y(_63__1_) );
OAI21X1 OAI21X1_234 ( .A(_795_), .B(_792_), .C(_797_), .Y(_65__2_) );
INVX1 INVX1_153 ( .A(_65__2_), .Y(_802_) );
OR2X2 OR2X2_83 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_803_) );
NAND2X1 NAND2X1_235 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_804_) );
NAND3X1 NAND3X1_83 ( .A(_802_), .B(_804_), .C(_803_), .Y(_805_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_799_) );
AND2X2 AND2X2_83 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_800_) );
OAI21X1 OAI21X1_235 ( .A(_799_), .B(_800_), .C(_65__2_), .Y(_801_) );
NAND2X1 NAND2X1_236 ( .A(_801_), .B(_805_), .Y(_63__2_) );
OAI21X1 OAI21X1_236 ( .A(_802_), .B(_799_), .C(_804_), .Y(_65__3_) );
INVX1 INVX1_154 ( .A(_65__3_), .Y(_809_) );
OR2X2 OR2X2_84 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_810_) );
NAND2X1 NAND2X1_237 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_811_) );
NAND3X1 NAND3X1_84 ( .A(_809_), .B(_811_), .C(_810_), .Y(_812_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_806_) );
AND2X2 AND2X2_84 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_807_) );
OAI21X1 OAI21X1_237 ( .A(_806_), .B(_807_), .C(_65__3_), .Y(_808_) );
NAND2X1 NAND2X1_238 ( .A(_808_), .B(_812_), .Y(_63__3_) );
OAI21X1 OAI21X1_238 ( .A(_809_), .B(_806_), .C(_811_), .Y(_61_) );
INVX1 INVX1_155 ( .A(1'b1), .Y(_816_) );
OR2X2 OR2X2_85 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_817_) );
NAND2X1 NAND2X1_239 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_818_) );
NAND3X1 NAND3X1_85 ( .A(_816_), .B(_818_), .C(_817_), .Y(_819_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_813_) );
AND2X2 AND2X2_85 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_814_) );
OAI21X1 OAI21X1_239 ( .A(_813_), .B(_814_), .C(1'b1), .Y(_815_) );
NAND2X1 NAND2X1_240 ( .A(_815_), .B(_819_), .Y(_64__0_) );
OAI21X1 OAI21X1_240 ( .A(_816_), .B(_813_), .C(_818_), .Y(_66__1_) );
INVX1 INVX1_156 ( .A(_66__1_), .Y(_823_) );
OR2X2 OR2X2_86 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_824_) );
NAND2X1 NAND2X1_241 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_825_) );
NAND3X1 NAND3X1_86 ( .A(_823_), .B(_825_), .C(_824_), .Y(_826_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_820_) );
AND2X2 AND2X2_86 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_821_) );
OAI21X1 OAI21X1_241 ( .A(_820_), .B(_821_), .C(_66__1_), .Y(_822_) );
NAND2X1 NAND2X1_242 ( .A(_822_), .B(_826_), .Y(_64__1_) );
OAI21X1 OAI21X1_242 ( .A(_823_), .B(_820_), .C(_825_), .Y(_66__2_) );
INVX1 INVX1_157 ( .A(_66__2_), .Y(_830_) );
OR2X2 OR2X2_87 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_831_) );
NAND2X1 NAND2X1_243 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_832_) );
NAND3X1 NAND3X1_87 ( .A(_830_), .B(_832_), .C(_831_), .Y(_833_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_827_) );
AND2X2 AND2X2_87 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_828_) );
OAI21X1 OAI21X1_243 ( .A(_827_), .B(_828_), .C(_66__2_), .Y(_829_) );
NAND2X1 NAND2X1_244 ( .A(_829_), .B(_833_), .Y(_64__2_) );
OAI21X1 OAI21X1_244 ( .A(_830_), .B(_827_), .C(_832_), .Y(_66__3_) );
INVX1 INVX1_158 ( .A(_66__3_), .Y(_837_) );
OR2X2 OR2X2_88 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_838_) );
NAND2X1 NAND2X1_245 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_839_) );
NAND3X1 NAND3X1_88 ( .A(_837_), .B(_839_), .C(_838_), .Y(_840_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_834_) );
AND2X2 AND2X2_88 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_835_) );
OAI21X1 OAI21X1_245 ( .A(_834_), .B(_835_), .C(_66__3_), .Y(_836_) );
NAND2X1 NAND2X1_246 ( .A(_836_), .B(_840_), .Y(_64__3_) );
OAI21X1 OAI21X1_246 ( .A(_837_), .B(_834_), .C(_839_), .Y(_62_) );
INVX1 INVX1_159 ( .A(1'b0), .Y(_844_) );
OR2X2 OR2X2_89 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_845_) );
NAND2X1 NAND2X1_247 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_846_) );
NAND3X1 NAND3X1_89 ( .A(_844_), .B(_846_), .C(_845_), .Y(_847_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_841_) );
AND2X2 AND2X2_89 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_842_) );
OAI21X1 OAI21X1_247 ( .A(_841_), .B(_842_), .C(1'b0), .Y(_843_) );
NAND2X1 NAND2X1_248 ( .A(_843_), .B(_847_), .Y(_69__0_) );
OAI21X1 OAI21X1_248 ( .A(_844_), .B(_841_), .C(_846_), .Y(_71__1_) );
INVX1 INVX1_160 ( .A(_71__1_), .Y(_851_) );
OR2X2 OR2X2_90 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_852_) );
NAND2X1 NAND2X1_249 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_853_) );
NAND3X1 NAND3X1_90 ( .A(_851_), .B(_853_), .C(_852_), .Y(_854_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_848_) );
AND2X2 AND2X2_90 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_849_) );
OAI21X1 OAI21X1_249 ( .A(_848_), .B(_849_), .C(_71__1_), .Y(_850_) );
NAND2X1 NAND2X1_250 ( .A(_850_), .B(_854_), .Y(_69__1_) );
OAI21X1 OAI21X1_250 ( .A(_851_), .B(_848_), .C(_853_), .Y(_71__2_) );
INVX1 INVX1_161 ( .A(_71__2_), .Y(_858_) );
OR2X2 OR2X2_91 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_859_) );
NAND2X1 NAND2X1_251 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_860_) );
NAND3X1 NAND3X1_91 ( .A(_858_), .B(_860_), .C(_859_), .Y(_861_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_855_) );
AND2X2 AND2X2_91 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_856_) );
OAI21X1 OAI21X1_251 ( .A(_855_), .B(_856_), .C(_71__2_), .Y(_857_) );
NAND2X1 NAND2X1_252 ( .A(_857_), .B(_861_), .Y(_69__2_) );
OAI21X1 OAI21X1_252 ( .A(_858_), .B(_855_), .C(_860_), .Y(_71__3_) );
INVX1 INVX1_162 ( .A(_71__3_), .Y(_865_) );
OR2X2 OR2X2_92 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_866_) );
NAND2X1 NAND2X1_253 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_867_) );
NAND3X1 NAND3X1_92 ( .A(_865_), .B(_867_), .C(_866_), .Y(_868_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_862_) );
AND2X2 AND2X2_92 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_863_) );
OAI21X1 OAI21X1_253 ( .A(_862_), .B(_863_), .C(_71__3_), .Y(_864_) );
NAND2X1 NAND2X1_254 ( .A(_864_), .B(_868_), .Y(_69__3_) );
OAI21X1 OAI21X1_254 ( .A(_865_), .B(_862_), .C(_867_), .Y(_67_) );
INVX1 INVX1_163 ( .A(1'b1), .Y(_872_) );
OR2X2 OR2X2_93 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_873_) );
NAND2X1 NAND2X1_255 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_874_) );
NAND3X1 NAND3X1_93 ( .A(_872_), .B(_874_), .C(_873_), .Y(_875_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_869_) );
AND2X2 AND2X2_93 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_870_) );
OAI21X1 OAI21X1_255 ( .A(_869_), .B(_870_), .C(1'b1), .Y(_871_) );
NAND2X1 NAND2X1_256 ( .A(_871_), .B(_875_), .Y(_70__0_) );
OAI21X1 OAI21X1_256 ( .A(_872_), .B(_869_), .C(_874_), .Y(_72__1_) );
INVX1 INVX1_164 ( .A(_72__1_), .Y(_879_) );
OR2X2 OR2X2_94 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_880_) );
NAND2X1 NAND2X1_257 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_881_) );
NAND3X1 NAND3X1_94 ( .A(_879_), .B(_881_), .C(_880_), .Y(_882_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_876_) );
AND2X2 AND2X2_94 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_877_) );
OAI21X1 OAI21X1_257 ( .A(_876_), .B(_877_), .C(_72__1_), .Y(_878_) );
NAND2X1 NAND2X1_258 ( .A(_878_), .B(_882_), .Y(_70__1_) );
OAI21X1 OAI21X1_258 ( .A(_879_), .B(_876_), .C(_881_), .Y(_72__2_) );
INVX1 INVX1_165 ( .A(_72__2_), .Y(_886_) );
OR2X2 OR2X2_95 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_887_) );
NAND2X1 NAND2X1_259 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_888_) );
NAND3X1 NAND3X1_95 ( .A(_886_), .B(_888_), .C(_887_), .Y(_889_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_883_) );
AND2X2 AND2X2_95 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_884_) );
OAI21X1 OAI21X1_259 ( .A(_883_), .B(_884_), .C(_72__2_), .Y(_885_) );
NAND2X1 NAND2X1_260 ( .A(_885_), .B(_889_), .Y(_70__2_) );
OAI21X1 OAI21X1_260 ( .A(_886_), .B(_883_), .C(_888_), .Y(_72__3_) );
INVX1 INVX1_166 ( .A(_72__3_), .Y(_893_) );
OR2X2 OR2X2_96 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_894_) );
NAND2X1 NAND2X1_261 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_895_) );
NAND3X1 NAND3X1_96 ( .A(_893_), .B(_895_), .C(_894_), .Y(_896_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_890_) );
AND2X2 AND2X2_96 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_891_) );
OAI21X1 OAI21X1_261 ( .A(_890_), .B(_891_), .C(_72__3_), .Y(_892_) );
NAND2X1 NAND2X1_262 ( .A(_892_), .B(_896_), .Y(_70__3_) );
OAI21X1 OAI21X1_262 ( .A(_893_), .B(_890_), .C(_895_), .Y(_68_) );
INVX1 INVX1_167 ( .A(1'b0), .Y(_900_) );
OR2X2 OR2X2_97 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_901_) );
NAND2X1 NAND2X1_263 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_902_) );
NAND3X1 NAND3X1_97 ( .A(_900_), .B(_902_), .C(_901_), .Y(_903_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_897_) );
AND2X2 AND2X2_97 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_898_) );
OAI21X1 OAI21X1_263 ( .A(_897_), .B(_898_), .C(1'b0), .Y(_899_) );
NAND2X1 NAND2X1_264 ( .A(_899_), .B(_903_), .Y(_75__0_) );
OAI21X1 OAI21X1_264 ( .A(_900_), .B(_897_), .C(_902_), .Y(_77__1_) );
INVX1 INVX1_168 ( .A(_77__1_), .Y(_907_) );
OR2X2 OR2X2_98 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_908_) );
NAND2X1 NAND2X1_265 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_909_) );
NAND3X1 NAND3X1_98 ( .A(_907_), .B(_909_), .C(_908_), .Y(_910_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_904_) );
AND2X2 AND2X2_98 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_905_) );
OAI21X1 OAI21X1_265 ( .A(_904_), .B(_905_), .C(_77__1_), .Y(_906_) );
NAND2X1 NAND2X1_266 ( .A(_906_), .B(_910_), .Y(_75__1_) );
OAI21X1 OAI21X1_266 ( .A(_907_), .B(_904_), .C(_909_), .Y(_77__2_) );
INVX1 INVX1_169 ( .A(_77__2_), .Y(_914_) );
OR2X2 OR2X2_99 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_915_) );
NAND2X1 NAND2X1_267 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_916_) );
NAND3X1 NAND3X1_99 ( .A(_914_), .B(_916_), .C(_915_), .Y(_917_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_911_) );
AND2X2 AND2X2_99 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_912_) );
OAI21X1 OAI21X1_267 ( .A(_911_), .B(_912_), .C(_77__2_), .Y(_913_) );
NAND2X1 NAND2X1_268 ( .A(_913_), .B(_917_), .Y(_75__2_) );
OAI21X1 OAI21X1_268 ( .A(_914_), .B(_911_), .C(_916_), .Y(_77__3_) );
INVX1 INVX1_170 ( .A(_77__3_), .Y(_921_) );
OR2X2 OR2X2_100 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_922_) );
NAND2X1 NAND2X1_269 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_923_) );
NAND3X1 NAND3X1_100 ( .A(_921_), .B(_923_), .C(_922_), .Y(_924_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_918_) );
AND2X2 AND2X2_100 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_919_) );
OAI21X1 OAI21X1_269 ( .A(_918_), .B(_919_), .C(_77__3_), .Y(_920_) );
NAND2X1 NAND2X1_270 ( .A(_920_), .B(_924_), .Y(_75__3_) );
OAI21X1 OAI21X1_270 ( .A(_921_), .B(_918_), .C(_923_), .Y(_73_) );
INVX1 INVX1_171 ( .A(1'b1), .Y(_928_) );
OR2X2 OR2X2_101 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_929_) );
NAND2X1 NAND2X1_271 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_930_) );
NAND3X1 NAND3X1_101 ( .A(_928_), .B(_930_), .C(_929_), .Y(_931_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_925_) );
AND2X2 AND2X2_101 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_926_) );
OAI21X1 OAI21X1_271 ( .A(_925_), .B(_926_), .C(1'b1), .Y(_927_) );
NAND2X1 NAND2X1_272 ( .A(_927_), .B(_931_), .Y(_76__0_) );
OAI21X1 OAI21X1_272 ( .A(_928_), .B(_925_), .C(_930_), .Y(_78__1_) );
INVX1 INVX1_172 ( .A(_78__1_), .Y(_935_) );
OR2X2 OR2X2_102 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_936_) );
NAND2X1 NAND2X1_273 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_937_) );
NAND3X1 NAND3X1_102 ( .A(_935_), .B(_937_), .C(_936_), .Y(_938_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_932_) );
AND2X2 AND2X2_102 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_933_) );
OAI21X1 OAI21X1_273 ( .A(_932_), .B(_933_), .C(_78__1_), .Y(_934_) );
NAND2X1 NAND2X1_274 ( .A(_934_), .B(_938_), .Y(_76__1_) );
OAI21X1 OAI21X1_274 ( .A(_935_), .B(_932_), .C(_937_), .Y(_78__2_) );
INVX1 INVX1_173 ( .A(_78__2_), .Y(_942_) );
OR2X2 OR2X2_103 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_943_) );
NAND2X1 NAND2X1_275 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_944_) );
NAND3X1 NAND3X1_103 ( .A(_942_), .B(_944_), .C(_943_), .Y(_945_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_939_) );
AND2X2 AND2X2_103 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_940_) );
OAI21X1 OAI21X1_275 ( .A(_939_), .B(_940_), .C(_78__2_), .Y(_941_) );
NAND2X1 NAND2X1_276 ( .A(_941_), .B(_945_), .Y(_76__2_) );
OAI21X1 OAI21X1_276 ( .A(_942_), .B(_939_), .C(_944_), .Y(_78__3_) );
INVX1 INVX1_174 ( .A(_78__3_), .Y(_949_) );
OR2X2 OR2X2_104 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_950_) );
NAND2X1 NAND2X1_277 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_951_) );
NAND3X1 NAND3X1_104 ( .A(_949_), .B(_951_), .C(_950_), .Y(_952_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_946_) );
AND2X2 AND2X2_104 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_947_) );
OAI21X1 OAI21X1_277 ( .A(_946_), .B(_947_), .C(_78__3_), .Y(_948_) );
NAND2X1 NAND2X1_278 ( .A(_948_), .B(_952_), .Y(_76__3_) );
OAI21X1 OAI21X1_278 ( .A(_949_), .B(_946_), .C(_951_), .Y(_74_) );
INVX1 INVX1_175 ( .A(1'b0), .Y(_956_) );
OR2X2 OR2X2_105 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_957_) );
NAND2X1 NAND2X1_279 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_958_) );
NAND3X1 NAND3X1_105 ( .A(_956_), .B(_958_), .C(_957_), .Y(_959_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_953_) );
AND2X2 AND2X2_105 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_954_) );
OAI21X1 OAI21X1_279 ( .A(_953_), .B(_954_), .C(1'b0), .Y(_955_) );
NAND2X1 NAND2X1_280 ( .A(_955_), .B(_959_), .Y(_81__0_) );
OAI21X1 OAI21X1_280 ( .A(_956_), .B(_953_), .C(_958_), .Y(_83__1_) );
INVX1 INVX1_176 ( .A(_83__1_), .Y(_963_) );
OR2X2 OR2X2_106 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_964_) );
NAND2X1 NAND2X1_281 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_965_) );
NAND3X1 NAND3X1_106 ( .A(_963_), .B(_965_), .C(_964_), .Y(_966_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_960_) );
AND2X2 AND2X2_106 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_961_) );
OAI21X1 OAI21X1_281 ( .A(_960_), .B(_961_), .C(_83__1_), .Y(_962_) );
NAND2X1 NAND2X1_282 ( .A(_962_), .B(_966_), .Y(_81__1_) );
OAI21X1 OAI21X1_282 ( .A(_963_), .B(_960_), .C(_965_), .Y(_83__2_) );
INVX1 INVX1_177 ( .A(_83__2_), .Y(_970_) );
OR2X2 OR2X2_107 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_971_) );
NAND2X1 NAND2X1_283 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_972_) );
NAND3X1 NAND3X1_107 ( .A(_970_), .B(_972_), .C(_971_), .Y(_973_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_967_) );
AND2X2 AND2X2_107 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_968_) );
OAI21X1 OAI21X1_283 ( .A(_967_), .B(_968_), .C(_83__2_), .Y(_969_) );
NAND2X1 NAND2X1_284 ( .A(_969_), .B(_973_), .Y(_81__2_) );
OAI21X1 OAI21X1_284 ( .A(_970_), .B(_967_), .C(_972_), .Y(_83__3_) );
INVX1 INVX1_178 ( .A(_83__3_), .Y(_977_) );
OR2X2 OR2X2_108 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_978_) );
NAND2X1 NAND2X1_285 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_979_) );
NAND3X1 NAND3X1_108 ( .A(_977_), .B(_979_), .C(_978_), .Y(_980_) );
NOR2X1 NOR2X1_108 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_974_) );
AND2X2 AND2X2_108 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_975_) );
OAI21X1 OAI21X1_285 ( .A(_974_), .B(_975_), .C(_83__3_), .Y(_976_) );
NAND2X1 NAND2X1_286 ( .A(_976_), .B(_980_), .Y(_81__3_) );
OAI21X1 OAI21X1_286 ( .A(_977_), .B(_974_), .C(_979_), .Y(_79_) );
INVX1 INVX1_179 ( .A(1'b1), .Y(_984_) );
OR2X2 OR2X2_109 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_985_) );
NAND2X1 NAND2X1_287 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_986_) );
NAND3X1 NAND3X1_109 ( .A(_984_), .B(_986_), .C(_985_), .Y(_987_) );
NOR2X1 NOR2X1_109 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_981_) );
AND2X2 AND2X2_109 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_982_) );
OAI21X1 OAI21X1_287 ( .A(_981_), .B(_982_), .C(1'b1), .Y(_983_) );
NAND2X1 NAND2X1_288 ( .A(_983_), .B(_987_), .Y(_82__0_) );
OAI21X1 OAI21X1_288 ( .A(_984_), .B(_981_), .C(_986_), .Y(_84__1_) );
INVX1 INVX1_180 ( .A(_84__1_), .Y(_991_) );
OR2X2 OR2X2_110 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_992_) );
NAND2X1 NAND2X1_289 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_993_) );
NAND3X1 NAND3X1_110 ( .A(_991_), .B(_993_), .C(_992_), .Y(_994_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_988_) );
AND2X2 AND2X2_110 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_989_) );
OAI21X1 OAI21X1_289 ( .A(_988_), .B(_989_), .C(_84__1_), .Y(_990_) );
NAND2X1 NAND2X1_290 ( .A(_990_), .B(_994_), .Y(_82__1_) );
OAI21X1 OAI21X1_290 ( .A(_991_), .B(_988_), .C(_993_), .Y(_84__2_) );
INVX1 INVX1_181 ( .A(_84__2_), .Y(_998_) );
OR2X2 OR2X2_111 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_999_) );
NAND2X1 NAND2X1_291 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_1000_) );
NAND3X1 NAND3X1_111 ( .A(_998_), .B(_1000_), .C(_999_), .Y(_1001_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_995_) );
AND2X2 AND2X2_111 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_996_) );
OAI21X1 OAI21X1_291 ( .A(_995_), .B(_996_), .C(_84__2_), .Y(_997_) );
NAND2X1 NAND2X1_292 ( .A(_997_), .B(_1001_), .Y(_82__2_) );
OAI21X1 OAI21X1_292 ( .A(_998_), .B(_995_), .C(_1000_), .Y(_84__3_) );
INVX1 INVX1_182 ( .A(_84__3_), .Y(_1005_) );
OR2X2 OR2X2_112 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_1006_) );
NAND2X1 NAND2X1_293 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_1007_) );
NAND3X1 NAND3X1_112 ( .A(_1005_), .B(_1007_), .C(_1006_), .Y(_1008_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_1002_) );
AND2X2 AND2X2_112 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_1003_) );
OAI21X1 OAI21X1_293 ( .A(_1002_), .B(_1003_), .C(_84__3_), .Y(_1004_) );
NAND2X1 NAND2X1_294 ( .A(_1004_), .B(_1008_), .Y(_82__3_) );
OAI21X1 OAI21X1_294 ( .A(_1005_), .B(_1002_), .C(_1007_), .Y(_80_) );
INVX1 INVX1_183 ( .A(1'b0), .Y(_1012_) );
OR2X2 OR2X2_113 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1013_) );
NAND2X1 NAND2X1_295 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1014_) );
NAND3X1 NAND3X1_113 ( .A(_1012_), .B(_1014_), .C(_1013_), .Y(_1015_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1009_) );
AND2X2 AND2X2_113 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1010_) );
OAI21X1 OAI21X1_295 ( .A(_1009_), .B(_1010_), .C(1'b0), .Y(_1011_) );
NAND2X1 NAND2X1_296 ( .A(_1011_), .B(_1015_), .Y(_0__0_) );
OAI21X1 OAI21X1_296 ( .A(_1012_), .B(_1009_), .C(_1014_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_184 ( .A(rca_inst_w_CARRY_1_), .Y(_1019_) );
OR2X2 OR2X2_114 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1020_) );
NAND2X1 NAND2X1_297 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1021_) );
NAND3X1 NAND3X1_114 ( .A(_1019_), .B(_1021_), .C(_1020_), .Y(_1022_) );
NOR2X1 NOR2X1_114 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1016_) );
AND2X2 AND2X2_114 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1017_) );
OAI21X1 OAI21X1_297 ( .A(_1016_), .B(_1017_), .C(rca_inst_w_CARRY_1_), .Y(_1018_) );
NAND2X1 NAND2X1_298 ( .A(_1018_), .B(_1022_), .Y(_0__1_) );
OAI21X1 OAI21X1_298 ( .A(_1019_), .B(_1016_), .C(_1021_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_185 ( .A(rca_inst_w_CARRY_2_), .Y(_1026_) );
OR2X2 OR2X2_115 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1027_) );
NAND2X1 NAND2X1_299 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1028_) );
NAND3X1 NAND3X1_115 ( .A(_1026_), .B(_1028_), .C(_1027_), .Y(_1029_) );
NOR2X1 NOR2X1_115 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1023_) );
AND2X2 AND2X2_115 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1024_) );
OAI21X1 OAI21X1_299 ( .A(_1023_), .B(_1024_), .C(rca_inst_w_CARRY_2_), .Y(_1025_) );
NAND2X1 NAND2X1_300 ( .A(_1025_), .B(_1029_), .Y(_0__2_) );
OAI21X1 OAI21X1_300 ( .A(_1026_), .B(_1023_), .C(_1028_), .Y(rca_inst_w_CARRY_3_) );
INVX1 INVX1_186 ( .A(rca_inst_w_CARRY_3_), .Y(_1033_) );
OR2X2 OR2X2_116 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_1034_) );
NAND2X1 NAND2X1_301 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_1035_) );
NAND3X1 NAND3X1_116 ( .A(_1033_), .B(_1035_), .C(_1034_), .Y(_1036_) );
NOR2X1 NOR2X1_116 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_1030_) );
AND2X2 AND2X2_116 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_1031_) );
OAI21X1 OAI21X1_301 ( .A(_1030_), .B(_1031_), .C(rca_inst_w_CARRY_3_), .Y(_1032_) );
NAND2X1 NAND2X1_302 ( .A(_1032_), .B(_1036_), .Y(_0__3_) );
OAI21X1 OAI21X1_302 ( .A(_1033_), .B(_1030_), .C(_1035_), .Y(rca_inst_cout) );
BUFX2 BUFX2_62 ( .A(1'b0), .Y(_5__0_) );
BUFX2 BUFX2_63 ( .A(_1_), .Y(_5__4_) );
BUFX2 BUFX2_64 ( .A(1'b1), .Y(_6__0_) );
BUFX2 BUFX2_65 ( .A(_2_), .Y(_6__4_) );
BUFX2 BUFX2_66 ( .A(1'b0), .Y(_11__0_) );
BUFX2 BUFX2_67 ( .A(_7_), .Y(_11__4_) );
BUFX2 BUFX2_68 ( .A(1'b1), .Y(_12__0_) );
BUFX2 BUFX2_69 ( .A(_8_), .Y(_12__4_) );
BUFX2 BUFX2_70 ( .A(1'b0), .Y(_17__0_) );
BUFX2 BUFX2_71 ( .A(_13_), .Y(_17__4_) );
BUFX2 BUFX2_72 ( .A(1'b1), .Y(_18__0_) );
BUFX2 BUFX2_73 ( .A(_14_), .Y(_18__4_) );
BUFX2 BUFX2_74 ( .A(1'b0), .Y(_23__0_) );
BUFX2 BUFX2_75 ( .A(_19_), .Y(_23__4_) );
BUFX2 BUFX2_76 ( .A(1'b1), .Y(_24__0_) );
BUFX2 BUFX2_77 ( .A(_20_), .Y(_24__4_) );
BUFX2 BUFX2_78 ( .A(1'b0), .Y(_29__0_) );
BUFX2 BUFX2_79 ( .A(_25_), .Y(_29__4_) );
BUFX2 BUFX2_80 ( .A(1'b1), .Y(_30__0_) );
BUFX2 BUFX2_81 ( .A(_26_), .Y(_30__4_) );
BUFX2 BUFX2_82 ( .A(1'b0), .Y(_35__0_) );
BUFX2 BUFX2_83 ( .A(_31_), .Y(_35__4_) );
BUFX2 BUFX2_84 ( .A(1'b1), .Y(_36__0_) );
BUFX2 BUFX2_85 ( .A(_32_), .Y(_36__4_) );
BUFX2 BUFX2_86 ( .A(1'b0), .Y(_41__0_) );
BUFX2 BUFX2_87 ( .A(_37_), .Y(_41__4_) );
BUFX2 BUFX2_88 ( .A(1'b1), .Y(_42__0_) );
BUFX2 BUFX2_89 ( .A(_38_), .Y(_42__4_) );
BUFX2 BUFX2_90 ( .A(1'b0), .Y(_47__0_) );
BUFX2 BUFX2_91 ( .A(_43_), .Y(_47__4_) );
BUFX2 BUFX2_92 ( .A(1'b1), .Y(_48__0_) );
BUFX2 BUFX2_93 ( .A(_44_), .Y(_48__4_) );
BUFX2 BUFX2_94 ( .A(1'b0), .Y(_53__0_) );
BUFX2 BUFX2_95 ( .A(_49_), .Y(_53__4_) );
BUFX2 BUFX2_96 ( .A(1'b1), .Y(_54__0_) );
BUFX2 BUFX2_97 ( .A(_50_), .Y(_54__4_) );
BUFX2 BUFX2_98 ( .A(1'b0), .Y(_59__0_) );
BUFX2 BUFX2_99 ( .A(_55_), .Y(_59__4_) );
BUFX2 BUFX2_100 ( .A(1'b1), .Y(_60__0_) );
BUFX2 BUFX2_101 ( .A(_56_), .Y(_60__4_) );
BUFX2 BUFX2_102 ( .A(1'b0), .Y(_65__0_) );
BUFX2 BUFX2_103 ( .A(_61_), .Y(_65__4_) );
BUFX2 BUFX2_104 ( .A(1'b1), .Y(_66__0_) );
BUFX2 BUFX2_105 ( .A(_62_), .Y(_66__4_) );
BUFX2 BUFX2_106 ( .A(1'b0), .Y(_71__0_) );
BUFX2 BUFX2_107 ( .A(_67_), .Y(_71__4_) );
BUFX2 BUFX2_108 ( .A(1'b1), .Y(_72__0_) );
BUFX2 BUFX2_109 ( .A(_68_), .Y(_72__4_) );
BUFX2 BUFX2_110 ( .A(1'b0), .Y(_77__0_) );
BUFX2 BUFX2_111 ( .A(_73_), .Y(_77__4_) );
BUFX2 BUFX2_112 ( .A(1'b1), .Y(_78__0_) );
BUFX2 BUFX2_113 ( .A(_74_), .Y(_78__4_) );
BUFX2 BUFX2_114 ( .A(1'b0), .Y(_83__0_) );
BUFX2 BUFX2_115 ( .A(_79_), .Y(_83__4_) );
BUFX2 BUFX2_116 ( .A(1'b1), .Y(_84__0_) );
BUFX2 BUFX2_117 ( .A(_80_), .Y(_84__4_) );
BUFX2 BUFX2_118 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_119 ( .A(rca_inst_cout), .Y(rca_inst_w_CARRY_4_) );
BUFX2 BUFX2_120 ( .A(rca_inst_cout), .Y(w_cout_0_) );
endmodule
