module csa_37bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output cout;

INVX1 INVX1_1 ( .A(_24__2_), .Y(_309_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_310_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_311_) );
NAND3X1 NAND3X1_1 ( .A(_309_), .B(_311_), .C(_310_), .Y(_312_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_306_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_307_) );
OAI21X1 OAI21X1_1 ( .A(_306_), .B(_307_), .C(_24__2_), .Y(_308_) );
NAND2X1 NAND2X1_2 ( .A(_308_), .B(_312_), .Y(_22__2_) );
OAI21X1 OAI21X1_2 ( .A(_309_), .B(_306_), .C(_311_), .Y(_24__3_) );
INVX1 INVX1_2 ( .A(_25_), .Y(_313_) );
NAND2X1 NAND2X1_3 ( .A(_26_), .B(w_cout_4_), .Y(_314_) );
OAI21X1 OAI21X1_3 ( .A(w_cout_4_), .B(_313_), .C(_314_), .Y(w_cout_5_) );
INVX1 INVX1_3 ( .A(_27__0_), .Y(_315_) );
NAND2X1 NAND2X1_4 ( .A(_28__0_), .B(w_cout_4_), .Y(_316_) );
OAI21X1 OAI21X1_4 ( .A(w_cout_4_), .B(_315_), .C(_316_), .Y(_0__20_) );
INVX1 INVX1_4 ( .A(_27__1_), .Y(_317_) );
NAND2X1 NAND2X1_5 ( .A(w_cout_4_), .B(_28__1_), .Y(_318_) );
OAI21X1 OAI21X1_5 ( .A(w_cout_4_), .B(_317_), .C(_318_), .Y(_0__21_) );
INVX1 INVX1_5 ( .A(_27__2_), .Y(_319_) );
NAND2X1 NAND2X1_6 ( .A(w_cout_4_), .B(_28__2_), .Y(_320_) );
OAI21X1 OAI21X1_6 ( .A(w_cout_4_), .B(_319_), .C(_320_), .Y(_0__22_) );
INVX1 INVX1_6 ( .A(_27__3_), .Y(_321_) );
NAND2X1 NAND2X1_7 ( .A(w_cout_4_), .B(_28__3_), .Y(_322_) );
OAI21X1 OAI21X1_7 ( .A(w_cout_4_), .B(_321_), .C(_322_), .Y(_0__23_) );
INVX1 INVX1_7 ( .A(1'b0), .Y(_326_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_327_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_328_) );
NAND3X1 NAND3X1_2 ( .A(_326_), .B(_328_), .C(_327_), .Y(_329_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_323_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_324_) );
OAI21X1 OAI21X1_8 ( .A(_323_), .B(_324_), .C(1'b0), .Y(_325_) );
NAND2X1 NAND2X1_9 ( .A(_325_), .B(_329_), .Y(_27__0_) );
OAI21X1 OAI21X1_9 ( .A(_326_), .B(_323_), .C(_328_), .Y(_29__1_) );
INVX1 INVX1_8 ( .A(_29__3_), .Y(_333_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_334_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_335_) );
NAND3X1 NAND3X1_3 ( .A(_333_), .B(_335_), .C(_334_), .Y(_336_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_330_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_331_) );
OAI21X1 OAI21X1_10 ( .A(_330_), .B(_331_), .C(_29__3_), .Y(_332_) );
NAND2X1 NAND2X1_11 ( .A(_332_), .B(_336_), .Y(_27__3_) );
OAI21X1 OAI21X1_11 ( .A(_333_), .B(_330_), .C(_335_), .Y(_25_) );
INVX1 INVX1_9 ( .A(_29__1_), .Y(_340_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_341_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_342_) );
NAND3X1 NAND3X1_4 ( .A(_340_), .B(_342_), .C(_341_), .Y(_343_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_337_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_338_) );
OAI21X1 OAI21X1_12 ( .A(_337_), .B(_338_), .C(_29__1_), .Y(_339_) );
NAND2X1 NAND2X1_13 ( .A(_339_), .B(_343_), .Y(_27__1_) );
OAI21X1 OAI21X1_13 ( .A(_340_), .B(_337_), .C(_342_), .Y(_29__2_) );
INVX1 INVX1_10 ( .A(_29__2_), .Y(_347_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_348_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_349_) );
NAND3X1 NAND3X1_5 ( .A(_347_), .B(_349_), .C(_348_), .Y(_350_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_344_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_345_) );
OAI21X1 OAI21X1_14 ( .A(_344_), .B(_345_), .C(_29__2_), .Y(_346_) );
NAND2X1 NAND2X1_15 ( .A(_346_), .B(_350_), .Y(_27__2_) );
OAI21X1 OAI21X1_15 ( .A(_347_), .B(_344_), .C(_349_), .Y(_29__3_) );
INVX1 INVX1_11 ( .A(1'b1), .Y(_354_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_355_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_356_) );
NAND3X1 NAND3X1_6 ( .A(_354_), .B(_356_), .C(_355_), .Y(_357_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_351_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_352_) );
OAI21X1 OAI21X1_16 ( .A(_351_), .B(_352_), .C(1'b1), .Y(_353_) );
NAND2X1 NAND2X1_17 ( .A(_353_), .B(_357_), .Y(_28__0_) );
OAI21X1 OAI21X1_17 ( .A(_354_), .B(_351_), .C(_356_), .Y(_30__1_) );
INVX1 INVX1_12 ( .A(_30__3_), .Y(_361_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_362_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_363_) );
NAND3X1 NAND3X1_7 ( .A(_361_), .B(_363_), .C(_362_), .Y(_364_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_358_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_359_) );
OAI21X1 OAI21X1_18 ( .A(_358_), .B(_359_), .C(_30__3_), .Y(_360_) );
NAND2X1 NAND2X1_19 ( .A(_360_), .B(_364_), .Y(_28__3_) );
OAI21X1 OAI21X1_19 ( .A(_361_), .B(_358_), .C(_363_), .Y(_26_) );
INVX1 INVX1_13 ( .A(_30__1_), .Y(_368_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_369_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_370_) );
NAND3X1 NAND3X1_8 ( .A(_368_), .B(_370_), .C(_369_), .Y(_371_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_365_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_366_) );
OAI21X1 OAI21X1_20 ( .A(_365_), .B(_366_), .C(_30__1_), .Y(_367_) );
NAND2X1 NAND2X1_21 ( .A(_367_), .B(_371_), .Y(_28__1_) );
OAI21X1 OAI21X1_21 ( .A(_368_), .B(_365_), .C(_370_), .Y(_30__2_) );
INVX1 INVX1_14 ( .A(_30__2_), .Y(_375_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_376_) );
NAND2X1 NAND2X1_22 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_377_) );
NAND3X1 NAND3X1_9 ( .A(_375_), .B(_377_), .C(_376_), .Y(_378_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_372_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_373_) );
OAI21X1 OAI21X1_22 ( .A(_372_), .B(_373_), .C(_30__2_), .Y(_374_) );
NAND2X1 NAND2X1_23 ( .A(_374_), .B(_378_), .Y(_28__2_) );
OAI21X1 OAI21X1_23 ( .A(_375_), .B(_372_), .C(_377_), .Y(_30__3_) );
INVX1 INVX1_15 ( .A(_31_), .Y(_379_) );
NAND2X1 NAND2X1_24 ( .A(_32_), .B(w_cout_5_), .Y(_380_) );
OAI21X1 OAI21X1_24 ( .A(w_cout_5_), .B(_379_), .C(_380_), .Y(w_cout_6_) );
INVX1 INVX1_16 ( .A(_33__0_), .Y(_381_) );
NAND2X1 NAND2X1_25 ( .A(_34__0_), .B(w_cout_5_), .Y(_382_) );
OAI21X1 OAI21X1_25 ( .A(w_cout_5_), .B(_381_), .C(_382_), .Y(_0__24_) );
INVX1 INVX1_17 ( .A(_33__1_), .Y(_383_) );
NAND2X1 NAND2X1_26 ( .A(w_cout_5_), .B(_34__1_), .Y(_384_) );
OAI21X1 OAI21X1_26 ( .A(w_cout_5_), .B(_383_), .C(_384_), .Y(_0__25_) );
INVX1 INVX1_18 ( .A(_33__2_), .Y(_385_) );
NAND2X1 NAND2X1_27 ( .A(w_cout_5_), .B(_34__2_), .Y(_386_) );
OAI21X1 OAI21X1_27 ( .A(w_cout_5_), .B(_385_), .C(_386_), .Y(_0__26_) );
INVX1 INVX1_19 ( .A(_33__3_), .Y(_387_) );
NAND2X1 NAND2X1_28 ( .A(w_cout_5_), .B(_34__3_), .Y(_388_) );
OAI21X1 OAI21X1_28 ( .A(w_cout_5_), .B(_387_), .C(_388_), .Y(_0__27_) );
INVX1 INVX1_20 ( .A(1'b0), .Y(_392_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_393_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_394_) );
NAND3X1 NAND3X1_10 ( .A(_392_), .B(_394_), .C(_393_), .Y(_395_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_389_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_390_) );
OAI21X1 OAI21X1_29 ( .A(_389_), .B(_390_), .C(1'b0), .Y(_391_) );
NAND2X1 NAND2X1_30 ( .A(_391_), .B(_395_), .Y(_33__0_) );
OAI21X1 OAI21X1_30 ( .A(_392_), .B(_389_), .C(_394_), .Y(_35__1_) );
INVX1 INVX1_21 ( .A(_35__3_), .Y(_399_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_400_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_401_) );
NAND3X1 NAND3X1_11 ( .A(_399_), .B(_401_), .C(_400_), .Y(_402_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_396_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_397_) );
OAI21X1 OAI21X1_31 ( .A(_396_), .B(_397_), .C(_35__3_), .Y(_398_) );
NAND2X1 NAND2X1_32 ( .A(_398_), .B(_402_), .Y(_33__3_) );
OAI21X1 OAI21X1_32 ( .A(_399_), .B(_396_), .C(_401_), .Y(_31_) );
INVX1 INVX1_22 ( .A(_35__1_), .Y(_406_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_407_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_408_) );
NAND3X1 NAND3X1_12 ( .A(_406_), .B(_408_), .C(_407_), .Y(_409_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_403_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_404_) );
OAI21X1 OAI21X1_33 ( .A(_403_), .B(_404_), .C(_35__1_), .Y(_405_) );
NAND2X1 NAND2X1_34 ( .A(_405_), .B(_409_), .Y(_33__1_) );
OAI21X1 OAI21X1_34 ( .A(_406_), .B(_403_), .C(_408_), .Y(_35__2_) );
INVX1 INVX1_23 ( .A(_35__2_), .Y(_413_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_414_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_415_) );
NAND3X1 NAND3X1_13 ( .A(_413_), .B(_415_), .C(_414_), .Y(_416_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_410_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_411_) );
OAI21X1 OAI21X1_35 ( .A(_410_), .B(_411_), .C(_35__2_), .Y(_412_) );
NAND2X1 NAND2X1_36 ( .A(_412_), .B(_416_), .Y(_33__2_) );
OAI21X1 OAI21X1_36 ( .A(_413_), .B(_410_), .C(_415_), .Y(_35__3_) );
INVX1 INVX1_24 ( .A(1'b1), .Y(_420_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_421_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_422_) );
NAND3X1 NAND3X1_14 ( .A(_420_), .B(_422_), .C(_421_), .Y(_423_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_417_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_418_) );
OAI21X1 OAI21X1_37 ( .A(_417_), .B(_418_), .C(1'b1), .Y(_419_) );
NAND2X1 NAND2X1_38 ( .A(_419_), .B(_423_), .Y(_34__0_) );
OAI21X1 OAI21X1_38 ( .A(_420_), .B(_417_), .C(_422_), .Y(_36__1_) );
INVX1 INVX1_25 ( .A(_36__3_), .Y(_427_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_428_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_429_) );
NAND3X1 NAND3X1_15 ( .A(_427_), .B(_429_), .C(_428_), .Y(_430_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_424_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_425_) );
OAI21X1 OAI21X1_39 ( .A(_424_), .B(_425_), .C(_36__3_), .Y(_426_) );
NAND2X1 NAND2X1_40 ( .A(_426_), .B(_430_), .Y(_34__3_) );
OAI21X1 OAI21X1_40 ( .A(_427_), .B(_424_), .C(_429_), .Y(_32_) );
INVX1 INVX1_26 ( .A(_36__1_), .Y(_434_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_435_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_436_) );
NAND3X1 NAND3X1_16 ( .A(_434_), .B(_436_), .C(_435_), .Y(_437_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_431_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_432_) );
OAI21X1 OAI21X1_41 ( .A(_431_), .B(_432_), .C(_36__1_), .Y(_433_) );
NAND2X1 NAND2X1_42 ( .A(_433_), .B(_437_), .Y(_34__1_) );
OAI21X1 OAI21X1_42 ( .A(_434_), .B(_431_), .C(_436_), .Y(_36__2_) );
INVX1 INVX1_27 ( .A(_36__2_), .Y(_441_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_442_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_443_) );
NAND3X1 NAND3X1_17 ( .A(_441_), .B(_443_), .C(_442_), .Y(_444_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_438_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_439_) );
OAI21X1 OAI21X1_43 ( .A(_438_), .B(_439_), .C(_36__2_), .Y(_440_) );
NAND2X1 NAND2X1_44 ( .A(_440_), .B(_444_), .Y(_34__2_) );
OAI21X1 OAI21X1_44 ( .A(_441_), .B(_438_), .C(_443_), .Y(_36__3_) );
INVX1 INVX1_28 ( .A(_37_), .Y(_445_) );
NAND2X1 NAND2X1_45 ( .A(_38_), .B(w_cout_6_), .Y(_446_) );
OAI21X1 OAI21X1_45 ( .A(w_cout_6_), .B(_445_), .C(_446_), .Y(w_cout_7_) );
INVX1 INVX1_29 ( .A(_39__0_), .Y(_447_) );
NAND2X1 NAND2X1_46 ( .A(_40__0_), .B(w_cout_6_), .Y(_448_) );
OAI21X1 OAI21X1_46 ( .A(w_cout_6_), .B(_447_), .C(_448_), .Y(_0__28_) );
INVX1 INVX1_30 ( .A(_39__1_), .Y(_449_) );
NAND2X1 NAND2X1_47 ( .A(w_cout_6_), .B(_40__1_), .Y(_450_) );
OAI21X1 OAI21X1_47 ( .A(w_cout_6_), .B(_449_), .C(_450_), .Y(_0__29_) );
INVX1 INVX1_31 ( .A(_39__2_), .Y(_451_) );
NAND2X1 NAND2X1_48 ( .A(w_cout_6_), .B(_40__2_), .Y(_452_) );
OAI21X1 OAI21X1_48 ( .A(w_cout_6_), .B(_451_), .C(_452_), .Y(_0__30_) );
INVX1 INVX1_32 ( .A(_39__3_), .Y(_453_) );
NAND2X1 NAND2X1_49 ( .A(w_cout_6_), .B(_40__3_), .Y(_454_) );
OAI21X1 OAI21X1_49 ( .A(w_cout_6_), .B(_453_), .C(_454_), .Y(_0__31_) );
INVX1 INVX1_33 ( .A(1'b0), .Y(_458_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_459_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_460_) );
NAND3X1 NAND3X1_18 ( .A(_458_), .B(_460_), .C(_459_), .Y(_461_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_455_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_456_) );
OAI21X1 OAI21X1_50 ( .A(_455_), .B(_456_), .C(1'b0), .Y(_457_) );
NAND2X1 NAND2X1_51 ( .A(_457_), .B(_461_), .Y(_39__0_) );
OAI21X1 OAI21X1_51 ( .A(_458_), .B(_455_), .C(_460_), .Y(_41__1_) );
INVX1 INVX1_34 ( .A(_41__3_), .Y(_465_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_466_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_467_) );
NAND3X1 NAND3X1_19 ( .A(_465_), .B(_467_), .C(_466_), .Y(_468_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_462_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_463_) );
OAI21X1 OAI21X1_52 ( .A(_462_), .B(_463_), .C(_41__3_), .Y(_464_) );
NAND2X1 NAND2X1_53 ( .A(_464_), .B(_468_), .Y(_39__3_) );
OAI21X1 OAI21X1_53 ( .A(_465_), .B(_462_), .C(_467_), .Y(_37_) );
INVX1 INVX1_35 ( .A(_41__1_), .Y(_472_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_473_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_474_) );
NAND3X1 NAND3X1_20 ( .A(_472_), .B(_474_), .C(_473_), .Y(_475_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_469_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_470_) );
OAI21X1 OAI21X1_54 ( .A(_469_), .B(_470_), .C(_41__1_), .Y(_471_) );
NAND2X1 NAND2X1_55 ( .A(_471_), .B(_475_), .Y(_39__1_) );
OAI21X1 OAI21X1_55 ( .A(_472_), .B(_469_), .C(_474_), .Y(_41__2_) );
INVX1 INVX1_36 ( .A(_41__2_), .Y(_479_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_480_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_481_) );
NAND3X1 NAND3X1_21 ( .A(_479_), .B(_481_), .C(_480_), .Y(_482_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_476_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_477_) );
OAI21X1 OAI21X1_56 ( .A(_476_), .B(_477_), .C(_41__2_), .Y(_478_) );
NAND2X1 NAND2X1_57 ( .A(_478_), .B(_482_), .Y(_39__2_) );
OAI21X1 OAI21X1_57 ( .A(_479_), .B(_476_), .C(_481_), .Y(_41__3_) );
INVX1 INVX1_37 ( .A(1'b1), .Y(_486_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_487_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_488_) );
NAND3X1 NAND3X1_22 ( .A(_486_), .B(_488_), .C(_487_), .Y(_489_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_483_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_484_) );
OAI21X1 OAI21X1_58 ( .A(_483_), .B(_484_), .C(1'b1), .Y(_485_) );
NAND2X1 NAND2X1_59 ( .A(_485_), .B(_489_), .Y(_40__0_) );
OAI21X1 OAI21X1_59 ( .A(_486_), .B(_483_), .C(_488_), .Y(_42__1_) );
INVX1 INVX1_38 ( .A(_42__3_), .Y(_493_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_494_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_495_) );
NAND3X1 NAND3X1_23 ( .A(_493_), .B(_495_), .C(_494_), .Y(_496_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_490_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_491_) );
OAI21X1 OAI21X1_60 ( .A(_490_), .B(_491_), .C(_42__3_), .Y(_492_) );
NAND2X1 NAND2X1_61 ( .A(_492_), .B(_496_), .Y(_40__3_) );
OAI21X1 OAI21X1_61 ( .A(_493_), .B(_490_), .C(_495_), .Y(_38_) );
INVX1 INVX1_39 ( .A(_42__1_), .Y(_500_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_501_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_502_) );
NAND3X1 NAND3X1_24 ( .A(_500_), .B(_502_), .C(_501_), .Y(_503_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_497_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_498_) );
OAI21X1 OAI21X1_62 ( .A(_497_), .B(_498_), .C(_42__1_), .Y(_499_) );
NAND2X1 NAND2X1_63 ( .A(_499_), .B(_503_), .Y(_40__1_) );
OAI21X1 OAI21X1_63 ( .A(_500_), .B(_497_), .C(_502_), .Y(_42__2_) );
INVX1 INVX1_40 ( .A(_42__2_), .Y(_507_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_508_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_509_) );
NAND3X1 NAND3X1_25 ( .A(_507_), .B(_509_), .C(_508_), .Y(_510_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_504_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_505_) );
OAI21X1 OAI21X1_64 ( .A(_504_), .B(_505_), .C(_42__2_), .Y(_506_) );
NAND2X1 NAND2X1_65 ( .A(_506_), .B(_510_), .Y(_40__2_) );
OAI21X1 OAI21X1_65 ( .A(_507_), .B(_504_), .C(_509_), .Y(_42__3_) );
INVX1 INVX1_41 ( .A(_43_), .Y(_511_) );
NAND2X1 NAND2X1_66 ( .A(_44_), .B(w_cout_7_), .Y(_512_) );
OAI21X1 OAI21X1_66 ( .A(w_cout_7_), .B(_511_), .C(_512_), .Y(csa_inst_cin) );
INVX1 INVX1_42 ( .A(_45__0_), .Y(_513_) );
NAND2X1 NAND2X1_67 ( .A(_46__0_), .B(w_cout_7_), .Y(_514_) );
OAI21X1 OAI21X1_67 ( .A(w_cout_7_), .B(_513_), .C(_514_), .Y(_0__32_) );
INVX1 INVX1_43 ( .A(_45__1_), .Y(_515_) );
NAND2X1 NAND2X1_68 ( .A(w_cout_7_), .B(_46__1_), .Y(_516_) );
OAI21X1 OAI21X1_68 ( .A(w_cout_7_), .B(_515_), .C(_516_), .Y(_0__33_) );
INVX1 INVX1_44 ( .A(_45__2_), .Y(_517_) );
NAND2X1 NAND2X1_69 ( .A(w_cout_7_), .B(_46__2_), .Y(_518_) );
OAI21X1 OAI21X1_69 ( .A(w_cout_7_), .B(_517_), .C(_518_), .Y(_0__34_) );
INVX1 INVX1_45 ( .A(_45__3_), .Y(_519_) );
NAND2X1 NAND2X1_70 ( .A(w_cout_7_), .B(_46__3_), .Y(_520_) );
OAI21X1 OAI21X1_70 ( .A(w_cout_7_), .B(_519_), .C(_520_), .Y(_0__35_) );
INVX1 INVX1_46 ( .A(1'b0), .Y(_524_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_525_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_526_) );
NAND3X1 NAND3X1_26 ( .A(_524_), .B(_526_), .C(_525_), .Y(_527_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_521_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_522_) );
OAI21X1 OAI21X1_71 ( .A(_521_), .B(_522_), .C(1'b0), .Y(_523_) );
NAND2X1 NAND2X1_72 ( .A(_523_), .B(_527_), .Y(_45__0_) );
OAI21X1 OAI21X1_72 ( .A(_524_), .B(_521_), .C(_526_), .Y(_47__1_) );
INVX1 INVX1_47 ( .A(_47__3_), .Y(_531_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_532_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_533_) );
NAND3X1 NAND3X1_27 ( .A(_531_), .B(_533_), .C(_532_), .Y(_534_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_528_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_529_) );
OAI21X1 OAI21X1_73 ( .A(_528_), .B(_529_), .C(_47__3_), .Y(_530_) );
NAND2X1 NAND2X1_74 ( .A(_530_), .B(_534_), .Y(_45__3_) );
OAI21X1 OAI21X1_74 ( .A(_531_), .B(_528_), .C(_533_), .Y(_43_) );
INVX1 INVX1_48 ( .A(_47__1_), .Y(_538_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_539_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_540_) );
NAND3X1 NAND3X1_28 ( .A(_538_), .B(_540_), .C(_539_), .Y(_541_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_535_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_536_) );
OAI21X1 OAI21X1_75 ( .A(_535_), .B(_536_), .C(_47__1_), .Y(_537_) );
NAND2X1 NAND2X1_76 ( .A(_537_), .B(_541_), .Y(_45__1_) );
OAI21X1 OAI21X1_76 ( .A(_538_), .B(_535_), .C(_540_), .Y(_47__2_) );
INVX1 INVX1_49 ( .A(_47__2_), .Y(_545_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_546_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_547_) );
NAND3X1 NAND3X1_29 ( .A(_545_), .B(_547_), .C(_546_), .Y(_548_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_542_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_543_) );
OAI21X1 OAI21X1_77 ( .A(_542_), .B(_543_), .C(_47__2_), .Y(_544_) );
NAND2X1 NAND2X1_78 ( .A(_544_), .B(_548_), .Y(_45__2_) );
OAI21X1 OAI21X1_78 ( .A(_545_), .B(_542_), .C(_547_), .Y(_47__3_) );
INVX1 INVX1_50 ( .A(1'b1), .Y(_552_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_553_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_554_) );
NAND3X1 NAND3X1_30 ( .A(_552_), .B(_554_), .C(_553_), .Y(_555_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_549_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_550_) );
OAI21X1 OAI21X1_79 ( .A(_549_), .B(_550_), .C(1'b1), .Y(_551_) );
NAND2X1 NAND2X1_80 ( .A(_551_), .B(_555_), .Y(_46__0_) );
OAI21X1 OAI21X1_80 ( .A(_552_), .B(_549_), .C(_554_), .Y(_48__1_) );
INVX1 INVX1_51 ( .A(_48__3_), .Y(_559_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_560_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_561_) );
NAND3X1 NAND3X1_31 ( .A(_559_), .B(_561_), .C(_560_), .Y(_562_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_556_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_557_) );
OAI21X1 OAI21X1_81 ( .A(_556_), .B(_557_), .C(_48__3_), .Y(_558_) );
NAND2X1 NAND2X1_82 ( .A(_558_), .B(_562_), .Y(_46__3_) );
OAI21X1 OAI21X1_82 ( .A(_559_), .B(_556_), .C(_561_), .Y(_44_) );
INVX1 INVX1_52 ( .A(_48__1_), .Y(_566_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_567_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_568_) );
NAND3X1 NAND3X1_32 ( .A(_566_), .B(_568_), .C(_567_), .Y(_569_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_563_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_564_) );
OAI21X1 OAI21X1_83 ( .A(_563_), .B(_564_), .C(_48__1_), .Y(_565_) );
NAND2X1 NAND2X1_84 ( .A(_565_), .B(_569_), .Y(_46__1_) );
OAI21X1 OAI21X1_84 ( .A(_566_), .B(_563_), .C(_568_), .Y(_48__2_) );
INVX1 INVX1_53 ( .A(_48__2_), .Y(_573_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_574_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_575_) );
NAND3X1 NAND3X1_33 ( .A(_573_), .B(_575_), .C(_574_), .Y(_576_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_570_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_571_) );
OAI21X1 OAI21X1_85 ( .A(_570_), .B(_571_), .C(_48__2_), .Y(_572_) );
NAND2X1 NAND2X1_86 ( .A(_572_), .B(_576_), .Y(_46__2_) );
OAI21X1 OAI21X1_86 ( .A(_573_), .B(_570_), .C(_575_), .Y(_48__3_) );
INVX1 INVX1_54 ( .A(csa_inst_cout0_0), .Y(_577_) );
NAND2X1 NAND2X1_87 ( .A(csa_inst_cout0_1), .B(csa_inst_cin), .Y(_578_) );
OAI21X1 OAI21X1_87 ( .A(csa_inst_cin), .B(_577_), .C(_578_), .Y(w_cout_9_) );
INVX1 INVX1_55 ( .A(csa_inst_mux0_sum_i0), .Y(_579_) );
NAND2X1 NAND2X1_88 ( .A(csa_inst_mux0_sum_i1), .B(csa_inst_cin), .Y(_580_) );
OAI21X1 OAI21X1_88 ( .A(csa_inst_cin), .B(_579_), .C(_580_), .Y(csa_inst_mux0_sum_y) );
INVX1 INVX1_56 ( .A(1'b0), .Y(_584_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_585_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_586_) );
NAND3X1 NAND3X1_34 ( .A(_584_), .B(_586_), .C(_585_), .Y(_587_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_581_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_582_) );
OAI21X1 OAI21X1_89 ( .A(_581_), .B(_582_), .C(1'b0), .Y(_583_) );
NAND2X1 NAND2X1_90 ( .A(_583_), .B(_587_), .Y(csa_inst_mux0_sum_i0) );
OAI21X1 OAI21X1_90 ( .A(_584_), .B(_581_), .C(_586_), .Y(csa_inst_cout0_0) );
INVX1 INVX1_57 ( .A(1'b1), .Y(_591_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_592_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_593_) );
NAND3X1 NAND3X1_35 ( .A(_591_), .B(_593_), .C(_592_), .Y(_594_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_588_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_589_) );
OAI21X1 OAI21X1_91 ( .A(_588_), .B(_589_), .C(1'b1), .Y(_590_) );
NAND2X1 NAND2X1_92 ( .A(_590_), .B(_594_), .Y(csa_inst_mux0_sum_i1) );
OAI21X1 OAI21X1_92 ( .A(_591_), .B(_588_), .C(_593_), .Y(csa_inst_cout0_1) );
INVX1 INVX1_58 ( .A(1'b0), .Y(_598_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_599_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_600_) );
NAND3X1 NAND3X1_36 ( .A(_598_), .B(_600_), .C(_599_), .Y(_601_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_595_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_596_) );
OAI21X1 OAI21X1_93 ( .A(_595_), .B(_596_), .C(1'b0), .Y(_597_) );
NAND2X1 NAND2X1_94 ( .A(_597_), .B(_601_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_94 ( .A(_598_), .B(_595_), .C(_600_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_59 ( .A(rca_inst_fa3_i_carry), .Y(_605_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_606_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_607_) );
NAND3X1 NAND3X1_37 ( .A(_605_), .B(_607_), .C(_606_), .Y(_608_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_602_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_603_) );
OAI21X1 OAI21X1_95 ( .A(_602_), .B(_603_), .C(rca_inst_fa3_i_carry), .Y(_604_) );
NAND2X1 NAND2X1_96 ( .A(_604_), .B(_608_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_96 ( .A(_605_), .B(_602_), .C(_607_), .Y(rca_inst_cout) );
INVX1 INVX1_60 ( .A(rca_inst_fa0_o_carry), .Y(_612_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_613_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_614_) );
NAND3X1 NAND3X1_38 ( .A(_612_), .B(_614_), .C(_613_), .Y(_615_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_609_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_610_) );
OAI21X1 OAI21X1_97 ( .A(_609_), .B(_610_), .C(rca_inst_fa0_o_carry), .Y(_611_) );
NAND2X1 NAND2X1_98 ( .A(_611_), .B(_615_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_98 ( .A(_612_), .B(_609_), .C(_614_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_61 ( .A(rca_inst_fa_1__o_carry), .Y(_619_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_620_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_621_) );
NAND3X1 NAND3X1_39 ( .A(_619_), .B(_621_), .C(_620_), .Y(_622_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_616_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_617_) );
OAI21X1 OAI21X1_99 ( .A(_616_), .B(_617_), .C(rca_inst_fa_1__o_carry), .Y(_618_) );
NAND2X1 NAND2X1_100 ( .A(_618_), .B(_622_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_100 ( .A(_619_), .B(_616_), .C(_621_), .Y(rca_inst_fa3_i_carry) );
BUFX2 BUFX2_1 ( .A(w_cout_9_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(csa_inst_mux0_sum_y), .Y(sum[36]) );
INVX1 INVX1_62 ( .A(_1_), .Y(_49_) );
NAND2X1 NAND2X1_101 ( .A(_2_), .B(rca_inst_cout), .Y(_50_) );
OAI21X1 OAI21X1_101 ( .A(rca_inst_cout), .B(_49_), .C(_50_), .Y(w_cout_1_) );
INVX1 INVX1_63 ( .A(_3__0_), .Y(_51_) );
NAND2X1 NAND2X1_102 ( .A(_4__0_), .B(rca_inst_cout), .Y(_52_) );
OAI21X1 OAI21X1_102 ( .A(rca_inst_cout), .B(_51_), .C(_52_), .Y(_0__4_) );
INVX1 INVX1_64 ( .A(_3__1_), .Y(_53_) );
NAND2X1 NAND2X1_103 ( .A(rca_inst_cout), .B(_4__1_), .Y(_54_) );
OAI21X1 OAI21X1_103 ( .A(rca_inst_cout), .B(_53_), .C(_54_), .Y(_0__5_) );
INVX1 INVX1_65 ( .A(_3__2_), .Y(_55_) );
NAND2X1 NAND2X1_104 ( .A(rca_inst_cout), .B(_4__2_), .Y(_56_) );
OAI21X1 OAI21X1_104 ( .A(rca_inst_cout), .B(_55_), .C(_56_), .Y(_0__6_) );
INVX1 INVX1_66 ( .A(_3__3_), .Y(_57_) );
NAND2X1 NAND2X1_105 ( .A(rca_inst_cout), .B(_4__3_), .Y(_58_) );
OAI21X1 OAI21X1_105 ( .A(rca_inst_cout), .B(_57_), .C(_58_), .Y(_0__7_) );
INVX1 INVX1_67 ( .A(1'b0), .Y(_62_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_63_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_64_) );
NAND3X1 NAND3X1_40 ( .A(_62_), .B(_64_), .C(_63_), .Y(_65_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_59_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_60_) );
OAI21X1 OAI21X1_106 ( .A(_59_), .B(_60_), .C(1'b0), .Y(_61_) );
NAND2X1 NAND2X1_107 ( .A(_61_), .B(_65_), .Y(_3__0_) );
OAI21X1 OAI21X1_107 ( .A(_62_), .B(_59_), .C(_64_), .Y(_5__1_) );
INVX1 INVX1_68 ( .A(_5__3_), .Y(_69_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_70_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_71_) );
NAND3X1 NAND3X1_41 ( .A(_69_), .B(_71_), .C(_70_), .Y(_72_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_66_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_67_) );
OAI21X1 OAI21X1_108 ( .A(_66_), .B(_67_), .C(_5__3_), .Y(_68_) );
NAND2X1 NAND2X1_109 ( .A(_68_), .B(_72_), .Y(_3__3_) );
OAI21X1 OAI21X1_109 ( .A(_69_), .B(_66_), .C(_71_), .Y(_1_) );
INVX1 INVX1_69 ( .A(_5__1_), .Y(_76_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_77_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_78_) );
NAND3X1 NAND3X1_42 ( .A(_76_), .B(_78_), .C(_77_), .Y(_79_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_73_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_74_) );
OAI21X1 OAI21X1_110 ( .A(_73_), .B(_74_), .C(_5__1_), .Y(_75_) );
NAND2X1 NAND2X1_111 ( .A(_75_), .B(_79_), .Y(_3__1_) );
OAI21X1 OAI21X1_111 ( .A(_76_), .B(_73_), .C(_78_), .Y(_5__2_) );
INVX1 INVX1_70 ( .A(_5__2_), .Y(_83_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_84_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_85_) );
NAND3X1 NAND3X1_43 ( .A(_83_), .B(_85_), .C(_84_), .Y(_86_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_80_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_81_) );
OAI21X1 OAI21X1_112 ( .A(_80_), .B(_81_), .C(_5__2_), .Y(_82_) );
NAND2X1 NAND2X1_113 ( .A(_82_), .B(_86_), .Y(_3__2_) );
OAI21X1 OAI21X1_113 ( .A(_83_), .B(_80_), .C(_85_), .Y(_5__3_) );
INVX1 INVX1_71 ( .A(1'b1), .Y(_90_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_91_) );
NAND2X1 NAND2X1_114 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_92_) );
NAND3X1 NAND3X1_44 ( .A(_90_), .B(_92_), .C(_91_), .Y(_93_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_87_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_88_) );
OAI21X1 OAI21X1_114 ( .A(_87_), .B(_88_), .C(1'b1), .Y(_89_) );
NAND2X1 NAND2X1_115 ( .A(_89_), .B(_93_), .Y(_4__0_) );
OAI21X1 OAI21X1_115 ( .A(_90_), .B(_87_), .C(_92_), .Y(_6__1_) );
INVX1 INVX1_72 ( .A(_6__3_), .Y(_97_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_98_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_99_) );
NAND3X1 NAND3X1_45 ( .A(_97_), .B(_99_), .C(_98_), .Y(_100_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_94_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_95_) );
OAI21X1 OAI21X1_116 ( .A(_94_), .B(_95_), .C(_6__3_), .Y(_96_) );
NAND2X1 NAND2X1_117 ( .A(_96_), .B(_100_), .Y(_4__3_) );
OAI21X1 OAI21X1_117 ( .A(_97_), .B(_94_), .C(_99_), .Y(_2_) );
INVX1 INVX1_73 ( .A(_6__1_), .Y(_104_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_105_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_106_) );
NAND3X1 NAND3X1_46 ( .A(_104_), .B(_106_), .C(_105_), .Y(_107_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_101_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_102_) );
OAI21X1 OAI21X1_118 ( .A(_101_), .B(_102_), .C(_6__1_), .Y(_103_) );
NAND2X1 NAND2X1_119 ( .A(_103_), .B(_107_), .Y(_4__1_) );
OAI21X1 OAI21X1_119 ( .A(_104_), .B(_101_), .C(_106_), .Y(_6__2_) );
INVX1 INVX1_74 ( .A(_6__2_), .Y(_111_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_112_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_113_) );
NAND3X1 NAND3X1_47 ( .A(_111_), .B(_113_), .C(_112_), .Y(_114_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_108_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_109_) );
OAI21X1 OAI21X1_120 ( .A(_108_), .B(_109_), .C(_6__2_), .Y(_110_) );
NAND2X1 NAND2X1_121 ( .A(_110_), .B(_114_), .Y(_4__2_) );
OAI21X1 OAI21X1_121 ( .A(_111_), .B(_108_), .C(_113_), .Y(_6__3_) );
INVX1 INVX1_75 ( .A(_7_), .Y(_115_) );
NAND2X1 NAND2X1_122 ( .A(_8_), .B(w_cout_1_), .Y(_116_) );
OAI21X1 OAI21X1_122 ( .A(w_cout_1_), .B(_115_), .C(_116_), .Y(w_cout_2_) );
INVX1 INVX1_76 ( .A(_9__0_), .Y(_117_) );
NAND2X1 NAND2X1_123 ( .A(_10__0_), .B(w_cout_1_), .Y(_118_) );
OAI21X1 OAI21X1_123 ( .A(w_cout_1_), .B(_117_), .C(_118_), .Y(_0__8_) );
INVX1 INVX1_77 ( .A(_9__1_), .Y(_119_) );
NAND2X1 NAND2X1_124 ( .A(w_cout_1_), .B(_10__1_), .Y(_120_) );
OAI21X1 OAI21X1_124 ( .A(w_cout_1_), .B(_119_), .C(_120_), .Y(_0__9_) );
INVX1 INVX1_78 ( .A(_9__2_), .Y(_121_) );
NAND2X1 NAND2X1_125 ( .A(w_cout_1_), .B(_10__2_), .Y(_122_) );
OAI21X1 OAI21X1_125 ( .A(w_cout_1_), .B(_121_), .C(_122_), .Y(_0__10_) );
INVX1 INVX1_79 ( .A(_9__3_), .Y(_123_) );
NAND2X1 NAND2X1_126 ( .A(w_cout_1_), .B(_10__3_), .Y(_124_) );
OAI21X1 OAI21X1_126 ( .A(w_cout_1_), .B(_123_), .C(_124_), .Y(_0__11_) );
INVX1 INVX1_80 ( .A(1'b0), .Y(_128_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_129_) );
NAND2X1 NAND2X1_127 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_130_) );
NAND3X1 NAND3X1_48 ( .A(_128_), .B(_130_), .C(_129_), .Y(_131_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_125_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_126_) );
OAI21X1 OAI21X1_127 ( .A(_125_), .B(_126_), .C(1'b0), .Y(_127_) );
NAND2X1 NAND2X1_128 ( .A(_127_), .B(_131_), .Y(_9__0_) );
OAI21X1 OAI21X1_128 ( .A(_128_), .B(_125_), .C(_130_), .Y(_11__1_) );
INVX1 INVX1_81 ( .A(_11__3_), .Y(_135_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_136_) );
NAND2X1 NAND2X1_129 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_137_) );
NAND3X1 NAND3X1_49 ( .A(_135_), .B(_137_), .C(_136_), .Y(_138_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_132_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_133_) );
OAI21X1 OAI21X1_129 ( .A(_132_), .B(_133_), .C(_11__3_), .Y(_134_) );
NAND2X1 NAND2X1_130 ( .A(_134_), .B(_138_), .Y(_9__3_) );
OAI21X1 OAI21X1_130 ( .A(_135_), .B(_132_), .C(_137_), .Y(_7_) );
INVX1 INVX1_82 ( .A(_11__1_), .Y(_142_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_143_) );
NAND2X1 NAND2X1_131 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_144_) );
NAND3X1 NAND3X1_50 ( .A(_142_), .B(_144_), .C(_143_), .Y(_145_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_139_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_140_) );
OAI21X1 OAI21X1_131 ( .A(_139_), .B(_140_), .C(_11__1_), .Y(_141_) );
NAND2X1 NAND2X1_132 ( .A(_141_), .B(_145_), .Y(_9__1_) );
OAI21X1 OAI21X1_132 ( .A(_142_), .B(_139_), .C(_144_), .Y(_11__2_) );
INVX1 INVX1_83 ( .A(_11__2_), .Y(_149_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_150_) );
NAND2X1 NAND2X1_133 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_151_) );
NAND3X1 NAND3X1_51 ( .A(_149_), .B(_151_), .C(_150_), .Y(_152_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_146_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_147_) );
OAI21X1 OAI21X1_133 ( .A(_146_), .B(_147_), .C(_11__2_), .Y(_148_) );
NAND2X1 NAND2X1_134 ( .A(_148_), .B(_152_), .Y(_9__2_) );
OAI21X1 OAI21X1_134 ( .A(_149_), .B(_146_), .C(_151_), .Y(_11__3_) );
INVX1 INVX1_84 ( .A(1'b1), .Y(_156_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_157_) );
NAND2X1 NAND2X1_135 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_158_) );
NAND3X1 NAND3X1_52 ( .A(_156_), .B(_158_), .C(_157_), .Y(_159_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_153_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_154_) );
OAI21X1 OAI21X1_135 ( .A(_153_), .B(_154_), .C(1'b1), .Y(_155_) );
NAND2X1 NAND2X1_136 ( .A(_155_), .B(_159_), .Y(_10__0_) );
OAI21X1 OAI21X1_136 ( .A(_156_), .B(_153_), .C(_158_), .Y(_12__1_) );
INVX1 INVX1_85 ( .A(_12__3_), .Y(_163_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_164_) );
NAND2X1 NAND2X1_137 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_165_) );
NAND3X1 NAND3X1_53 ( .A(_163_), .B(_165_), .C(_164_), .Y(_166_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_160_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_161_) );
OAI21X1 OAI21X1_137 ( .A(_160_), .B(_161_), .C(_12__3_), .Y(_162_) );
NAND2X1 NAND2X1_138 ( .A(_162_), .B(_166_), .Y(_10__3_) );
OAI21X1 OAI21X1_138 ( .A(_163_), .B(_160_), .C(_165_), .Y(_8_) );
INVX1 INVX1_86 ( .A(_12__1_), .Y(_170_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_171_) );
NAND2X1 NAND2X1_139 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_172_) );
NAND3X1 NAND3X1_54 ( .A(_170_), .B(_172_), .C(_171_), .Y(_173_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_167_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_168_) );
OAI21X1 OAI21X1_139 ( .A(_167_), .B(_168_), .C(_12__1_), .Y(_169_) );
NAND2X1 NAND2X1_140 ( .A(_169_), .B(_173_), .Y(_10__1_) );
OAI21X1 OAI21X1_140 ( .A(_170_), .B(_167_), .C(_172_), .Y(_12__2_) );
INVX1 INVX1_87 ( .A(_12__2_), .Y(_177_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_178_) );
NAND2X1 NAND2X1_141 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_179_) );
NAND3X1 NAND3X1_55 ( .A(_177_), .B(_179_), .C(_178_), .Y(_180_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_174_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_175_) );
OAI21X1 OAI21X1_141 ( .A(_174_), .B(_175_), .C(_12__2_), .Y(_176_) );
NAND2X1 NAND2X1_142 ( .A(_176_), .B(_180_), .Y(_10__2_) );
OAI21X1 OAI21X1_142 ( .A(_177_), .B(_174_), .C(_179_), .Y(_12__3_) );
INVX1 INVX1_88 ( .A(_13_), .Y(_181_) );
NAND2X1 NAND2X1_143 ( .A(_14_), .B(w_cout_2_), .Y(_182_) );
OAI21X1 OAI21X1_143 ( .A(w_cout_2_), .B(_181_), .C(_182_), .Y(w_cout_3_) );
INVX1 INVX1_89 ( .A(_15__0_), .Y(_183_) );
NAND2X1 NAND2X1_144 ( .A(_16__0_), .B(w_cout_2_), .Y(_184_) );
OAI21X1 OAI21X1_144 ( .A(w_cout_2_), .B(_183_), .C(_184_), .Y(_0__12_) );
INVX1 INVX1_90 ( .A(_15__1_), .Y(_185_) );
NAND2X1 NAND2X1_145 ( .A(w_cout_2_), .B(_16__1_), .Y(_186_) );
OAI21X1 OAI21X1_145 ( .A(w_cout_2_), .B(_185_), .C(_186_), .Y(_0__13_) );
INVX1 INVX1_91 ( .A(_15__2_), .Y(_187_) );
NAND2X1 NAND2X1_146 ( .A(w_cout_2_), .B(_16__2_), .Y(_188_) );
OAI21X1 OAI21X1_146 ( .A(w_cout_2_), .B(_187_), .C(_188_), .Y(_0__14_) );
INVX1 INVX1_92 ( .A(_15__3_), .Y(_189_) );
NAND2X1 NAND2X1_147 ( .A(w_cout_2_), .B(_16__3_), .Y(_190_) );
OAI21X1 OAI21X1_147 ( .A(w_cout_2_), .B(_189_), .C(_190_), .Y(_0__15_) );
INVX1 INVX1_93 ( .A(1'b0), .Y(_194_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_195_) );
NAND2X1 NAND2X1_148 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_196_) );
NAND3X1 NAND3X1_56 ( .A(_194_), .B(_196_), .C(_195_), .Y(_197_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_191_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_192_) );
OAI21X1 OAI21X1_148 ( .A(_191_), .B(_192_), .C(1'b0), .Y(_193_) );
NAND2X1 NAND2X1_149 ( .A(_193_), .B(_197_), .Y(_15__0_) );
OAI21X1 OAI21X1_149 ( .A(_194_), .B(_191_), .C(_196_), .Y(_17__1_) );
INVX1 INVX1_94 ( .A(_17__3_), .Y(_201_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_202_) );
NAND2X1 NAND2X1_150 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_203_) );
NAND3X1 NAND3X1_57 ( .A(_201_), .B(_203_), .C(_202_), .Y(_204_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_198_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_199_) );
OAI21X1 OAI21X1_150 ( .A(_198_), .B(_199_), .C(_17__3_), .Y(_200_) );
NAND2X1 NAND2X1_151 ( .A(_200_), .B(_204_), .Y(_15__3_) );
OAI21X1 OAI21X1_151 ( .A(_201_), .B(_198_), .C(_203_), .Y(_13_) );
INVX1 INVX1_95 ( .A(_17__1_), .Y(_208_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_209_) );
NAND2X1 NAND2X1_152 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_210_) );
NAND3X1 NAND3X1_58 ( .A(_208_), .B(_210_), .C(_209_), .Y(_211_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_205_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_206_) );
OAI21X1 OAI21X1_152 ( .A(_205_), .B(_206_), .C(_17__1_), .Y(_207_) );
NAND2X1 NAND2X1_153 ( .A(_207_), .B(_211_), .Y(_15__1_) );
OAI21X1 OAI21X1_153 ( .A(_208_), .B(_205_), .C(_210_), .Y(_17__2_) );
INVX1 INVX1_96 ( .A(_17__2_), .Y(_215_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_216_) );
NAND2X1 NAND2X1_154 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_217_) );
NAND3X1 NAND3X1_59 ( .A(_215_), .B(_217_), .C(_216_), .Y(_218_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_212_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_213_) );
OAI21X1 OAI21X1_154 ( .A(_212_), .B(_213_), .C(_17__2_), .Y(_214_) );
NAND2X1 NAND2X1_155 ( .A(_214_), .B(_218_), .Y(_15__2_) );
OAI21X1 OAI21X1_155 ( .A(_215_), .B(_212_), .C(_217_), .Y(_17__3_) );
INVX1 INVX1_97 ( .A(1'b1), .Y(_222_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_223_) );
NAND2X1 NAND2X1_156 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_224_) );
NAND3X1 NAND3X1_60 ( .A(_222_), .B(_224_), .C(_223_), .Y(_225_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_219_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_220_) );
OAI21X1 OAI21X1_156 ( .A(_219_), .B(_220_), .C(1'b1), .Y(_221_) );
NAND2X1 NAND2X1_157 ( .A(_221_), .B(_225_), .Y(_16__0_) );
OAI21X1 OAI21X1_157 ( .A(_222_), .B(_219_), .C(_224_), .Y(_18__1_) );
INVX1 INVX1_98 ( .A(_18__3_), .Y(_229_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_230_) );
NAND2X1 NAND2X1_158 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_231_) );
NAND3X1 NAND3X1_61 ( .A(_229_), .B(_231_), .C(_230_), .Y(_232_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_226_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_227_) );
OAI21X1 OAI21X1_158 ( .A(_226_), .B(_227_), .C(_18__3_), .Y(_228_) );
NAND2X1 NAND2X1_159 ( .A(_228_), .B(_232_), .Y(_16__3_) );
OAI21X1 OAI21X1_159 ( .A(_229_), .B(_226_), .C(_231_), .Y(_14_) );
INVX1 INVX1_99 ( .A(_18__1_), .Y(_236_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_237_) );
NAND2X1 NAND2X1_160 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_238_) );
NAND3X1 NAND3X1_62 ( .A(_236_), .B(_238_), .C(_237_), .Y(_239_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_233_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_234_) );
OAI21X1 OAI21X1_160 ( .A(_233_), .B(_234_), .C(_18__1_), .Y(_235_) );
NAND2X1 NAND2X1_161 ( .A(_235_), .B(_239_), .Y(_16__1_) );
OAI21X1 OAI21X1_161 ( .A(_236_), .B(_233_), .C(_238_), .Y(_18__2_) );
INVX1 INVX1_100 ( .A(_18__2_), .Y(_243_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_244_) );
NAND2X1 NAND2X1_162 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_245_) );
NAND3X1 NAND3X1_63 ( .A(_243_), .B(_245_), .C(_244_), .Y(_246_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_240_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_241_) );
OAI21X1 OAI21X1_162 ( .A(_240_), .B(_241_), .C(_18__2_), .Y(_242_) );
NAND2X1 NAND2X1_163 ( .A(_242_), .B(_246_), .Y(_16__2_) );
OAI21X1 OAI21X1_163 ( .A(_243_), .B(_240_), .C(_245_), .Y(_18__3_) );
INVX1 INVX1_101 ( .A(_19_), .Y(_247_) );
NAND2X1 NAND2X1_164 ( .A(_20_), .B(w_cout_3_), .Y(_248_) );
OAI21X1 OAI21X1_164 ( .A(w_cout_3_), .B(_247_), .C(_248_), .Y(w_cout_4_) );
INVX1 INVX1_102 ( .A(_21__0_), .Y(_249_) );
NAND2X1 NAND2X1_165 ( .A(_22__0_), .B(w_cout_3_), .Y(_250_) );
OAI21X1 OAI21X1_165 ( .A(w_cout_3_), .B(_249_), .C(_250_), .Y(_0__16_) );
INVX1 INVX1_103 ( .A(_21__1_), .Y(_251_) );
NAND2X1 NAND2X1_166 ( .A(w_cout_3_), .B(_22__1_), .Y(_252_) );
OAI21X1 OAI21X1_166 ( .A(w_cout_3_), .B(_251_), .C(_252_), .Y(_0__17_) );
INVX1 INVX1_104 ( .A(_21__2_), .Y(_253_) );
NAND2X1 NAND2X1_167 ( .A(w_cout_3_), .B(_22__2_), .Y(_254_) );
OAI21X1 OAI21X1_167 ( .A(w_cout_3_), .B(_253_), .C(_254_), .Y(_0__18_) );
INVX1 INVX1_105 ( .A(_21__3_), .Y(_255_) );
NAND2X1 NAND2X1_168 ( .A(w_cout_3_), .B(_22__3_), .Y(_256_) );
OAI21X1 OAI21X1_168 ( .A(w_cout_3_), .B(_255_), .C(_256_), .Y(_0__19_) );
INVX1 INVX1_106 ( .A(1'b0), .Y(_260_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_261_) );
NAND2X1 NAND2X1_169 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_262_) );
NAND3X1 NAND3X1_64 ( .A(_260_), .B(_262_), .C(_261_), .Y(_263_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_257_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_258_) );
OAI21X1 OAI21X1_169 ( .A(_257_), .B(_258_), .C(1'b0), .Y(_259_) );
NAND2X1 NAND2X1_170 ( .A(_259_), .B(_263_), .Y(_21__0_) );
OAI21X1 OAI21X1_170 ( .A(_260_), .B(_257_), .C(_262_), .Y(_23__1_) );
INVX1 INVX1_107 ( .A(_23__3_), .Y(_267_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_268_) );
NAND2X1 NAND2X1_171 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_269_) );
NAND3X1 NAND3X1_65 ( .A(_267_), .B(_269_), .C(_268_), .Y(_270_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_264_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_265_) );
OAI21X1 OAI21X1_171 ( .A(_264_), .B(_265_), .C(_23__3_), .Y(_266_) );
NAND2X1 NAND2X1_172 ( .A(_266_), .B(_270_), .Y(_21__3_) );
OAI21X1 OAI21X1_172 ( .A(_267_), .B(_264_), .C(_269_), .Y(_19_) );
INVX1 INVX1_108 ( .A(_23__1_), .Y(_274_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_275_) );
NAND2X1 NAND2X1_173 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_276_) );
NAND3X1 NAND3X1_66 ( .A(_274_), .B(_276_), .C(_275_), .Y(_277_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_271_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_272_) );
OAI21X1 OAI21X1_173 ( .A(_271_), .B(_272_), .C(_23__1_), .Y(_273_) );
NAND2X1 NAND2X1_174 ( .A(_273_), .B(_277_), .Y(_21__1_) );
OAI21X1 OAI21X1_174 ( .A(_274_), .B(_271_), .C(_276_), .Y(_23__2_) );
INVX1 INVX1_109 ( .A(_23__2_), .Y(_281_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_282_) );
NAND2X1 NAND2X1_175 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_283_) );
NAND3X1 NAND3X1_67 ( .A(_281_), .B(_283_), .C(_282_), .Y(_284_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_278_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_279_) );
OAI21X1 OAI21X1_175 ( .A(_278_), .B(_279_), .C(_23__2_), .Y(_280_) );
NAND2X1 NAND2X1_176 ( .A(_280_), .B(_284_), .Y(_21__2_) );
OAI21X1 OAI21X1_176 ( .A(_281_), .B(_278_), .C(_283_), .Y(_23__3_) );
INVX1 INVX1_110 ( .A(1'b1), .Y(_288_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_289_) );
NAND2X1 NAND2X1_177 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_290_) );
NAND3X1 NAND3X1_68 ( .A(_288_), .B(_290_), .C(_289_), .Y(_291_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_285_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_286_) );
OAI21X1 OAI21X1_177 ( .A(_285_), .B(_286_), .C(1'b1), .Y(_287_) );
NAND2X1 NAND2X1_178 ( .A(_287_), .B(_291_), .Y(_22__0_) );
OAI21X1 OAI21X1_178 ( .A(_288_), .B(_285_), .C(_290_), .Y(_24__1_) );
INVX1 INVX1_111 ( .A(_24__3_), .Y(_295_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_296_) );
NAND2X1 NAND2X1_179 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_297_) );
NAND3X1 NAND3X1_69 ( .A(_295_), .B(_297_), .C(_296_), .Y(_298_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_292_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_293_) );
OAI21X1 OAI21X1_179 ( .A(_292_), .B(_293_), .C(_24__3_), .Y(_294_) );
NAND2X1 NAND2X1_180 ( .A(_294_), .B(_298_), .Y(_22__3_) );
OAI21X1 OAI21X1_180 ( .A(_295_), .B(_292_), .C(_297_), .Y(_20_) );
INVX1 INVX1_112 ( .A(_24__1_), .Y(_302_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_303_) );
NAND2X1 NAND2X1_181 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_304_) );
NAND3X1 NAND3X1_70 ( .A(_302_), .B(_304_), .C(_303_), .Y(_305_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_299_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_300_) );
OAI21X1 OAI21X1_181 ( .A(_299_), .B(_300_), .C(_24__1_), .Y(_301_) );
NAND2X1 NAND2X1_182 ( .A(_301_), .B(_305_), .Y(_22__1_) );
OAI21X1 OAI21X1_182 ( .A(_302_), .B(_299_), .C(_304_), .Y(_24__2_) );
BUFX2 BUFX2_39 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_40 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_41 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_42 ( .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_43 ( .A(csa_inst_mux0_sum_y), .Y(_0__36_) );
BUFX2 BUFX2_44 ( .A(rca_inst_cout), .Y(w_cout_0_) );
BUFX2 BUFX2_45 ( .A(csa_inst_cin), .Y(w_cout_8_) );
endmodule
