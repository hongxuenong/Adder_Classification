module cla_18bit (i_add1, i_add2, o_result);

input [17:0] i_add1;
input [17:0] i_add2;
output [18:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_49_) );
INVX1 INVX1_1 ( .A(_49_), .Y(w_C_1_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_50_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_51_) );
NOR2X1 NOR2X1_2 ( .A(_50_), .B(_51_), .Y(w_C_2_) );
INVX1 INVX1_2 ( .A(i_add2[2]), .Y(_52_) );
INVX1 INVX1_3 ( .A(i_add1[2]), .Y(_53_) );
NAND2X1 NAND2X1_2 ( .A(_52_), .B(_53_), .Y(_54_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_55_) );
OAI21X1 OAI21X1_1 ( .A(_50_), .B(_51_), .C(_55_), .Y(_56_) );
AND2X2 AND2X2_1 ( .A(_56_), .B(_54_), .Y(w_C_3_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_57_) );
OR2X2 OR2X2_1 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_58_) );
NAND3X1 NAND3X1_1 ( .A(_54_), .B(_58_), .C(_56_), .Y(_59_) );
NAND2X1 NAND2X1_5 ( .A(_57_), .B(_59_), .Y(w_C_4_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_60_) );
NAND3X1 NAND3X1_2 ( .A(_57_), .B(_60_), .C(_59_), .Y(_61_) );
OAI21X1 OAI21X1_2 ( .A(i_add2[4]), .B(i_add1[4]), .C(_61_), .Y(_62_) );
INVX1 INVX1_4 ( .A(_62_), .Y(w_C_5_) );
INVX1 INVX1_5 ( .A(i_add2[5]), .Y(_63_) );
INVX1 INVX1_6 ( .A(i_add1[5]), .Y(_64_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_65_) );
INVX1 INVX1_7 ( .A(_65_), .Y(_66_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_67_) );
INVX1 INVX1_8 ( .A(_67_), .Y(_68_) );
NAND3X1 NAND3X1_3 ( .A(_66_), .B(_68_), .C(_61_), .Y(_69_) );
OAI21X1 OAI21X1_3 ( .A(_63_), .B(_64_), .C(_69_), .Y(w_C_6_) );
NOR2X1 NOR2X1_5 ( .A(_63_), .B(_64_), .Y(_70_) );
INVX1 INVX1_9 ( .A(_70_), .Y(_71_) );
AND2X2 AND2X2_2 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_72_) );
INVX1 INVX1_10 ( .A(_72_), .Y(_73_) );
NAND3X1 NAND3X1_4 ( .A(_71_), .B(_73_), .C(_69_), .Y(_74_) );
OAI21X1 OAI21X1_4 ( .A(i_add2[6]), .B(i_add1[6]), .C(_74_), .Y(_75_) );
INVX1 INVX1_11 ( .A(_75_), .Y(w_C_7_) );
INVX1 INVX1_12 ( .A(i_add2[7]), .Y(_76_) );
INVX1 INVX1_13 ( .A(i_add1[7]), .Y(_77_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_78_) );
INVX1 INVX1_14 ( .A(_78_), .Y(_79_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_80_) );
INVX1 INVX1_15 ( .A(_80_), .Y(_81_) );
NAND3X1 NAND3X1_5 ( .A(_79_), .B(_81_), .C(_74_), .Y(_82_) );
OAI21X1 OAI21X1_5 ( .A(_76_), .B(_77_), .C(_82_), .Y(w_C_8_) );
NOR2X1 NOR2X1_8 ( .A(_76_), .B(_77_), .Y(_83_) );
INVX1 INVX1_16 ( .A(_83_), .Y(_84_) );
AND2X2 AND2X2_3 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_85_) );
INVX1 INVX1_17 ( .A(_85_), .Y(_0_) );
NAND3X1 NAND3X1_6 ( .A(_84_), .B(_0_), .C(_82_), .Y(_1_) );
OAI21X1 OAI21X1_6 ( .A(i_add2[8]), .B(i_add1[8]), .C(_1_), .Y(_2_) );
INVX1 INVX1_18 ( .A(_2_), .Y(w_C_9_) );
INVX1 INVX1_19 ( .A(i_add2[9]), .Y(_3_) );
INVX1 INVX1_20 ( .A(i_add1[9]), .Y(_4_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_5_) );
INVX1 INVX1_21 ( .A(_5_), .Y(_6_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_7_) );
INVX1 INVX1_22 ( .A(_7_), .Y(_8_) );
NAND3X1 NAND3X1_7 ( .A(_6_), .B(_8_), .C(_1_), .Y(_9_) );
OAI21X1 OAI21X1_7 ( .A(_3_), .B(_4_), .C(_9_), .Y(w_C_10_) );
NOR2X1 NOR2X1_11 ( .A(_3_), .B(_4_), .Y(_10_) );
INVX1 INVX1_23 ( .A(_10_), .Y(_11_) );
AND2X2 AND2X2_4 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_12_) );
INVX1 INVX1_24 ( .A(_12_), .Y(_13_) );
NAND3X1 NAND3X1_8 ( .A(_11_), .B(_13_), .C(_9_), .Y(_14_) );
OAI21X1 OAI21X1_8 ( .A(i_add2[10]), .B(i_add1[10]), .C(_14_), .Y(_15_) );
INVX1 INVX1_25 ( .A(_15_), .Y(w_C_11_) );
INVX1 INVX1_26 ( .A(i_add2[11]), .Y(_16_) );
INVX1 INVX1_27 ( .A(i_add1[11]), .Y(_17_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_18_) );
INVX1 INVX1_28 ( .A(_18_), .Y(_19_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_20_) );
INVX1 INVX1_29 ( .A(_20_), .Y(_21_) );
NAND3X1 NAND3X1_9 ( .A(_19_), .B(_21_), .C(_14_), .Y(_22_) );
OAI21X1 OAI21X1_9 ( .A(_16_), .B(_17_), .C(_22_), .Y(w_C_12_) );
NOR2X1 NOR2X1_14 ( .A(_16_), .B(_17_), .Y(_23_) );
INVX1 INVX1_30 ( .A(_23_), .Y(_24_) );
AND2X2 AND2X2_5 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_25_) );
INVX1 INVX1_31 ( .A(_25_), .Y(_26_) );
NAND3X1 NAND3X1_10 ( .A(_24_), .B(_26_), .C(_22_), .Y(_27_) );
OAI21X1 OAI21X1_10 ( .A(i_add2[12]), .B(i_add1[12]), .C(_27_), .Y(_28_) );
INVX1 INVX1_32 ( .A(_28_), .Y(w_C_13_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_29_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_30_) );
OAI21X1 OAI21X1_11 ( .A(_30_), .B(_28_), .C(_29_), .Y(w_C_14_) );
OR2X2 OR2X2_2 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_31_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_32_) );
INVX1 INVX1_33 ( .A(_32_), .Y(_33_) );
INVX1 INVX1_34 ( .A(_30_), .Y(_34_) );
NAND3X1 NAND3X1_11 ( .A(_33_), .B(_34_), .C(_27_), .Y(_35_) );
NAND2X1 NAND2X1_8 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_36_) );
NAND3X1 NAND3X1_12 ( .A(_29_), .B(_36_), .C(_35_), .Y(_37_) );
AND2X2 AND2X2_6 ( .A(_37_), .B(_31_), .Y(w_C_15_) );
INVX1 INVX1_35 ( .A(i_add2[15]), .Y(_38_) );
INVX1 INVX1_36 ( .A(i_add1[15]), .Y(_39_) );
NAND2X1 NAND2X1_9 ( .A(_38_), .B(_39_), .Y(_40_) );
NAND3X1 NAND3X1_13 ( .A(_31_), .B(_40_), .C(_37_), .Y(_41_) );
OAI21X1 OAI21X1_12 ( .A(_38_), .B(_39_), .C(_41_), .Y(w_C_16_) );
OR2X2 OR2X2_3 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_42_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_43_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_44_) );
NAND3X1 NAND3X1_14 ( .A(_43_), .B(_44_), .C(_41_), .Y(_45_) );
AND2X2 AND2X2_7 ( .A(_45_), .B(_42_), .Y(w_C_17_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_46_) );
OR2X2 OR2X2_4 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_47_) );
NAND3X1 NAND3X1_15 ( .A(_42_), .B(_47_), .C(_45_), .Y(_48_) );
NAND2X1 NAND2X1_13 ( .A(_46_), .B(_48_), .Y(w_C_18_) );
BUFX2 BUFX2_1 ( .A(_86__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_86__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_86__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_86__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_86__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_86__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_86__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_86__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_86__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_86__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_86__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_86__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_86__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_86__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_86__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_86__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_86__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_86__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(w_C_18_), .Y(o_result[18]) );
INVX1 INVX1_37 ( .A(w_C_4_), .Y(_90_) );
OR2X2 OR2X2_5 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_91_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_92_) );
NAND3X1 NAND3X1_16 ( .A(_90_), .B(_92_), .C(_91_), .Y(_93_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_87_) );
AND2X2 AND2X2_8 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_88_) );
OAI21X1 OAI21X1_13 ( .A(_87_), .B(_88_), .C(w_C_4_), .Y(_89_) );
NAND2X1 NAND2X1_15 ( .A(_89_), .B(_93_), .Y(_86__4_) );
INVX1 INVX1_38 ( .A(w_C_5_), .Y(_97_) );
OR2X2 OR2X2_6 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_98_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_99_) );
NAND3X1 NAND3X1_17 ( .A(_97_), .B(_99_), .C(_98_), .Y(_100_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_94_) );
AND2X2 AND2X2_9 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_95_) );
OAI21X1 OAI21X1_14 ( .A(_94_), .B(_95_), .C(w_C_5_), .Y(_96_) );
NAND2X1 NAND2X1_17 ( .A(_96_), .B(_100_), .Y(_86__5_) );
INVX1 INVX1_39 ( .A(w_C_6_), .Y(_104_) );
OR2X2 OR2X2_7 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_105_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_106_) );
NAND3X1 NAND3X1_18 ( .A(_104_), .B(_106_), .C(_105_), .Y(_107_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_101_) );
AND2X2 AND2X2_10 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_102_) );
OAI21X1 OAI21X1_15 ( .A(_101_), .B(_102_), .C(w_C_6_), .Y(_103_) );
NAND2X1 NAND2X1_19 ( .A(_103_), .B(_107_), .Y(_86__6_) );
INVX1 INVX1_40 ( .A(w_C_7_), .Y(_111_) );
OR2X2 OR2X2_8 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_112_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_113_) );
NAND3X1 NAND3X1_19 ( .A(_111_), .B(_113_), .C(_112_), .Y(_114_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_108_) );
AND2X2 AND2X2_11 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_109_) );
OAI21X1 OAI21X1_16 ( .A(_108_), .B(_109_), .C(w_C_7_), .Y(_110_) );
NAND2X1 NAND2X1_21 ( .A(_110_), .B(_114_), .Y(_86__7_) );
INVX1 INVX1_41 ( .A(w_C_8_), .Y(_118_) );
OR2X2 OR2X2_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_119_) );
NAND2X1 NAND2X1_22 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_120_) );
NAND3X1 NAND3X1_20 ( .A(_118_), .B(_120_), .C(_119_), .Y(_121_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_115_) );
AND2X2 AND2X2_12 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_116_) );
OAI21X1 OAI21X1_17 ( .A(_115_), .B(_116_), .C(w_C_8_), .Y(_117_) );
NAND2X1 NAND2X1_23 ( .A(_117_), .B(_121_), .Y(_86__8_) );
INVX1 INVX1_42 ( .A(w_C_9_), .Y(_125_) );
OR2X2 OR2X2_10 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_126_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_127_) );
NAND3X1 NAND3X1_21 ( .A(_125_), .B(_127_), .C(_126_), .Y(_128_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_122_) );
AND2X2 AND2X2_13 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_123_) );
OAI21X1 OAI21X1_18 ( .A(_122_), .B(_123_), .C(w_C_9_), .Y(_124_) );
NAND2X1 NAND2X1_25 ( .A(_124_), .B(_128_), .Y(_86__9_) );
INVX1 INVX1_43 ( .A(w_C_10_), .Y(_132_) );
OR2X2 OR2X2_11 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_133_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_134_) );
NAND3X1 NAND3X1_22 ( .A(_132_), .B(_134_), .C(_133_), .Y(_135_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_129_) );
AND2X2 AND2X2_14 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_130_) );
OAI21X1 OAI21X1_19 ( .A(_129_), .B(_130_), .C(w_C_10_), .Y(_131_) );
NAND2X1 NAND2X1_27 ( .A(_131_), .B(_135_), .Y(_86__10_) );
INVX1 INVX1_44 ( .A(w_C_11_), .Y(_139_) );
OR2X2 OR2X2_12 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_140_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_141_) );
NAND3X1 NAND3X1_23 ( .A(_139_), .B(_141_), .C(_140_), .Y(_142_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_136_) );
AND2X2 AND2X2_15 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_137_) );
OAI21X1 OAI21X1_20 ( .A(_136_), .B(_137_), .C(w_C_11_), .Y(_138_) );
NAND2X1 NAND2X1_29 ( .A(_138_), .B(_142_), .Y(_86__11_) );
INVX1 INVX1_45 ( .A(w_C_12_), .Y(_146_) );
OR2X2 OR2X2_13 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_147_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_148_) );
NAND3X1 NAND3X1_24 ( .A(_146_), .B(_148_), .C(_147_), .Y(_149_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_143_) );
AND2X2 AND2X2_16 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_144_) );
OAI21X1 OAI21X1_21 ( .A(_143_), .B(_144_), .C(w_C_12_), .Y(_145_) );
NAND2X1 NAND2X1_31 ( .A(_145_), .B(_149_), .Y(_86__12_) );
INVX1 INVX1_46 ( .A(w_C_13_), .Y(_153_) );
OR2X2 OR2X2_14 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_154_) );
NAND2X1 NAND2X1_32 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_155_) );
NAND3X1 NAND3X1_25 ( .A(_153_), .B(_155_), .C(_154_), .Y(_156_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_150_) );
AND2X2 AND2X2_17 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_151_) );
OAI21X1 OAI21X1_22 ( .A(_150_), .B(_151_), .C(w_C_13_), .Y(_152_) );
NAND2X1 NAND2X1_33 ( .A(_152_), .B(_156_), .Y(_86__13_) );
INVX1 INVX1_47 ( .A(w_C_14_), .Y(_160_) );
OR2X2 OR2X2_15 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_161_) );
NAND2X1 NAND2X1_34 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_162_) );
NAND3X1 NAND3X1_26 ( .A(_160_), .B(_162_), .C(_161_), .Y(_163_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_157_) );
AND2X2 AND2X2_18 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_158_) );
OAI21X1 OAI21X1_23 ( .A(_157_), .B(_158_), .C(w_C_14_), .Y(_159_) );
NAND2X1 NAND2X1_35 ( .A(_159_), .B(_163_), .Y(_86__14_) );
INVX1 INVX1_48 ( .A(w_C_15_), .Y(_167_) );
OR2X2 OR2X2_16 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_168_) );
NAND2X1 NAND2X1_36 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_169_) );
NAND3X1 NAND3X1_27 ( .A(_167_), .B(_169_), .C(_168_), .Y(_170_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_164_) );
AND2X2 AND2X2_19 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_165_) );
OAI21X1 OAI21X1_24 ( .A(_164_), .B(_165_), .C(w_C_15_), .Y(_166_) );
NAND2X1 NAND2X1_37 ( .A(_166_), .B(_170_), .Y(_86__15_) );
INVX1 INVX1_49 ( .A(w_C_16_), .Y(_174_) );
OR2X2 OR2X2_17 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_175_) );
NAND2X1 NAND2X1_38 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_176_) );
NAND3X1 NAND3X1_28 ( .A(_174_), .B(_176_), .C(_175_), .Y(_177_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_171_) );
AND2X2 AND2X2_20 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_172_) );
OAI21X1 OAI21X1_25 ( .A(_171_), .B(_172_), .C(w_C_16_), .Y(_173_) );
NAND2X1 NAND2X1_39 ( .A(_173_), .B(_177_), .Y(_86__16_) );
INVX1 INVX1_50 ( .A(w_C_17_), .Y(_181_) );
OR2X2 OR2X2_18 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_182_) );
NAND2X1 NAND2X1_40 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_183_) );
NAND3X1 NAND3X1_29 ( .A(_181_), .B(_183_), .C(_182_), .Y(_184_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_178_) );
AND2X2 AND2X2_21 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_179_) );
OAI21X1 OAI21X1_26 ( .A(_178_), .B(_179_), .C(w_C_17_), .Y(_180_) );
NAND2X1 NAND2X1_41 ( .A(_180_), .B(_184_), .Y(_86__17_) );
INVX1 INVX1_51 ( .A(gnd), .Y(_188_) );
OR2X2 OR2X2_19 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_189_) );
NAND2X1 NAND2X1_42 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_190_) );
NAND3X1 NAND3X1_30 ( .A(_188_), .B(_190_), .C(_189_), .Y(_191_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_185_) );
AND2X2 AND2X2_22 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_186_) );
OAI21X1 OAI21X1_27 ( .A(_185_), .B(_186_), .C(gnd), .Y(_187_) );
NAND2X1 NAND2X1_43 ( .A(_187_), .B(_191_), .Y(_86__0_) );
INVX1 INVX1_52 ( .A(w_C_1_), .Y(_195_) );
OR2X2 OR2X2_20 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_196_) );
NAND2X1 NAND2X1_44 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_197_) );
NAND3X1 NAND3X1_31 ( .A(_195_), .B(_197_), .C(_196_), .Y(_198_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_192_) );
AND2X2 AND2X2_23 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_193_) );
OAI21X1 OAI21X1_28 ( .A(_192_), .B(_193_), .C(w_C_1_), .Y(_194_) );
NAND2X1 NAND2X1_45 ( .A(_194_), .B(_198_), .Y(_86__1_) );
INVX1 INVX1_53 ( .A(w_C_2_), .Y(_202_) );
OR2X2 OR2X2_21 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_203_) );
NAND2X1 NAND2X1_46 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_204_) );
NAND3X1 NAND3X1_32 ( .A(_202_), .B(_204_), .C(_203_), .Y(_205_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_199_) );
AND2X2 AND2X2_24 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_200_) );
OAI21X1 OAI21X1_29 ( .A(_199_), .B(_200_), .C(w_C_2_), .Y(_201_) );
NAND2X1 NAND2X1_47 ( .A(_201_), .B(_205_), .Y(_86__2_) );
INVX1 INVX1_54 ( .A(w_C_3_), .Y(_209_) );
OR2X2 OR2X2_22 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_210_) );
NAND2X1 NAND2X1_48 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_211_) );
NAND3X1 NAND3X1_33 ( .A(_209_), .B(_211_), .C(_210_), .Y(_212_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_206_) );
AND2X2 AND2X2_25 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_207_) );
OAI21X1 OAI21X1_30 ( .A(_206_), .B(_207_), .C(w_C_3_), .Y(_208_) );
NAND2X1 NAND2X1_49 ( .A(_208_), .B(_212_), .Y(_86__3_) );
BUFX2 BUFX2_20 ( .A(w_C_18_), .Y(_86__18_) );
BUFX2 BUFX2_21 ( .A(gnd), .Y(w_C_0_) );
endmodule
