module csa_47bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term1[45], i_add_term1[46], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], i_add_term2[45], i_add_term2[46], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], sum[45], sum[46], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term1[45];
input i_add_term1[46];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
input i_add_term2[45];
input i_add_term2[46];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output sum[45];
output sum[46];
output cout;

INVX1 INVX1_1 ( .A(_57__0_), .Y(_159_) );
NAND2X1 NAND2X1_1 ( .A(_58__0_), .B(w_cout_9_), .Y(_160_) );
OAI21X1 OAI21X1_1 ( .A(w_cout_9_), .B(_159_), .C(_160_), .Y(_0__39_) );
INVX1 INVX1_2 ( .A(_57__1_), .Y(_161_) );
NAND2X1 NAND2X1_2 ( .A(w_cout_9_), .B(_58__1_), .Y(_162_) );
OAI21X1 OAI21X1_2 ( .A(w_cout_9_), .B(_161_), .C(_162_), .Y(_0__40_) );
INVX1 INVX1_3 ( .A(_57__2_), .Y(_163_) );
NAND2X1 NAND2X1_3 ( .A(w_cout_9_), .B(_58__2_), .Y(_164_) );
OAI21X1 OAI21X1_3 ( .A(w_cout_9_), .B(_163_), .C(_164_), .Y(_0__41_) );
INVX1 INVX1_4 ( .A(_57__3_), .Y(_165_) );
NAND2X1 NAND2X1_4 ( .A(w_cout_9_), .B(_58__3_), .Y(_166_) );
OAI21X1 OAI21X1_4 ( .A(w_cout_9_), .B(_165_), .C(_166_), .Y(_0__42_) );
INVX1 INVX1_5 ( .A(_61_), .Y(_167_) );
NAND2X1 NAND2X1_5 ( .A(_62_), .B(w_cout_10_), .Y(_168_) );
OAI21X1 OAI21X1_5 ( .A(w_cout_10_), .B(_167_), .C(_168_), .Y(w_cout_11_) );
INVX1 INVX1_6 ( .A(_63__0_), .Y(_169_) );
NAND2X1 NAND2X1_6 ( .A(_64__0_), .B(w_cout_10_), .Y(_170_) );
OAI21X1 OAI21X1_6 ( .A(w_cout_10_), .B(_169_), .C(_170_), .Y(_0__43_) );
INVX1 INVX1_7 ( .A(_63__1_), .Y(_171_) );
NAND2X1 NAND2X1_7 ( .A(w_cout_10_), .B(_64__1_), .Y(_172_) );
OAI21X1 OAI21X1_7 ( .A(w_cout_10_), .B(_171_), .C(_172_), .Y(_0__44_) );
INVX1 INVX1_8 ( .A(_63__2_), .Y(_173_) );
NAND2X1 NAND2X1_8 ( .A(w_cout_10_), .B(_64__2_), .Y(_174_) );
OAI21X1 OAI21X1_8 ( .A(w_cout_10_), .B(_173_), .C(_174_), .Y(_0__45_) );
INVX1 INVX1_9 ( .A(_63__3_), .Y(_175_) );
NAND2X1 NAND2X1_9 ( .A(w_cout_10_), .B(_64__3_), .Y(_176_) );
OAI21X1 OAI21X1_9 ( .A(w_cout_10_), .B(_175_), .C(_176_), .Y(_0__46_) );
INVX1 INVX1_10 ( .A(1'b0), .Y(_180_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_181_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_182_) );
NAND3X1 NAND3X1_1 ( .A(_180_), .B(_182_), .C(_181_), .Y(_183_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_177_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_178_) );
OAI21X1 OAI21X1_10 ( .A(_177_), .B(_178_), .C(1'b0), .Y(_179_) );
NAND2X1 NAND2X1_11 ( .A(_179_), .B(_183_), .Y(_3__0_) );
OAI21X1 OAI21X1_11 ( .A(_180_), .B(_177_), .C(_182_), .Y(_5__1_) );
INVX1 INVX1_11 ( .A(_5__1_), .Y(_187_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_188_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_189_) );
NAND3X1 NAND3X1_2 ( .A(_187_), .B(_189_), .C(_188_), .Y(_190_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_184_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_185_) );
OAI21X1 OAI21X1_12 ( .A(_184_), .B(_185_), .C(_5__1_), .Y(_186_) );
NAND2X1 NAND2X1_13 ( .A(_186_), .B(_190_), .Y(_3__1_) );
OAI21X1 OAI21X1_13 ( .A(_187_), .B(_184_), .C(_189_), .Y(_5__2_) );
INVX1 INVX1_12 ( .A(_5__2_), .Y(_194_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_195_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_196_) );
NAND3X1 NAND3X1_3 ( .A(_194_), .B(_196_), .C(_195_), .Y(_197_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_191_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_192_) );
OAI21X1 OAI21X1_14 ( .A(_191_), .B(_192_), .C(_5__2_), .Y(_193_) );
NAND2X1 NAND2X1_15 ( .A(_193_), .B(_197_), .Y(_3__2_) );
OAI21X1 OAI21X1_15 ( .A(_194_), .B(_191_), .C(_196_), .Y(_5__3_) );
INVX1 INVX1_13 ( .A(_5__3_), .Y(_201_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_202_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_203_) );
NAND3X1 NAND3X1_4 ( .A(_201_), .B(_203_), .C(_202_), .Y(_204_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_198_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_199_) );
OAI21X1 OAI21X1_16 ( .A(_198_), .B(_199_), .C(_5__3_), .Y(_200_) );
NAND2X1 NAND2X1_17 ( .A(_200_), .B(_204_), .Y(_3__3_) );
OAI21X1 OAI21X1_17 ( .A(_201_), .B(_198_), .C(_203_), .Y(_1_) );
INVX1 INVX1_14 ( .A(1'b1), .Y(_208_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_209_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_210_) );
NAND3X1 NAND3X1_5 ( .A(_208_), .B(_210_), .C(_209_), .Y(_211_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_205_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_206_) );
OAI21X1 OAI21X1_18 ( .A(_205_), .B(_206_), .C(1'b1), .Y(_207_) );
NAND2X1 NAND2X1_19 ( .A(_207_), .B(_211_), .Y(_4__0_) );
OAI21X1 OAI21X1_19 ( .A(_208_), .B(_205_), .C(_210_), .Y(_6__1_) );
INVX1 INVX1_15 ( .A(_6__1_), .Y(_215_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_216_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_217_) );
NAND3X1 NAND3X1_6 ( .A(_215_), .B(_217_), .C(_216_), .Y(_218_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_212_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_213_) );
OAI21X1 OAI21X1_20 ( .A(_212_), .B(_213_), .C(_6__1_), .Y(_214_) );
NAND2X1 NAND2X1_21 ( .A(_214_), .B(_218_), .Y(_4__1_) );
OAI21X1 OAI21X1_21 ( .A(_215_), .B(_212_), .C(_217_), .Y(_6__2_) );
INVX1 INVX1_16 ( .A(_6__2_), .Y(_222_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_223_) );
NAND2X1 NAND2X1_22 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_224_) );
NAND3X1 NAND3X1_7 ( .A(_222_), .B(_224_), .C(_223_), .Y(_225_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_219_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_220_) );
OAI21X1 OAI21X1_22 ( .A(_219_), .B(_220_), .C(_6__2_), .Y(_221_) );
NAND2X1 NAND2X1_23 ( .A(_221_), .B(_225_), .Y(_4__2_) );
OAI21X1 OAI21X1_23 ( .A(_222_), .B(_219_), .C(_224_), .Y(_6__3_) );
INVX1 INVX1_17 ( .A(_6__3_), .Y(_229_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_230_) );
NAND2X1 NAND2X1_24 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_231_) );
NAND3X1 NAND3X1_8 ( .A(_229_), .B(_231_), .C(_230_), .Y(_232_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_226_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_227_) );
OAI21X1 OAI21X1_24 ( .A(_226_), .B(_227_), .C(_6__3_), .Y(_228_) );
NAND2X1 NAND2X1_25 ( .A(_228_), .B(_232_), .Y(_4__3_) );
OAI21X1 OAI21X1_25 ( .A(_229_), .B(_226_), .C(_231_), .Y(_2_) );
INVX1 INVX1_18 ( .A(1'b0), .Y(_236_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_237_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_238_) );
NAND3X1 NAND3X1_9 ( .A(_236_), .B(_238_), .C(_237_), .Y(_239_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_233_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_234_) );
OAI21X1 OAI21X1_26 ( .A(_233_), .B(_234_), .C(1'b0), .Y(_235_) );
NAND2X1 NAND2X1_27 ( .A(_235_), .B(_239_), .Y(_9__0_) );
OAI21X1 OAI21X1_27 ( .A(_236_), .B(_233_), .C(_238_), .Y(_11__1_) );
INVX1 INVX1_19 ( .A(_11__1_), .Y(_243_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_244_) );
NAND2X1 NAND2X1_28 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_245_) );
NAND3X1 NAND3X1_10 ( .A(_243_), .B(_245_), .C(_244_), .Y(_246_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_240_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_241_) );
OAI21X1 OAI21X1_28 ( .A(_240_), .B(_241_), .C(_11__1_), .Y(_242_) );
NAND2X1 NAND2X1_29 ( .A(_242_), .B(_246_), .Y(_9__1_) );
OAI21X1 OAI21X1_29 ( .A(_243_), .B(_240_), .C(_245_), .Y(_11__2_) );
INVX1 INVX1_20 ( .A(_11__2_), .Y(_250_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_251_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_252_) );
NAND3X1 NAND3X1_11 ( .A(_250_), .B(_252_), .C(_251_), .Y(_253_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_247_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_248_) );
OAI21X1 OAI21X1_30 ( .A(_247_), .B(_248_), .C(_11__2_), .Y(_249_) );
NAND2X1 NAND2X1_31 ( .A(_249_), .B(_253_), .Y(_9__2_) );
OAI21X1 OAI21X1_31 ( .A(_250_), .B(_247_), .C(_252_), .Y(_11__3_) );
INVX1 INVX1_21 ( .A(_11__3_), .Y(_257_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_258_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_259_) );
NAND3X1 NAND3X1_12 ( .A(_257_), .B(_259_), .C(_258_), .Y(_260_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_254_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_255_) );
OAI21X1 OAI21X1_32 ( .A(_254_), .B(_255_), .C(_11__3_), .Y(_256_) );
NAND2X1 NAND2X1_33 ( .A(_256_), .B(_260_), .Y(_9__3_) );
OAI21X1 OAI21X1_33 ( .A(_257_), .B(_254_), .C(_259_), .Y(_7_) );
INVX1 INVX1_22 ( .A(1'b1), .Y(_264_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_265_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_266_) );
NAND3X1 NAND3X1_13 ( .A(_264_), .B(_266_), .C(_265_), .Y(_267_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_261_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_262_) );
OAI21X1 OAI21X1_34 ( .A(_261_), .B(_262_), .C(1'b1), .Y(_263_) );
NAND2X1 NAND2X1_35 ( .A(_263_), .B(_267_), .Y(_10__0_) );
OAI21X1 OAI21X1_35 ( .A(_264_), .B(_261_), .C(_266_), .Y(_12__1_) );
INVX1 INVX1_23 ( .A(_12__1_), .Y(_271_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_272_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_273_) );
NAND3X1 NAND3X1_14 ( .A(_271_), .B(_273_), .C(_272_), .Y(_274_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_268_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_269_) );
OAI21X1 OAI21X1_36 ( .A(_268_), .B(_269_), .C(_12__1_), .Y(_270_) );
NAND2X1 NAND2X1_37 ( .A(_270_), .B(_274_), .Y(_10__1_) );
OAI21X1 OAI21X1_37 ( .A(_271_), .B(_268_), .C(_273_), .Y(_12__2_) );
INVX1 INVX1_24 ( .A(_12__2_), .Y(_278_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_279_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_280_) );
NAND3X1 NAND3X1_15 ( .A(_278_), .B(_280_), .C(_279_), .Y(_281_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_275_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_276_) );
OAI21X1 OAI21X1_38 ( .A(_275_), .B(_276_), .C(_12__2_), .Y(_277_) );
NAND2X1 NAND2X1_39 ( .A(_277_), .B(_281_), .Y(_10__2_) );
OAI21X1 OAI21X1_39 ( .A(_278_), .B(_275_), .C(_280_), .Y(_12__3_) );
INVX1 INVX1_25 ( .A(_12__3_), .Y(_285_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_286_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_287_) );
NAND3X1 NAND3X1_16 ( .A(_285_), .B(_287_), .C(_286_), .Y(_288_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_282_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_283_) );
OAI21X1 OAI21X1_40 ( .A(_282_), .B(_283_), .C(_12__3_), .Y(_284_) );
NAND2X1 NAND2X1_41 ( .A(_284_), .B(_288_), .Y(_10__3_) );
OAI21X1 OAI21X1_41 ( .A(_285_), .B(_282_), .C(_287_), .Y(_8_) );
INVX1 INVX1_26 ( .A(1'b0), .Y(_292_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_293_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_294_) );
NAND3X1 NAND3X1_17 ( .A(_292_), .B(_294_), .C(_293_), .Y(_295_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_289_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_290_) );
OAI21X1 OAI21X1_42 ( .A(_289_), .B(_290_), .C(1'b0), .Y(_291_) );
NAND2X1 NAND2X1_43 ( .A(_291_), .B(_295_), .Y(_15__0_) );
OAI21X1 OAI21X1_43 ( .A(_292_), .B(_289_), .C(_294_), .Y(_17__1_) );
INVX1 INVX1_27 ( .A(_17__1_), .Y(_299_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_300_) );
NAND2X1 NAND2X1_44 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_301_) );
NAND3X1 NAND3X1_18 ( .A(_299_), .B(_301_), .C(_300_), .Y(_302_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_296_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_297_) );
OAI21X1 OAI21X1_44 ( .A(_296_), .B(_297_), .C(_17__1_), .Y(_298_) );
NAND2X1 NAND2X1_45 ( .A(_298_), .B(_302_), .Y(_15__1_) );
OAI21X1 OAI21X1_45 ( .A(_299_), .B(_296_), .C(_301_), .Y(_17__2_) );
INVX1 INVX1_28 ( .A(_17__2_), .Y(_306_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_307_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_308_) );
NAND3X1 NAND3X1_19 ( .A(_306_), .B(_308_), .C(_307_), .Y(_309_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_303_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_304_) );
OAI21X1 OAI21X1_46 ( .A(_303_), .B(_304_), .C(_17__2_), .Y(_305_) );
NAND2X1 NAND2X1_47 ( .A(_305_), .B(_309_), .Y(_15__2_) );
OAI21X1 OAI21X1_47 ( .A(_306_), .B(_303_), .C(_308_), .Y(_17__3_) );
INVX1 INVX1_29 ( .A(_17__3_), .Y(_313_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_314_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_315_) );
NAND3X1 NAND3X1_20 ( .A(_313_), .B(_315_), .C(_314_), .Y(_316_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_310_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_311_) );
OAI21X1 OAI21X1_48 ( .A(_310_), .B(_311_), .C(_17__3_), .Y(_312_) );
NAND2X1 NAND2X1_49 ( .A(_312_), .B(_316_), .Y(_15__3_) );
OAI21X1 OAI21X1_49 ( .A(_313_), .B(_310_), .C(_315_), .Y(_13_) );
INVX1 INVX1_30 ( .A(1'b1), .Y(_320_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_321_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_322_) );
NAND3X1 NAND3X1_21 ( .A(_320_), .B(_322_), .C(_321_), .Y(_323_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_317_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_318_) );
OAI21X1 OAI21X1_50 ( .A(_317_), .B(_318_), .C(1'b1), .Y(_319_) );
NAND2X1 NAND2X1_51 ( .A(_319_), .B(_323_), .Y(_16__0_) );
OAI21X1 OAI21X1_51 ( .A(_320_), .B(_317_), .C(_322_), .Y(_18__1_) );
INVX1 INVX1_31 ( .A(_18__1_), .Y(_327_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_328_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_329_) );
NAND3X1 NAND3X1_22 ( .A(_327_), .B(_329_), .C(_328_), .Y(_330_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_324_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_325_) );
OAI21X1 OAI21X1_52 ( .A(_324_), .B(_325_), .C(_18__1_), .Y(_326_) );
NAND2X1 NAND2X1_53 ( .A(_326_), .B(_330_), .Y(_16__1_) );
OAI21X1 OAI21X1_53 ( .A(_327_), .B(_324_), .C(_329_), .Y(_18__2_) );
INVX1 INVX1_32 ( .A(_18__2_), .Y(_334_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_335_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_336_) );
NAND3X1 NAND3X1_23 ( .A(_334_), .B(_336_), .C(_335_), .Y(_337_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_331_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_332_) );
OAI21X1 OAI21X1_54 ( .A(_331_), .B(_332_), .C(_18__2_), .Y(_333_) );
NAND2X1 NAND2X1_55 ( .A(_333_), .B(_337_), .Y(_16__2_) );
OAI21X1 OAI21X1_55 ( .A(_334_), .B(_331_), .C(_336_), .Y(_18__3_) );
INVX1 INVX1_33 ( .A(_18__3_), .Y(_341_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_342_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_343_) );
NAND3X1 NAND3X1_24 ( .A(_341_), .B(_343_), .C(_342_), .Y(_344_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_338_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_339_) );
OAI21X1 OAI21X1_56 ( .A(_338_), .B(_339_), .C(_18__3_), .Y(_340_) );
NAND2X1 NAND2X1_57 ( .A(_340_), .B(_344_), .Y(_16__3_) );
OAI21X1 OAI21X1_57 ( .A(_341_), .B(_338_), .C(_343_), .Y(_14_) );
INVX1 INVX1_34 ( .A(1'b0), .Y(_348_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_349_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_350_) );
NAND3X1 NAND3X1_25 ( .A(_348_), .B(_350_), .C(_349_), .Y(_351_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_345_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_346_) );
OAI21X1 OAI21X1_58 ( .A(_345_), .B(_346_), .C(1'b0), .Y(_347_) );
NAND2X1 NAND2X1_59 ( .A(_347_), .B(_351_), .Y(_21__0_) );
OAI21X1 OAI21X1_59 ( .A(_348_), .B(_345_), .C(_350_), .Y(_23__1_) );
INVX1 INVX1_35 ( .A(_23__1_), .Y(_355_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_356_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_357_) );
NAND3X1 NAND3X1_26 ( .A(_355_), .B(_357_), .C(_356_), .Y(_358_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_352_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_353_) );
OAI21X1 OAI21X1_60 ( .A(_352_), .B(_353_), .C(_23__1_), .Y(_354_) );
NAND2X1 NAND2X1_61 ( .A(_354_), .B(_358_), .Y(_21__1_) );
OAI21X1 OAI21X1_61 ( .A(_355_), .B(_352_), .C(_357_), .Y(_23__2_) );
INVX1 INVX1_36 ( .A(_23__2_), .Y(_362_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_363_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_364_) );
NAND3X1 NAND3X1_27 ( .A(_362_), .B(_364_), .C(_363_), .Y(_365_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_359_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_360_) );
OAI21X1 OAI21X1_62 ( .A(_359_), .B(_360_), .C(_23__2_), .Y(_361_) );
NAND2X1 NAND2X1_63 ( .A(_361_), .B(_365_), .Y(_21__2_) );
OAI21X1 OAI21X1_63 ( .A(_362_), .B(_359_), .C(_364_), .Y(_23__3_) );
INVX1 INVX1_37 ( .A(_23__3_), .Y(_369_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_370_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_371_) );
NAND3X1 NAND3X1_28 ( .A(_369_), .B(_371_), .C(_370_), .Y(_372_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_366_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_367_) );
OAI21X1 OAI21X1_64 ( .A(_366_), .B(_367_), .C(_23__3_), .Y(_368_) );
NAND2X1 NAND2X1_65 ( .A(_368_), .B(_372_), .Y(_21__3_) );
OAI21X1 OAI21X1_65 ( .A(_369_), .B(_366_), .C(_371_), .Y(_19_) );
INVX1 INVX1_38 ( .A(1'b1), .Y(_376_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_377_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_378_) );
NAND3X1 NAND3X1_29 ( .A(_376_), .B(_378_), .C(_377_), .Y(_379_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_373_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_374_) );
OAI21X1 OAI21X1_66 ( .A(_373_), .B(_374_), .C(1'b1), .Y(_375_) );
NAND2X1 NAND2X1_67 ( .A(_375_), .B(_379_), .Y(_22__0_) );
OAI21X1 OAI21X1_67 ( .A(_376_), .B(_373_), .C(_378_), .Y(_24__1_) );
INVX1 INVX1_39 ( .A(_24__1_), .Y(_383_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_384_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_385_) );
NAND3X1 NAND3X1_30 ( .A(_383_), .B(_385_), .C(_384_), .Y(_386_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_380_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_381_) );
OAI21X1 OAI21X1_68 ( .A(_380_), .B(_381_), .C(_24__1_), .Y(_382_) );
NAND2X1 NAND2X1_69 ( .A(_382_), .B(_386_), .Y(_22__1_) );
OAI21X1 OAI21X1_69 ( .A(_383_), .B(_380_), .C(_385_), .Y(_24__2_) );
INVX1 INVX1_40 ( .A(_24__2_), .Y(_390_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_391_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_392_) );
NAND3X1 NAND3X1_31 ( .A(_390_), .B(_392_), .C(_391_), .Y(_393_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_387_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_388_) );
OAI21X1 OAI21X1_70 ( .A(_387_), .B(_388_), .C(_24__2_), .Y(_389_) );
NAND2X1 NAND2X1_71 ( .A(_389_), .B(_393_), .Y(_22__2_) );
OAI21X1 OAI21X1_71 ( .A(_390_), .B(_387_), .C(_392_), .Y(_24__3_) );
INVX1 INVX1_41 ( .A(_24__3_), .Y(_397_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_398_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_399_) );
NAND3X1 NAND3X1_32 ( .A(_397_), .B(_399_), .C(_398_), .Y(_400_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_394_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_395_) );
OAI21X1 OAI21X1_72 ( .A(_394_), .B(_395_), .C(_24__3_), .Y(_396_) );
NAND2X1 NAND2X1_73 ( .A(_396_), .B(_400_), .Y(_22__3_) );
OAI21X1 OAI21X1_73 ( .A(_397_), .B(_394_), .C(_399_), .Y(_20_) );
INVX1 INVX1_42 ( .A(1'b0), .Y(_404_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_405_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_406_) );
NAND3X1 NAND3X1_33 ( .A(_404_), .B(_406_), .C(_405_), .Y(_407_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_401_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_402_) );
OAI21X1 OAI21X1_74 ( .A(_401_), .B(_402_), .C(1'b0), .Y(_403_) );
NAND2X1 NAND2X1_75 ( .A(_403_), .B(_407_), .Y(_27__0_) );
OAI21X1 OAI21X1_75 ( .A(_404_), .B(_401_), .C(_406_), .Y(_29__1_) );
INVX1 INVX1_43 ( .A(_29__1_), .Y(_411_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_412_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_413_) );
NAND3X1 NAND3X1_34 ( .A(_411_), .B(_413_), .C(_412_), .Y(_414_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_408_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_409_) );
OAI21X1 OAI21X1_76 ( .A(_408_), .B(_409_), .C(_29__1_), .Y(_410_) );
NAND2X1 NAND2X1_77 ( .A(_410_), .B(_414_), .Y(_27__1_) );
OAI21X1 OAI21X1_77 ( .A(_411_), .B(_408_), .C(_413_), .Y(_29__2_) );
INVX1 INVX1_44 ( .A(_29__2_), .Y(_418_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_419_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_420_) );
NAND3X1 NAND3X1_35 ( .A(_418_), .B(_420_), .C(_419_), .Y(_421_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_415_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_416_) );
OAI21X1 OAI21X1_78 ( .A(_415_), .B(_416_), .C(_29__2_), .Y(_417_) );
NAND2X1 NAND2X1_79 ( .A(_417_), .B(_421_), .Y(_27__2_) );
OAI21X1 OAI21X1_79 ( .A(_418_), .B(_415_), .C(_420_), .Y(_29__3_) );
INVX1 INVX1_45 ( .A(_29__3_), .Y(_425_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_426_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_427_) );
NAND3X1 NAND3X1_36 ( .A(_425_), .B(_427_), .C(_426_), .Y(_428_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_422_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_423_) );
OAI21X1 OAI21X1_80 ( .A(_422_), .B(_423_), .C(_29__3_), .Y(_424_) );
NAND2X1 NAND2X1_81 ( .A(_424_), .B(_428_), .Y(_27__3_) );
OAI21X1 OAI21X1_81 ( .A(_425_), .B(_422_), .C(_427_), .Y(_25_) );
INVX1 INVX1_46 ( .A(1'b1), .Y(_432_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_433_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_434_) );
NAND3X1 NAND3X1_37 ( .A(_432_), .B(_434_), .C(_433_), .Y(_435_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_429_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_430_) );
OAI21X1 OAI21X1_82 ( .A(_429_), .B(_430_), .C(1'b1), .Y(_431_) );
NAND2X1 NAND2X1_83 ( .A(_431_), .B(_435_), .Y(_28__0_) );
OAI21X1 OAI21X1_83 ( .A(_432_), .B(_429_), .C(_434_), .Y(_30__1_) );
INVX1 INVX1_47 ( .A(_30__1_), .Y(_439_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_440_) );
NAND2X1 NAND2X1_84 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_441_) );
NAND3X1 NAND3X1_38 ( .A(_439_), .B(_441_), .C(_440_), .Y(_442_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_436_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_437_) );
OAI21X1 OAI21X1_84 ( .A(_436_), .B(_437_), .C(_30__1_), .Y(_438_) );
NAND2X1 NAND2X1_85 ( .A(_438_), .B(_442_), .Y(_28__1_) );
OAI21X1 OAI21X1_85 ( .A(_439_), .B(_436_), .C(_441_), .Y(_30__2_) );
INVX1 INVX1_48 ( .A(_30__2_), .Y(_446_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_447_) );
NAND2X1 NAND2X1_86 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_448_) );
NAND3X1 NAND3X1_39 ( .A(_446_), .B(_448_), .C(_447_), .Y(_449_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_443_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_444_) );
OAI21X1 OAI21X1_86 ( .A(_443_), .B(_444_), .C(_30__2_), .Y(_445_) );
NAND2X1 NAND2X1_87 ( .A(_445_), .B(_449_), .Y(_28__2_) );
OAI21X1 OAI21X1_87 ( .A(_446_), .B(_443_), .C(_448_), .Y(_30__3_) );
INVX1 INVX1_49 ( .A(_30__3_), .Y(_453_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_454_) );
NAND2X1 NAND2X1_88 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_455_) );
NAND3X1 NAND3X1_40 ( .A(_453_), .B(_455_), .C(_454_), .Y(_456_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_450_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_451_) );
OAI21X1 OAI21X1_88 ( .A(_450_), .B(_451_), .C(_30__3_), .Y(_452_) );
NAND2X1 NAND2X1_89 ( .A(_452_), .B(_456_), .Y(_28__3_) );
OAI21X1 OAI21X1_89 ( .A(_453_), .B(_450_), .C(_455_), .Y(_26_) );
INVX1 INVX1_50 ( .A(1'b0), .Y(_460_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_461_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_462_) );
NAND3X1 NAND3X1_41 ( .A(_460_), .B(_462_), .C(_461_), .Y(_463_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_457_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_458_) );
OAI21X1 OAI21X1_90 ( .A(_457_), .B(_458_), .C(1'b0), .Y(_459_) );
NAND2X1 NAND2X1_91 ( .A(_459_), .B(_463_), .Y(_33__0_) );
OAI21X1 OAI21X1_91 ( .A(_460_), .B(_457_), .C(_462_), .Y(_35__1_) );
INVX1 INVX1_51 ( .A(_35__1_), .Y(_467_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_468_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_469_) );
NAND3X1 NAND3X1_42 ( .A(_467_), .B(_469_), .C(_468_), .Y(_470_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_464_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_465_) );
OAI21X1 OAI21X1_92 ( .A(_464_), .B(_465_), .C(_35__1_), .Y(_466_) );
NAND2X1 NAND2X1_93 ( .A(_466_), .B(_470_), .Y(_33__1_) );
OAI21X1 OAI21X1_93 ( .A(_467_), .B(_464_), .C(_469_), .Y(_35__2_) );
INVX1 INVX1_52 ( .A(_35__2_), .Y(_474_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_475_) );
NAND2X1 NAND2X1_94 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_476_) );
NAND3X1 NAND3X1_43 ( .A(_474_), .B(_476_), .C(_475_), .Y(_477_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_471_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_472_) );
OAI21X1 OAI21X1_94 ( .A(_471_), .B(_472_), .C(_35__2_), .Y(_473_) );
NAND2X1 NAND2X1_95 ( .A(_473_), .B(_477_), .Y(_33__2_) );
OAI21X1 OAI21X1_95 ( .A(_474_), .B(_471_), .C(_476_), .Y(_35__3_) );
INVX1 INVX1_53 ( .A(_35__3_), .Y(_481_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_482_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_483_) );
NAND3X1 NAND3X1_44 ( .A(_481_), .B(_483_), .C(_482_), .Y(_484_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_478_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_479_) );
OAI21X1 OAI21X1_96 ( .A(_478_), .B(_479_), .C(_35__3_), .Y(_480_) );
NAND2X1 NAND2X1_97 ( .A(_480_), .B(_484_), .Y(_33__3_) );
OAI21X1 OAI21X1_97 ( .A(_481_), .B(_478_), .C(_483_), .Y(_31_) );
INVX1 INVX1_54 ( .A(1'b1), .Y(_488_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_489_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_490_) );
NAND3X1 NAND3X1_45 ( .A(_488_), .B(_490_), .C(_489_), .Y(_491_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_485_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_486_) );
OAI21X1 OAI21X1_98 ( .A(_485_), .B(_486_), .C(1'b1), .Y(_487_) );
NAND2X1 NAND2X1_99 ( .A(_487_), .B(_491_), .Y(_34__0_) );
OAI21X1 OAI21X1_99 ( .A(_488_), .B(_485_), .C(_490_), .Y(_36__1_) );
INVX1 INVX1_55 ( .A(_36__1_), .Y(_495_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_496_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_497_) );
NAND3X1 NAND3X1_46 ( .A(_495_), .B(_497_), .C(_496_), .Y(_498_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_492_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_493_) );
OAI21X1 OAI21X1_100 ( .A(_492_), .B(_493_), .C(_36__1_), .Y(_494_) );
NAND2X1 NAND2X1_101 ( .A(_494_), .B(_498_), .Y(_34__1_) );
OAI21X1 OAI21X1_101 ( .A(_495_), .B(_492_), .C(_497_), .Y(_36__2_) );
INVX1 INVX1_56 ( .A(_36__2_), .Y(_502_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_503_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_504_) );
NAND3X1 NAND3X1_47 ( .A(_502_), .B(_504_), .C(_503_), .Y(_505_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_499_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_500_) );
OAI21X1 OAI21X1_102 ( .A(_499_), .B(_500_), .C(_36__2_), .Y(_501_) );
NAND2X1 NAND2X1_103 ( .A(_501_), .B(_505_), .Y(_34__2_) );
OAI21X1 OAI21X1_103 ( .A(_502_), .B(_499_), .C(_504_), .Y(_36__3_) );
INVX1 INVX1_57 ( .A(_36__3_), .Y(_509_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_510_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_511_) );
NAND3X1 NAND3X1_48 ( .A(_509_), .B(_511_), .C(_510_), .Y(_512_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_506_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_507_) );
OAI21X1 OAI21X1_104 ( .A(_506_), .B(_507_), .C(_36__3_), .Y(_508_) );
NAND2X1 NAND2X1_105 ( .A(_508_), .B(_512_), .Y(_34__3_) );
OAI21X1 OAI21X1_105 ( .A(_509_), .B(_506_), .C(_511_), .Y(_32_) );
INVX1 INVX1_58 ( .A(1'b0), .Y(_516_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_517_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_518_) );
NAND3X1 NAND3X1_49 ( .A(_516_), .B(_518_), .C(_517_), .Y(_519_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_513_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_514_) );
OAI21X1 OAI21X1_106 ( .A(_513_), .B(_514_), .C(1'b0), .Y(_515_) );
NAND2X1 NAND2X1_107 ( .A(_515_), .B(_519_), .Y(_39__0_) );
OAI21X1 OAI21X1_107 ( .A(_516_), .B(_513_), .C(_518_), .Y(_41__1_) );
INVX1 INVX1_59 ( .A(_41__1_), .Y(_523_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_524_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_525_) );
NAND3X1 NAND3X1_50 ( .A(_523_), .B(_525_), .C(_524_), .Y(_526_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_520_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_521_) );
OAI21X1 OAI21X1_108 ( .A(_520_), .B(_521_), .C(_41__1_), .Y(_522_) );
NAND2X1 NAND2X1_109 ( .A(_522_), .B(_526_), .Y(_39__1_) );
OAI21X1 OAI21X1_109 ( .A(_523_), .B(_520_), .C(_525_), .Y(_41__2_) );
INVX1 INVX1_60 ( .A(_41__2_), .Y(_530_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_531_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_532_) );
NAND3X1 NAND3X1_51 ( .A(_530_), .B(_532_), .C(_531_), .Y(_533_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_527_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_528_) );
OAI21X1 OAI21X1_110 ( .A(_527_), .B(_528_), .C(_41__2_), .Y(_529_) );
NAND2X1 NAND2X1_111 ( .A(_529_), .B(_533_), .Y(_39__2_) );
OAI21X1 OAI21X1_111 ( .A(_530_), .B(_527_), .C(_532_), .Y(_41__3_) );
INVX1 INVX1_61 ( .A(_41__3_), .Y(_537_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_538_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_539_) );
NAND3X1 NAND3X1_52 ( .A(_537_), .B(_539_), .C(_538_), .Y(_540_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_534_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_535_) );
OAI21X1 OAI21X1_112 ( .A(_534_), .B(_535_), .C(_41__3_), .Y(_536_) );
NAND2X1 NAND2X1_113 ( .A(_536_), .B(_540_), .Y(_39__3_) );
OAI21X1 OAI21X1_113 ( .A(_537_), .B(_534_), .C(_539_), .Y(_37_) );
INVX1 INVX1_62 ( .A(1'b1), .Y(_544_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_545_) );
NAND2X1 NAND2X1_114 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_546_) );
NAND3X1 NAND3X1_53 ( .A(_544_), .B(_546_), .C(_545_), .Y(_547_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_541_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_542_) );
OAI21X1 OAI21X1_114 ( .A(_541_), .B(_542_), .C(1'b1), .Y(_543_) );
NAND2X1 NAND2X1_115 ( .A(_543_), .B(_547_), .Y(_40__0_) );
OAI21X1 OAI21X1_115 ( .A(_544_), .B(_541_), .C(_546_), .Y(_42__1_) );
INVX1 INVX1_63 ( .A(_42__1_), .Y(_551_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_552_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_553_) );
NAND3X1 NAND3X1_54 ( .A(_551_), .B(_553_), .C(_552_), .Y(_554_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_548_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_549_) );
OAI21X1 OAI21X1_116 ( .A(_548_), .B(_549_), .C(_42__1_), .Y(_550_) );
NAND2X1 NAND2X1_117 ( .A(_550_), .B(_554_), .Y(_40__1_) );
OAI21X1 OAI21X1_117 ( .A(_551_), .B(_548_), .C(_553_), .Y(_42__2_) );
INVX1 INVX1_64 ( .A(_42__2_), .Y(_558_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_559_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_560_) );
NAND3X1 NAND3X1_55 ( .A(_558_), .B(_560_), .C(_559_), .Y(_561_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_555_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_556_) );
OAI21X1 OAI21X1_118 ( .A(_555_), .B(_556_), .C(_42__2_), .Y(_557_) );
NAND2X1 NAND2X1_119 ( .A(_557_), .B(_561_), .Y(_40__2_) );
OAI21X1 OAI21X1_119 ( .A(_558_), .B(_555_), .C(_560_), .Y(_42__3_) );
INVX1 INVX1_65 ( .A(_42__3_), .Y(_565_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_566_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_567_) );
NAND3X1 NAND3X1_56 ( .A(_565_), .B(_567_), .C(_566_), .Y(_568_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_562_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_563_) );
OAI21X1 OAI21X1_120 ( .A(_562_), .B(_563_), .C(_42__3_), .Y(_564_) );
NAND2X1 NAND2X1_121 ( .A(_564_), .B(_568_), .Y(_40__3_) );
OAI21X1 OAI21X1_121 ( .A(_565_), .B(_562_), .C(_567_), .Y(_38_) );
INVX1 INVX1_66 ( .A(1'b0), .Y(_572_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_573_) );
NAND2X1 NAND2X1_122 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_574_) );
NAND3X1 NAND3X1_57 ( .A(_572_), .B(_574_), .C(_573_), .Y(_575_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_569_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_570_) );
OAI21X1 OAI21X1_122 ( .A(_569_), .B(_570_), .C(1'b0), .Y(_571_) );
NAND2X1 NAND2X1_123 ( .A(_571_), .B(_575_), .Y(_45__0_) );
OAI21X1 OAI21X1_123 ( .A(_572_), .B(_569_), .C(_574_), .Y(_47__1_) );
INVX1 INVX1_67 ( .A(_47__1_), .Y(_579_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_580_) );
NAND2X1 NAND2X1_124 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_581_) );
NAND3X1 NAND3X1_58 ( .A(_579_), .B(_581_), .C(_580_), .Y(_582_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_576_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_577_) );
OAI21X1 OAI21X1_124 ( .A(_576_), .B(_577_), .C(_47__1_), .Y(_578_) );
NAND2X1 NAND2X1_125 ( .A(_578_), .B(_582_), .Y(_45__1_) );
OAI21X1 OAI21X1_125 ( .A(_579_), .B(_576_), .C(_581_), .Y(_47__2_) );
INVX1 INVX1_68 ( .A(_47__2_), .Y(_586_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_587_) );
NAND2X1 NAND2X1_126 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_588_) );
NAND3X1 NAND3X1_59 ( .A(_586_), .B(_588_), .C(_587_), .Y(_589_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_583_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_584_) );
OAI21X1 OAI21X1_126 ( .A(_583_), .B(_584_), .C(_47__2_), .Y(_585_) );
NAND2X1 NAND2X1_127 ( .A(_585_), .B(_589_), .Y(_45__2_) );
OAI21X1 OAI21X1_127 ( .A(_586_), .B(_583_), .C(_588_), .Y(_47__3_) );
INVX1 INVX1_69 ( .A(_47__3_), .Y(_593_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_594_) );
NAND2X1 NAND2X1_128 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_595_) );
NAND3X1 NAND3X1_60 ( .A(_593_), .B(_595_), .C(_594_), .Y(_596_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_590_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_591_) );
OAI21X1 OAI21X1_128 ( .A(_590_), .B(_591_), .C(_47__3_), .Y(_592_) );
NAND2X1 NAND2X1_129 ( .A(_592_), .B(_596_), .Y(_45__3_) );
OAI21X1 OAI21X1_129 ( .A(_593_), .B(_590_), .C(_595_), .Y(_43_) );
INVX1 INVX1_70 ( .A(1'b1), .Y(_600_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_601_) );
NAND2X1 NAND2X1_130 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_602_) );
NAND3X1 NAND3X1_61 ( .A(_600_), .B(_602_), .C(_601_), .Y(_603_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_597_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_598_) );
OAI21X1 OAI21X1_130 ( .A(_597_), .B(_598_), .C(1'b1), .Y(_599_) );
NAND2X1 NAND2X1_131 ( .A(_599_), .B(_603_), .Y(_46__0_) );
OAI21X1 OAI21X1_131 ( .A(_600_), .B(_597_), .C(_602_), .Y(_48__1_) );
INVX1 INVX1_71 ( .A(_48__1_), .Y(_607_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_608_) );
NAND2X1 NAND2X1_132 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_609_) );
NAND3X1 NAND3X1_62 ( .A(_607_), .B(_609_), .C(_608_), .Y(_610_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_604_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_605_) );
OAI21X1 OAI21X1_132 ( .A(_604_), .B(_605_), .C(_48__1_), .Y(_606_) );
NAND2X1 NAND2X1_133 ( .A(_606_), .B(_610_), .Y(_46__1_) );
OAI21X1 OAI21X1_133 ( .A(_607_), .B(_604_), .C(_609_), .Y(_48__2_) );
INVX1 INVX1_72 ( .A(_48__2_), .Y(_614_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_615_) );
NAND2X1 NAND2X1_134 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_616_) );
NAND3X1 NAND3X1_63 ( .A(_614_), .B(_616_), .C(_615_), .Y(_617_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_611_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_612_) );
OAI21X1 OAI21X1_134 ( .A(_611_), .B(_612_), .C(_48__2_), .Y(_613_) );
NAND2X1 NAND2X1_135 ( .A(_613_), .B(_617_), .Y(_46__2_) );
OAI21X1 OAI21X1_135 ( .A(_614_), .B(_611_), .C(_616_), .Y(_48__3_) );
INVX1 INVX1_73 ( .A(_48__3_), .Y(_621_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_622_) );
NAND2X1 NAND2X1_136 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_623_) );
NAND3X1 NAND3X1_64 ( .A(_621_), .B(_623_), .C(_622_), .Y(_624_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_618_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_619_) );
OAI21X1 OAI21X1_136 ( .A(_618_), .B(_619_), .C(_48__3_), .Y(_620_) );
NAND2X1 NAND2X1_137 ( .A(_620_), .B(_624_), .Y(_46__3_) );
OAI21X1 OAI21X1_137 ( .A(_621_), .B(_618_), .C(_623_), .Y(_44_) );
INVX1 INVX1_74 ( .A(1'b0), .Y(_628_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_629_) );
NAND2X1 NAND2X1_138 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_630_) );
NAND3X1 NAND3X1_65 ( .A(_628_), .B(_630_), .C(_629_), .Y(_631_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_625_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_626_) );
OAI21X1 OAI21X1_138 ( .A(_625_), .B(_626_), .C(1'b0), .Y(_627_) );
NAND2X1 NAND2X1_139 ( .A(_627_), .B(_631_), .Y(_51__0_) );
OAI21X1 OAI21X1_139 ( .A(_628_), .B(_625_), .C(_630_), .Y(_53__1_) );
INVX1 INVX1_75 ( .A(_53__1_), .Y(_635_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_636_) );
NAND2X1 NAND2X1_140 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_637_) );
NAND3X1 NAND3X1_66 ( .A(_635_), .B(_637_), .C(_636_), .Y(_638_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_632_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_633_) );
OAI21X1 OAI21X1_140 ( .A(_632_), .B(_633_), .C(_53__1_), .Y(_634_) );
NAND2X1 NAND2X1_141 ( .A(_634_), .B(_638_), .Y(_51__1_) );
OAI21X1 OAI21X1_141 ( .A(_635_), .B(_632_), .C(_637_), .Y(_53__2_) );
INVX1 INVX1_76 ( .A(_53__2_), .Y(_642_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_643_) );
NAND2X1 NAND2X1_142 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_644_) );
NAND3X1 NAND3X1_67 ( .A(_642_), .B(_644_), .C(_643_), .Y(_645_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_639_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_640_) );
OAI21X1 OAI21X1_142 ( .A(_639_), .B(_640_), .C(_53__2_), .Y(_641_) );
NAND2X1 NAND2X1_143 ( .A(_641_), .B(_645_), .Y(_51__2_) );
OAI21X1 OAI21X1_143 ( .A(_642_), .B(_639_), .C(_644_), .Y(_53__3_) );
INVX1 INVX1_77 ( .A(_53__3_), .Y(_649_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_650_) );
NAND2X1 NAND2X1_144 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_651_) );
NAND3X1 NAND3X1_68 ( .A(_649_), .B(_651_), .C(_650_), .Y(_652_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_646_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_647_) );
OAI21X1 OAI21X1_144 ( .A(_646_), .B(_647_), .C(_53__3_), .Y(_648_) );
NAND2X1 NAND2X1_145 ( .A(_648_), .B(_652_), .Y(_51__3_) );
OAI21X1 OAI21X1_145 ( .A(_649_), .B(_646_), .C(_651_), .Y(_49_) );
INVX1 INVX1_78 ( .A(1'b1), .Y(_656_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_657_) );
NAND2X1 NAND2X1_146 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_658_) );
NAND3X1 NAND3X1_69 ( .A(_656_), .B(_658_), .C(_657_), .Y(_659_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_653_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_654_) );
OAI21X1 OAI21X1_146 ( .A(_653_), .B(_654_), .C(1'b1), .Y(_655_) );
NAND2X1 NAND2X1_147 ( .A(_655_), .B(_659_), .Y(_52__0_) );
OAI21X1 OAI21X1_147 ( .A(_656_), .B(_653_), .C(_658_), .Y(_54__1_) );
INVX1 INVX1_79 ( .A(_54__1_), .Y(_663_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_664_) );
NAND2X1 NAND2X1_148 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_665_) );
NAND3X1 NAND3X1_70 ( .A(_663_), .B(_665_), .C(_664_), .Y(_666_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_660_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_661_) );
OAI21X1 OAI21X1_148 ( .A(_660_), .B(_661_), .C(_54__1_), .Y(_662_) );
NAND2X1 NAND2X1_149 ( .A(_662_), .B(_666_), .Y(_52__1_) );
OAI21X1 OAI21X1_149 ( .A(_663_), .B(_660_), .C(_665_), .Y(_54__2_) );
INVX1 INVX1_80 ( .A(_54__2_), .Y(_670_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_671_) );
NAND2X1 NAND2X1_150 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_672_) );
NAND3X1 NAND3X1_71 ( .A(_670_), .B(_672_), .C(_671_), .Y(_673_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_667_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_668_) );
OAI21X1 OAI21X1_150 ( .A(_667_), .B(_668_), .C(_54__2_), .Y(_669_) );
NAND2X1 NAND2X1_151 ( .A(_669_), .B(_673_), .Y(_52__2_) );
OAI21X1 OAI21X1_151 ( .A(_670_), .B(_667_), .C(_672_), .Y(_54__3_) );
INVX1 INVX1_81 ( .A(_54__3_), .Y(_677_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_678_) );
NAND2X1 NAND2X1_152 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_679_) );
NAND3X1 NAND3X1_72 ( .A(_677_), .B(_679_), .C(_678_), .Y(_680_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_674_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_675_) );
OAI21X1 OAI21X1_152 ( .A(_674_), .B(_675_), .C(_54__3_), .Y(_676_) );
NAND2X1 NAND2X1_153 ( .A(_676_), .B(_680_), .Y(_52__3_) );
OAI21X1 OAI21X1_153 ( .A(_677_), .B(_674_), .C(_679_), .Y(_50_) );
INVX1 INVX1_82 ( .A(1'b0), .Y(_684_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_685_) );
NAND2X1 NAND2X1_154 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_686_) );
NAND3X1 NAND3X1_73 ( .A(_684_), .B(_686_), .C(_685_), .Y(_687_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_681_) );
AND2X2 AND2X2_73 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_682_) );
OAI21X1 OAI21X1_154 ( .A(_681_), .B(_682_), .C(1'b0), .Y(_683_) );
NAND2X1 NAND2X1_155 ( .A(_683_), .B(_687_), .Y(_57__0_) );
OAI21X1 OAI21X1_155 ( .A(_684_), .B(_681_), .C(_686_), .Y(_59__1_) );
INVX1 INVX1_83 ( .A(_59__1_), .Y(_691_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_692_) );
NAND2X1 NAND2X1_156 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_693_) );
NAND3X1 NAND3X1_74 ( .A(_691_), .B(_693_), .C(_692_), .Y(_694_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_688_) );
AND2X2 AND2X2_74 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_689_) );
OAI21X1 OAI21X1_156 ( .A(_688_), .B(_689_), .C(_59__1_), .Y(_690_) );
NAND2X1 NAND2X1_157 ( .A(_690_), .B(_694_), .Y(_57__1_) );
OAI21X1 OAI21X1_157 ( .A(_691_), .B(_688_), .C(_693_), .Y(_59__2_) );
INVX1 INVX1_84 ( .A(_59__2_), .Y(_698_) );
OR2X2 OR2X2_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_699_) );
NAND2X1 NAND2X1_158 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_700_) );
NAND3X1 NAND3X1_75 ( .A(_698_), .B(_700_), .C(_699_), .Y(_701_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_695_) );
AND2X2 AND2X2_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_696_) );
OAI21X1 OAI21X1_158 ( .A(_695_), .B(_696_), .C(_59__2_), .Y(_697_) );
NAND2X1 NAND2X1_159 ( .A(_697_), .B(_701_), .Y(_57__2_) );
OAI21X1 OAI21X1_159 ( .A(_698_), .B(_695_), .C(_700_), .Y(_59__3_) );
INVX1 INVX1_85 ( .A(_59__3_), .Y(_705_) );
OR2X2 OR2X2_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_706_) );
NAND2X1 NAND2X1_160 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_707_) );
NAND3X1 NAND3X1_76 ( .A(_705_), .B(_707_), .C(_706_), .Y(_708_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_702_) );
AND2X2 AND2X2_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_703_) );
OAI21X1 OAI21X1_160 ( .A(_702_), .B(_703_), .C(_59__3_), .Y(_704_) );
NAND2X1 NAND2X1_161 ( .A(_704_), .B(_708_), .Y(_57__3_) );
OAI21X1 OAI21X1_161 ( .A(_705_), .B(_702_), .C(_707_), .Y(_55_) );
INVX1 INVX1_86 ( .A(1'b1), .Y(_712_) );
OR2X2 OR2X2_77 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_713_) );
NAND2X1 NAND2X1_162 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_714_) );
NAND3X1 NAND3X1_77 ( .A(_712_), .B(_714_), .C(_713_), .Y(_715_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_709_) );
AND2X2 AND2X2_77 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_710_) );
OAI21X1 OAI21X1_162 ( .A(_709_), .B(_710_), .C(1'b1), .Y(_711_) );
NAND2X1 NAND2X1_163 ( .A(_711_), .B(_715_), .Y(_58__0_) );
OAI21X1 OAI21X1_163 ( .A(_712_), .B(_709_), .C(_714_), .Y(_60__1_) );
INVX1 INVX1_87 ( .A(_60__1_), .Y(_719_) );
OR2X2 OR2X2_78 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_720_) );
NAND2X1 NAND2X1_164 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_721_) );
NAND3X1 NAND3X1_78 ( .A(_719_), .B(_721_), .C(_720_), .Y(_722_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_716_) );
AND2X2 AND2X2_78 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_717_) );
OAI21X1 OAI21X1_164 ( .A(_716_), .B(_717_), .C(_60__1_), .Y(_718_) );
NAND2X1 NAND2X1_165 ( .A(_718_), .B(_722_), .Y(_58__1_) );
OAI21X1 OAI21X1_165 ( .A(_719_), .B(_716_), .C(_721_), .Y(_60__2_) );
INVX1 INVX1_88 ( .A(_60__2_), .Y(_726_) );
OR2X2 OR2X2_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_727_) );
NAND2X1 NAND2X1_166 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_728_) );
NAND3X1 NAND3X1_79 ( .A(_726_), .B(_728_), .C(_727_), .Y(_729_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_723_) );
AND2X2 AND2X2_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_724_) );
OAI21X1 OAI21X1_166 ( .A(_723_), .B(_724_), .C(_60__2_), .Y(_725_) );
NAND2X1 NAND2X1_167 ( .A(_725_), .B(_729_), .Y(_58__2_) );
OAI21X1 OAI21X1_167 ( .A(_726_), .B(_723_), .C(_728_), .Y(_60__3_) );
INVX1 INVX1_89 ( .A(_60__3_), .Y(_733_) );
OR2X2 OR2X2_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_734_) );
NAND2X1 NAND2X1_168 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_735_) );
NAND3X1 NAND3X1_80 ( .A(_733_), .B(_735_), .C(_734_), .Y(_736_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_730_) );
AND2X2 AND2X2_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_731_) );
OAI21X1 OAI21X1_168 ( .A(_730_), .B(_731_), .C(_60__3_), .Y(_732_) );
NAND2X1 NAND2X1_169 ( .A(_732_), .B(_736_), .Y(_58__3_) );
OAI21X1 OAI21X1_169 ( .A(_733_), .B(_730_), .C(_735_), .Y(_56_) );
INVX1 INVX1_90 ( .A(1'b0), .Y(_740_) );
OR2X2 OR2X2_81 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_741_) );
NAND2X1 NAND2X1_170 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_742_) );
NAND3X1 NAND3X1_81 ( .A(_740_), .B(_742_), .C(_741_), .Y(_743_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_737_) );
AND2X2 AND2X2_81 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_738_) );
OAI21X1 OAI21X1_170 ( .A(_737_), .B(_738_), .C(1'b0), .Y(_739_) );
NAND2X1 NAND2X1_171 ( .A(_739_), .B(_743_), .Y(_63__0_) );
OAI21X1 OAI21X1_171 ( .A(_740_), .B(_737_), .C(_742_), .Y(_65__1_) );
INVX1 INVX1_91 ( .A(_65__1_), .Y(_747_) );
OR2X2 OR2X2_82 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_748_) );
NAND2X1 NAND2X1_172 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_749_) );
NAND3X1 NAND3X1_82 ( .A(_747_), .B(_749_), .C(_748_), .Y(_750_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_744_) );
AND2X2 AND2X2_82 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_745_) );
OAI21X1 OAI21X1_172 ( .A(_744_), .B(_745_), .C(_65__1_), .Y(_746_) );
NAND2X1 NAND2X1_173 ( .A(_746_), .B(_750_), .Y(_63__1_) );
OAI21X1 OAI21X1_173 ( .A(_747_), .B(_744_), .C(_749_), .Y(_65__2_) );
INVX1 INVX1_92 ( .A(_65__2_), .Y(_754_) );
OR2X2 OR2X2_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_755_) );
NAND2X1 NAND2X1_174 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_756_) );
NAND3X1 NAND3X1_83 ( .A(_754_), .B(_756_), .C(_755_), .Y(_757_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_751_) );
AND2X2 AND2X2_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_752_) );
OAI21X1 OAI21X1_174 ( .A(_751_), .B(_752_), .C(_65__2_), .Y(_753_) );
NAND2X1 NAND2X1_175 ( .A(_753_), .B(_757_), .Y(_63__2_) );
OAI21X1 OAI21X1_175 ( .A(_754_), .B(_751_), .C(_756_), .Y(_65__3_) );
INVX1 INVX1_93 ( .A(_65__3_), .Y(_761_) );
OR2X2 OR2X2_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_762_) );
NAND2X1 NAND2X1_176 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_763_) );
NAND3X1 NAND3X1_84 ( .A(_761_), .B(_763_), .C(_762_), .Y(_764_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_758_) );
AND2X2 AND2X2_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_759_) );
OAI21X1 OAI21X1_176 ( .A(_758_), .B(_759_), .C(_65__3_), .Y(_760_) );
NAND2X1 NAND2X1_177 ( .A(_760_), .B(_764_), .Y(_63__3_) );
OAI21X1 OAI21X1_177 ( .A(_761_), .B(_758_), .C(_763_), .Y(_61_) );
INVX1 INVX1_94 ( .A(1'b1), .Y(_768_) );
OR2X2 OR2X2_85 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_769_) );
NAND2X1 NAND2X1_178 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_770_) );
NAND3X1 NAND3X1_85 ( .A(_768_), .B(_770_), .C(_769_), .Y(_771_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_765_) );
AND2X2 AND2X2_85 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_766_) );
OAI21X1 OAI21X1_178 ( .A(_765_), .B(_766_), .C(1'b1), .Y(_767_) );
NAND2X1 NAND2X1_179 ( .A(_767_), .B(_771_), .Y(_64__0_) );
OAI21X1 OAI21X1_179 ( .A(_768_), .B(_765_), .C(_770_), .Y(_66__1_) );
INVX1 INVX1_95 ( .A(_66__1_), .Y(_775_) );
OR2X2 OR2X2_86 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_776_) );
NAND2X1 NAND2X1_180 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_777_) );
NAND3X1 NAND3X1_86 ( .A(_775_), .B(_777_), .C(_776_), .Y(_778_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_772_) );
AND2X2 AND2X2_86 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_773_) );
OAI21X1 OAI21X1_180 ( .A(_772_), .B(_773_), .C(_66__1_), .Y(_774_) );
NAND2X1 NAND2X1_181 ( .A(_774_), .B(_778_), .Y(_64__1_) );
OAI21X1 OAI21X1_181 ( .A(_775_), .B(_772_), .C(_777_), .Y(_66__2_) );
INVX1 INVX1_96 ( .A(_66__2_), .Y(_782_) );
OR2X2 OR2X2_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_783_) );
NAND2X1 NAND2X1_182 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_784_) );
NAND3X1 NAND3X1_87 ( .A(_782_), .B(_784_), .C(_783_), .Y(_785_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_779_) );
AND2X2 AND2X2_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_780_) );
OAI21X1 OAI21X1_182 ( .A(_779_), .B(_780_), .C(_66__2_), .Y(_781_) );
NAND2X1 NAND2X1_183 ( .A(_781_), .B(_785_), .Y(_64__2_) );
OAI21X1 OAI21X1_183 ( .A(_782_), .B(_779_), .C(_784_), .Y(_66__3_) );
INVX1 INVX1_97 ( .A(_66__3_), .Y(_789_) );
OR2X2 OR2X2_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_790_) );
NAND2X1 NAND2X1_184 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_791_) );
NAND3X1 NAND3X1_88 ( .A(_789_), .B(_791_), .C(_790_), .Y(_792_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_786_) );
AND2X2 AND2X2_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_787_) );
OAI21X1 OAI21X1_184 ( .A(_786_), .B(_787_), .C(_66__3_), .Y(_788_) );
NAND2X1 NAND2X1_185 ( .A(_788_), .B(_792_), .Y(_64__3_) );
OAI21X1 OAI21X1_185 ( .A(_789_), .B(_786_), .C(_791_), .Y(_62_) );
INVX1 INVX1_98 ( .A(1'b0), .Y(_796_) );
OR2X2 OR2X2_89 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_797_) );
NAND2X1 NAND2X1_186 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_798_) );
NAND3X1 NAND3X1_89 ( .A(_796_), .B(_798_), .C(_797_), .Y(_799_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_793_) );
AND2X2 AND2X2_89 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_794_) );
OAI21X1 OAI21X1_186 ( .A(_793_), .B(_794_), .C(1'b0), .Y(_795_) );
NAND2X1 NAND2X1_187 ( .A(_795_), .B(_799_), .Y(_0__0_) );
OAI21X1 OAI21X1_187 ( .A(_796_), .B(_793_), .C(_798_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_99 ( .A(rca_inst_w_CARRY_1_), .Y(_803_) );
OR2X2 OR2X2_90 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_804_) );
NAND2X1 NAND2X1_188 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_805_) );
NAND3X1 NAND3X1_90 ( .A(_803_), .B(_805_), .C(_804_), .Y(_806_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_800_) );
AND2X2 AND2X2_90 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_801_) );
OAI21X1 OAI21X1_188 ( .A(_800_), .B(_801_), .C(rca_inst_w_CARRY_1_), .Y(_802_) );
NAND2X1 NAND2X1_189 ( .A(_802_), .B(_806_), .Y(_0__1_) );
OAI21X1 OAI21X1_189 ( .A(_803_), .B(_800_), .C(_805_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_100 ( .A(rca_inst_w_CARRY_2_), .Y(_810_) );
OR2X2 OR2X2_91 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_811_) );
NAND2X1 NAND2X1_190 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_812_) );
NAND3X1 NAND3X1_91 ( .A(_810_), .B(_812_), .C(_811_), .Y(_813_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_807_) );
AND2X2 AND2X2_91 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_808_) );
OAI21X1 OAI21X1_190 ( .A(_807_), .B(_808_), .C(rca_inst_w_CARRY_2_), .Y(_809_) );
NAND2X1 NAND2X1_191 ( .A(_809_), .B(_813_), .Y(_0__2_) );
BUFX2 BUFX2_1 ( .A(w_cout_11_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
INVX1 INVX1_101 ( .A(_1_), .Y(_67_) );
NAND2X1 NAND2X1_192 ( .A(_2_), .B(1'b0), .Y(_68_) );
OAI21X1 OAI21X1_191 ( .A(1'b0), .B(_67_), .C(_68_), .Y(w_cout_1_) );
INVX1 INVX1_102 ( .A(_3__0_), .Y(_69_) );
NAND2X1 NAND2X1_193 ( .A(_4__0_), .B(1'b0), .Y(_70_) );
OAI21X1 OAI21X1_192 ( .A(1'b0), .B(_69_), .C(_70_), .Y(_0__3_) );
INVX1 INVX1_103 ( .A(_3__1_), .Y(_71_) );
NAND2X1 NAND2X1_194 ( .A(1'b0), .B(_4__1_), .Y(_72_) );
OAI21X1 OAI21X1_193 ( .A(1'b0), .B(_71_), .C(_72_), .Y(_0__4_) );
INVX1 INVX1_104 ( .A(_3__2_), .Y(_73_) );
NAND2X1 NAND2X1_195 ( .A(1'b0), .B(_4__2_), .Y(_74_) );
OAI21X1 OAI21X1_194 ( .A(1'b0), .B(_73_), .C(_74_), .Y(_0__5_) );
INVX1 INVX1_105 ( .A(_3__3_), .Y(_75_) );
NAND2X1 NAND2X1_196 ( .A(1'b0), .B(_4__3_), .Y(_76_) );
OAI21X1 OAI21X1_195 ( .A(1'b0), .B(_75_), .C(_76_), .Y(_0__6_) );
INVX1 INVX1_106 ( .A(_7_), .Y(_77_) );
NAND2X1 NAND2X1_197 ( .A(_8_), .B(w_cout_1_), .Y(_78_) );
OAI21X1 OAI21X1_196 ( .A(w_cout_1_), .B(_77_), .C(_78_), .Y(w_cout_2_) );
INVX1 INVX1_107 ( .A(_9__0_), .Y(_79_) );
NAND2X1 NAND2X1_198 ( .A(_10__0_), .B(w_cout_1_), .Y(_80_) );
OAI21X1 OAI21X1_197 ( .A(w_cout_1_), .B(_79_), .C(_80_), .Y(_0__7_) );
INVX1 INVX1_108 ( .A(_9__1_), .Y(_81_) );
NAND2X1 NAND2X1_199 ( .A(w_cout_1_), .B(_10__1_), .Y(_82_) );
OAI21X1 OAI21X1_198 ( .A(w_cout_1_), .B(_81_), .C(_82_), .Y(_0__8_) );
INVX1 INVX1_109 ( .A(_9__2_), .Y(_83_) );
NAND2X1 NAND2X1_200 ( .A(w_cout_1_), .B(_10__2_), .Y(_84_) );
OAI21X1 OAI21X1_199 ( .A(w_cout_1_), .B(_83_), .C(_84_), .Y(_0__9_) );
INVX1 INVX1_110 ( .A(_9__3_), .Y(_85_) );
NAND2X1 NAND2X1_201 ( .A(w_cout_1_), .B(_10__3_), .Y(_86_) );
OAI21X1 OAI21X1_200 ( .A(w_cout_1_), .B(_85_), .C(_86_), .Y(_0__10_) );
INVX1 INVX1_111 ( .A(_13_), .Y(_87_) );
NAND2X1 NAND2X1_202 ( .A(_14_), .B(w_cout_2_), .Y(_88_) );
OAI21X1 OAI21X1_201 ( .A(w_cout_2_), .B(_87_), .C(_88_), .Y(w_cout_3_) );
INVX1 INVX1_112 ( .A(_15__0_), .Y(_89_) );
NAND2X1 NAND2X1_203 ( .A(_16__0_), .B(w_cout_2_), .Y(_90_) );
OAI21X1 OAI21X1_202 ( .A(w_cout_2_), .B(_89_), .C(_90_), .Y(_0__11_) );
INVX1 INVX1_113 ( .A(_15__1_), .Y(_91_) );
NAND2X1 NAND2X1_204 ( .A(w_cout_2_), .B(_16__1_), .Y(_92_) );
OAI21X1 OAI21X1_203 ( .A(w_cout_2_), .B(_91_), .C(_92_), .Y(_0__12_) );
INVX1 INVX1_114 ( .A(_15__2_), .Y(_93_) );
NAND2X1 NAND2X1_205 ( .A(w_cout_2_), .B(_16__2_), .Y(_94_) );
OAI21X1 OAI21X1_204 ( .A(w_cout_2_), .B(_93_), .C(_94_), .Y(_0__13_) );
INVX1 INVX1_115 ( .A(_15__3_), .Y(_95_) );
NAND2X1 NAND2X1_206 ( .A(w_cout_2_), .B(_16__3_), .Y(_96_) );
OAI21X1 OAI21X1_205 ( .A(w_cout_2_), .B(_95_), .C(_96_), .Y(_0__14_) );
INVX1 INVX1_116 ( .A(_19_), .Y(_97_) );
NAND2X1 NAND2X1_207 ( .A(_20_), .B(w_cout_3_), .Y(_98_) );
OAI21X1 OAI21X1_206 ( .A(w_cout_3_), .B(_97_), .C(_98_), .Y(w_cout_4_) );
INVX1 INVX1_117 ( .A(_21__0_), .Y(_99_) );
NAND2X1 NAND2X1_208 ( .A(_22__0_), .B(w_cout_3_), .Y(_100_) );
OAI21X1 OAI21X1_207 ( .A(w_cout_3_), .B(_99_), .C(_100_), .Y(_0__15_) );
INVX1 INVX1_118 ( .A(_21__1_), .Y(_101_) );
NAND2X1 NAND2X1_209 ( .A(w_cout_3_), .B(_22__1_), .Y(_102_) );
OAI21X1 OAI21X1_208 ( .A(w_cout_3_), .B(_101_), .C(_102_), .Y(_0__16_) );
INVX1 INVX1_119 ( .A(_21__2_), .Y(_103_) );
NAND2X1 NAND2X1_210 ( .A(w_cout_3_), .B(_22__2_), .Y(_104_) );
OAI21X1 OAI21X1_209 ( .A(w_cout_3_), .B(_103_), .C(_104_), .Y(_0__17_) );
INVX1 INVX1_120 ( .A(_21__3_), .Y(_105_) );
NAND2X1 NAND2X1_211 ( .A(w_cout_3_), .B(_22__3_), .Y(_106_) );
OAI21X1 OAI21X1_210 ( .A(w_cout_3_), .B(_105_), .C(_106_), .Y(_0__18_) );
INVX1 INVX1_121 ( .A(_25_), .Y(_107_) );
NAND2X1 NAND2X1_212 ( .A(_26_), .B(w_cout_4_), .Y(_108_) );
OAI21X1 OAI21X1_211 ( .A(w_cout_4_), .B(_107_), .C(_108_), .Y(w_cout_5_) );
INVX1 INVX1_122 ( .A(_27__0_), .Y(_109_) );
NAND2X1 NAND2X1_213 ( .A(_28__0_), .B(w_cout_4_), .Y(_110_) );
OAI21X1 OAI21X1_212 ( .A(w_cout_4_), .B(_109_), .C(_110_), .Y(_0__19_) );
INVX1 INVX1_123 ( .A(_27__1_), .Y(_111_) );
NAND2X1 NAND2X1_214 ( .A(w_cout_4_), .B(_28__1_), .Y(_112_) );
OAI21X1 OAI21X1_213 ( .A(w_cout_4_), .B(_111_), .C(_112_), .Y(_0__20_) );
INVX1 INVX1_124 ( .A(_27__2_), .Y(_113_) );
NAND2X1 NAND2X1_215 ( .A(w_cout_4_), .B(_28__2_), .Y(_114_) );
OAI21X1 OAI21X1_214 ( .A(w_cout_4_), .B(_113_), .C(_114_), .Y(_0__21_) );
INVX1 INVX1_125 ( .A(_27__3_), .Y(_115_) );
NAND2X1 NAND2X1_216 ( .A(w_cout_4_), .B(_28__3_), .Y(_116_) );
OAI21X1 OAI21X1_215 ( .A(w_cout_4_), .B(_115_), .C(_116_), .Y(_0__22_) );
INVX1 INVX1_126 ( .A(_31_), .Y(_117_) );
NAND2X1 NAND2X1_217 ( .A(_32_), .B(w_cout_5_), .Y(_118_) );
OAI21X1 OAI21X1_216 ( .A(w_cout_5_), .B(_117_), .C(_118_), .Y(w_cout_6_) );
INVX1 INVX1_127 ( .A(_33__0_), .Y(_119_) );
NAND2X1 NAND2X1_218 ( .A(_34__0_), .B(w_cout_5_), .Y(_120_) );
OAI21X1 OAI21X1_217 ( .A(w_cout_5_), .B(_119_), .C(_120_), .Y(_0__23_) );
INVX1 INVX1_128 ( .A(_33__1_), .Y(_121_) );
NAND2X1 NAND2X1_219 ( .A(w_cout_5_), .B(_34__1_), .Y(_122_) );
OAI21X1 OAI21X1_218 ( .A(w_cout_5_), .B(_121_), .C(_122_), .Y(_0__24_) );
INVX1 INVX1_129 ( .A(_33__2_), .Y(_123_) );
NAND2X1 NAND2X1_220 ( .A(w_cout_5_), .B(_34__2_), .Y(_124_) );
OAI21X1 OAI21X1_219 ( .A(w_cout_5_), .B(_123_), .C(_124_), .Y(_0__25_) );
INVX1 INVX1_130 ( .A(_33__3_), .Y(_125_) );
NAND2X1 NAND2X1_221 ( .A(w_cout_5_), .B(_34__3_), .Y(_126_) );
OAI21X1 OAI21X1_220 ( .A(w_cout_5_), .B(_125_), .C(_126_), .Y(_0__26_) );
INVX1 INVX1_131 ( .A(_37_), .Y(_127_) );
NAND2X1 NAND2X1_222 ( .A(_38_), .B(w_cout_6_), .Y(_128_) );
OAI21X1 OAI21X1_221 ( .A(w_cout_6_), .B(_127_), .C(_128_), .Y(w_cout_7_) );
INVX1 INVX1_132 ( .A(_39__0_), .Y(_129_) );
NAND2X1 NAND2X1_223 ( .A(_40__0_), .B(w_cout_6_), .Y(_130_) );
OAI21X1 OAI21X1_222 ( .A(w_cout_6_), .B(_129_), .C(_130_), .Y(_0__27_) );
INVX1 INVX1_133 ( .A(_39__1_), .Y(_131_) );
NAND2X1 NAND2X1_224 ( .A(w_cout_6_), .B(_40__1_), .Y(_132_) );
OAI21X1 OAI21X1_223 ( .A(w_cout_6_), .B(_131_), .C(_132_), .Y(_0__28_) );
INVX1 INVX1_134 ( .A(_39__2_), .Y(_133_) );
NAND2X1 NAND2X1_225 ( .A(w_cout_6_), .B(_40__2_), .Y(_134_) );
OAI21X1 OAI21X1_224 ( .A(w_cout_6_), .B(_133_), .C(_134_), .Y(_0__29_) );
INVX1 INVX1_135 ( .A(_39__3_), .Y(_135_) );
NAND2X1 NAND2X1_226 ( .A(w_cout_6_), .B(_40__3_), .Y(_136_) );
OAI21X1 OAI21X1_225 ( .A(w_cout_6_), .B(_135_), .C(_136_), .Y(_0__30_) );
INVX1 INVX1_136 ( .A(_43_), .Y(_137_) );
NAND2X1 NAND2X1_227 ( .A(_44_), .B(w_cout_7_), .Y(_138_) );
OAI21X1 OAI21X1_226 ( .A(w_cout_7_), .B(_137_), .C(_138_), .Y(w_cout_8_) );
INVX1 INVX1_137 ( .A(_45__0_), .Y(_139_) );
NAND2X1 NAND2X1_228 ( .A(_46__0_), .B(w_cout_7_), .Y(_140_) );
OAI21X1 OAI21X1_227 ( .A(w_cout_7_), .B(_139_), .C(_140_), .Y(_0__31_) );
INVX1 INVX1_138 ( .A(_45__1_), .Y(_141_) );
NAND2X1 NAND2X1_229 ( .A(w_cout_7_), .B(_46__1_), .Y(_142_) );
OAI21X1 OAI21X1_228 ( .A(w_cout_7_), .B(_141_), .C(_142_), .Y(_0__32_) );
INVX1 INVX1_139 ( .A(_45__2_), .Y(_143_) );
NAND2X1 NAND2X1_230 ( .A(w_cout_7_), .B(_46__2_), .Y(_144_) );
OAI21X1 OAI21X1_229 ( .A(w_cout_7_), .B(_143_), .C(_144_), .Y(_0__33_) );
INVX1 INVX1_140 ( .A(_45__3_), .Y(_145_) );
NAND2X1 NAND2X1_231 ( .A(w_cout_7_), .B(_46__3_), .Y(_146_) );
OAI21X1 OAI21X1_230 ( .A(w_cout_7_), .B(_145_), .C(_146_), .Y(_0__34_) );
INVX1 INVX1_141 ( .A(_49_), .Y(_147_) );
NAND2X1 NAND2X1_232 ( .A(_50_), .B(w_cout_8_), .Y(_148_) );
OAI21X1 OAI21X1_231 ( .A(w_cout_8_), .B(_147_), .C(_148_), .Y(w_cout_9_) );
INVX1 INVX1_142 ( .A(_51__0_), .Y(_149_) );
NAND2X1 NAND2X1_233 ( .A(_52__0_), .B(w_cout_8_), .Y(_150_) );
OAI21X1 OAI21X1_232 ( .A(w_cout_8_), .B(_149_), .C(_150_), .Y(_0__35_) );
INVX1 INVX1_143 ( .A(_51__1_), .Y(_151_) );
NAND2X1 NAND2X1_234 ( .A(w_cout_8_), .B(_52__1_), .Y(_152_) );
OAI21X1 OAI21X1_233 ( .A(w_cout_8_), .B(_151_), .C(_152_), .Y(_0__36_) );
INVX1 INVX1_144 ( .A(_51__2_), .Y(_153_) );
NAND2X1 NAND2X1_235 ( .A(w_cout_8_), .B(_52__2_), .Y(_154_) );
OAI21X1 OAI21X1_234 ( .A(w_cout_8_), .B(_153_), .C(_154_), .Y(_0__37_) );
INVX1 INVX1_145 ( .A(_51__3_), .Y(_155_) );
NAND2X1 NAND2X1_236 ( .A(w_cout_8_), .B(_52__3_), .Y(_156_) );
OAI21X1 OAI21X1_235 ( .A(w_cout_8_), .B(_155_), .C(_156_), .Y(_0__38_) );
INVX1 INVX1_146 ( .A(_55_), .Y(_157_) );
NAND2X1 NAND2X1_237 ( .A(_56_), .B(w_cout_9_), .Y(_158_) );
OAI21X1 OAI21X1_236 ( .A(w_cout_9_), .B(_157_), .C(_158_), .Y(w_cout_10_) );
BUFX2 BUFX2_49 ( .A(1'b0), .Y(_5__0_) );
BUFX2 BUFX2_50 ( .A(_1_), .Y(_5__4_) );
BUFX2 BUFX2_51 ( .A(1'b1), .Y(_6__0_) );
BUFX2 BUFX2_52 ( .A(_2_), .Y(_6__4_) );
BUFX2 BUFX2_53 ( .A(1'b0), .Y(_11__0_) );
BUFX2 BUFX2_54 ( .A(_7_), .Y(_11__4_) );
BUFX2 BUFX2_55 ( .A(1'b1), .Y(_12__0_) );
BUFX2 BUFX2_56 ( .A(_8_), .Y(_12__4_) );
BUFX2 BUFX2_57 ( .A(1'b0), .Y(_17__0_) );
BUFX2 BUFX2_58 ( .A(_13_), .Y(_17__4_) );
BUFX2 BUFX2_59 ( .A(1'b1), .Y(_18__0_) );
BUFX2 BUFX2_60 ( .A(_14_), .Y(_18__4_) );
BUFX2 BUFX2_61 ( .A(1'b0), .Y(_23__0_) );
BUFX2 BUFX2_62 ( .A(_19_), .Y(_23__4_) );
BUFX2 BUFX2_63 ( .A(1'b1), .Y(_24__0_) );
BUFX2 BUFX2_64 ( .A(_20_), .Y(_24__4_) );
BUFX2 BUFX2_65 ( .A(1'b0), .Y(_29__0_) );
BUFX2 BUFX2_66 ( .A(_25_), .Y(_29__4_) );
BUFX2 BUFX2_67 ( .A(1'b1), .Y(_30__0_) );
BUFX2 BUFX2_68 ( .A(_26_), .Y(_30__4_) );
BUFX2 BUFX2_69 ( .A(1'b0), .Y(_35__0_) );
BUFX2 BUFX2_70 ( .A(_31_), .Y(_35__4_) );
BUFX2 BUFX2_71 ( .A(1'b1), .Y(_36__0_) );
BUFX2 BUFX2_72 ( .A(_32_), .Y(_36__4_) );
BUFX2 BUFX2_73 ( .A(1'b0), .Y(_41__0_) );
BUFX2 BUFX2_74 ( .A(_37_), .Y(_41__4_) );
BUFX2 BUFX2_75 ( .A(1'b1), .Y(_42__0_) );
BUFX2 BUFX2_76 ( .A(_38_), .Y(_42__4_) );
BUFX2 BUFX2_77 ( .A(1'b0), .Y(_47__0_) );
BUFX2 BUFX2_78 ( .A(_43_), .Y(_47__4_) );
BUFX2 BUFX2_79 ( .A(1'b1), .Y(_48__0_) );
BUFX2 BUFX2_80 ( .A(_44_), .Y(_48__4_) );
BUFX2 BUFX2_81 ( .A(1'b0), .Y(_53__0_) );
BUFX2 BUFX2_82 ( .A(_49_), .Y(_53__4_) );
BUFX2 BUFX2_83 ( .A(1'b1), .Y(_54__0_) );
BUFX2 BUFX2_84 ( .A(_50_), .Y(_54__4_) );
BUFX2 BUFX2_85 ( .A(1'b0), .Y(_59__0_) );
BUFX2 BUFX2_86 ( .A(_55_), .Y(_59__4_) );
BUFX2 BUFX2_87 ( .A(1'b1), .Y(_60__0_) );
BUFX2 BUFX2_88 ( .A(_56_), .Y(_60__4_) );
BUFX2 BUFX2_89 ( .A(1'b0), .Y(_65__0_) );
BUFX2 BUFX2_90 ( .A(_61_), .Y(_65__4_) );
BUFX2 BUFX2_91 ( .A(1'b1), .Y(_66__0_) );
BUFX2 BUFX2_92 ( .A(_62_), .Y(_66__4_) );
BUFX2 BUFX2_93 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_94 ( .A(1'b0), .Y(w_cout_0_) );
endmodule
