module cla_4bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [3:0] i_add1;
input [3:0] i_add2;
output [4:0] o_result;

NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_0_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_1_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_1_), .Y(w_C_2_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_2_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_3_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_1_), .C(_3_), .Y(_4_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_2_), .Y(w_C_3_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_5_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_6_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(_6_), .C(_4_), .Y(_7_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_7_), .Y(w_C_4_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_8_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_8_), .Y(w_C_1_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_9__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_9__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_9__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_9__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(o_result[4]) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_13_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_14_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_15_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_15_), .C(_14_), .Y(_16_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_10_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_11_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_11_), .C(gnd), .Y(_12_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_16_), .Y(_9__0_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_20_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_21_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_22_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_22_), .C(_21_), .Y(_23_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_17_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_18_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_18_), .C(w_C_1_), .Y(_19_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_23_), .Y(_9__1_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_27_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_28_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_29_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_29_), .C(_28_), .Y(_30_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_24_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_25_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_25_), .C(w_C_2_), .Y(_26_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_30_), .Y(_9__2_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_34_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_35_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_36_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_36_), .C(_35_), .Y(_37_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_31_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_32_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_32_), .C(w_C_3_), .Y(_33_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_37_), .Y(_9__3_) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_9__4_) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
