module cla_15bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [14:0] i_add1;
input [14:0] i_add2;
output [15:0] o_result;

NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_18_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_18_), .Y(w_C_1_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_19_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_19_), .Y(_20_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .C(_20_), .Y(_21_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_21_), .Y(w_C_2_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_22_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_23_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_24_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_24_), .C(_20_), .Y(_25_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_25_), .Y(w_C_3_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_26_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_27_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_27_), .C(_25_), .Y(_28_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_26_), .Y(w_C_4_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_29_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_30_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_30_), .C(_28_), .Y(_31_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_31_), .Y(w_C_5_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_32_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_32_), .Y(_33_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_34_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_34_), .C(_31_), .Y(_35_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_33_), .Y(w_C_6_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .Y(_36_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add1[6]), .Y(_37_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_38_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_38_), .Y(_39_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_39_), .C(_35_), .Y(_40_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_37_), .C(_40_), .Y(w_C_7_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_41_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_41_), .Y(_42_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_37_), .Y(_43_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(_44_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_45_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_45_), .Y(_46_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_46_), .C(_40_), .Y(_47_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_42_), .Y(w_C_8_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_48_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_48_), .Y(_49_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_50_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_50_), .Y(_51_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_51_), .C(_47_), .Y(_52_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_49_), .Y(_53_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_53_), .Y(w_C_9_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_54_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_54_), .Y(_55_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_56_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_53_), .C(_55_), .Y(w_C_10_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_57_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_57_), .Y(_58_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_56_), .Y(_59_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_55_), .C(_52_), .Y(_60_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_61_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_61_), .Y(_0_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_0_), .C(_60_), .Y(_1_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_58_), .Y(_2_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_2_), .Y(w_C_11_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_3_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_4_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_2_), .C(_3_), .Y(w_C_12_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .Y(_5_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add1[12]), .Y(_6_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(_7_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_3_), .C(_1_), .Y(_8_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_6_), .Y(_9_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_9_), .C(_8_), .Y(_10_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_6_), .C(_10_), .Y(w_C_13_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_11_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_12_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_13_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_13_), .C(_10_), .Y(_14_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_11_), .Y(w_C_14_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_15_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_16_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_16_), .C(_14_), .Y(_17_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_17_), .Y(w_C_15_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_62__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_62__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_62__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_62__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_62__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_62__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_62__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_62__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_62__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_62__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_62__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_62__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_62__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_62__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_62__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(o_result[15]) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_66_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_67_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_68_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_68_), .C(_67_), .Y(_69_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_63_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_64_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_64_), .C(w_C_4_), .Y(_65_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_69_), .Y(_62__4_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_73_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_74_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_75_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_75_), .C(_74_), .Y(_76_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_70_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_71_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_71_), .C(w_C_5_), .Y(_72_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_76_), .Y(_62__5_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_80_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_81_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_82_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_82_), .C(_81_), .Y(_83_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_77_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_78_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_78_), .C(w_C_6_), .Y(_79_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_83_), .Y(_62__6_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_87_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_88_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_89_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_89_), .C(_88_), .Y(_90_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_84_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_85_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_85_), .C(w_C_7_), .Y(_86_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_90_), .Y(_62__7_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_94_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_95_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_96_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_96_), .C(_95_), .Y(_97_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_91_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_92_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_92_), .C(w_C_8_), .Y(_93_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_97_), .Y(_62__8_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_101_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_102_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_103_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_103_), .C(_102_), .Y(_104_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_98_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_99_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_99_), .C(w_C_9_), .Y(_100_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_104_), .Y(_62__9_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_108_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_109_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_110_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_110_), .C(_109_), .Y(_111_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_105_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_106_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_106_), .C(w_C_10_), .Y(_107_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_111_), .Y(_62__10_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_115_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_116_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_117_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_117_), .C(_116_), .Y(_118_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_112_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_113_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_113_), .C(w_C_11_), .Y(_114_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_118_), .Y(_62__11_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(w_C_12_), .Y(_122_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_123_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_124_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_124_), .C(_123_), .Y(_125_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_119_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_120_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_120_), .C(w_C_12_), .Y(_121_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_125_), .Y(_62__12_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(w_C_13_), .Y(_129_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_130_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_131_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_129_), .B(_131_), .C(_130_), .Y(_132_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_126_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_127_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_127_), .C(w_C_13_), .Y(_128_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_132_), .Y(_62__13_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(w_C_14_), .Y(_136_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_137_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_138_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_138_), .C(_137_), .Y(_139_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_133_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_134_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_134_), .C(w_C_14_), .Y(_135_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_139_), .Y(_62__14_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_143_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_144_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_145_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_145_), .C(_144_), .Y(_146_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_140_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_141_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_141_), .C(gnd), .Y(_142_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_146_), .Y(_62__0_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_150_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_151_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_152_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_152_), .C(_151_), .Y(_153_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_147_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_148_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_148_), .C(w_C_1_), .Y(_149_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_153_), .Y(_62__1_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_157_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_158_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_159_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_159_), .C(_158_), .Y(_160_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_154_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_155_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_155_), .C(w_C_2_), .Y(_156_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_160_), .Y(_62__2_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_164_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_165_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_166_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_166_), .C(_165_), .Y(_167_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_161_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_162_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_162_), .C(w_C_3_), .Y(_163_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_167_), .Y(_62__3_) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(_62__15_) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
