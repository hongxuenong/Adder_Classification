module CSkipA_15bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_4_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
INVX1 INVX1_1 ( .A(i_add_term1[0]), .Y(_10_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[0]), .B(_10_), .Y(_11_) );
INVX1 INVX1_2 ( .A(i_add_term2[0]), .Y(_12_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term1[0]), .B(_12_), .Y(_13_) );
INVX1 INVX1_3 ( .A(i_add_term1[1]), .Y(_14_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[1]), .B(_14_), .Y(_15_) );
INVX1 INVX1_4 ( .A(i_add_term2[1]), .Y(_16_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term1[1]), .B(_16_), .Y(_17_) );
OAI22X1 OAI22X1_1 ( .A(_11_), .B(_13_), .C(_15_), .D(_17_), .Y(_18_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_19_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_20_) );
NOR2X1 NOR2X1_6 ( .A(_19_), .B(_20_), .Y(_21_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_22_) );
NAND2X1 NAND2X1_1 ( .A(_21_), .B(_22_), .Y(_23_) );
NOR2X1 NOR2X1_7 ( .A(_18_), .B(_23_), .Y(_3_) );
INVX1 INVX1_5 ( .A(_1_), .Y(_24_) );
NAND2X1 NAND2X1_2 ( .A(1'b0), .B(_3_), .Y(_25_) );
OAI21X1 OAI21X1_1 ( .A(_3_), .B(_24_), .C(_25_), .Y(w_cout_1_) );
INVX1 INVX1_6 ( .A(i_add_term1[4]), .Y(_26_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[4]), .B(_26_), .Y(_27_) );
INVX1 INVX1_7 ( .A(i_add_term2[4]), .Y(_28_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term1[4]), .B(_28_), .Y(_29_) );
INVX1 INVX1_8 ( .A(i_add_term1[5]), .Y(_30_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[5]), .B(_30_), .Y(_31_) );
INVX1 INVX1_9 ( .A(i_add_term2[5]), .Y(_32_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term1[5]), .B(_32_), .Y(_33_) );
OAI22X1 OAI22X1_2 ( .A(_27_), .B(_29_), .C(_31_), .D(_33_), .Y(_34_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_35_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_36_) );
NOR2X1 NOR2X1_13 ( .A(_35_), .B(_36_), .Y(_37_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_38_) );
NAND2X1 NAND2X1_3 ( .A(_37_), .B(_38_), .Y(_39_) );
NOR2X1 NOR2X1_14 ( .A(_34_), .B(_39_), .Y(_6_) );
INVX1 INVX1_10 ( .A(_4_), .Y(_40_) );
NAND2X1 NAND2X1_4 ( .A(1'b0), .B(_6_), .Y(_41_) );
OAI21X1 OAI21X1_2 ( .A(_6_), .B(_40_), .C(_41_), .Y(w_cout_2_) );
INVX1 INVX1_11 ( .A(i_add_term1[8]), .Y(_42_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[8]), .B(_42_), .Y(_43_) );
INVX1 INVX1_12 ( .A(i_add_term2[8]), .Y(_44_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term1[8]), .B(_44_), .Y(_45_) );
INVX1 INVX1_13 ( .A(i_add_term1[9]), .Y(_46_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[9]), .B(_46_), .Y(_47_) );
INVX1 INVX1_14 ( .A(i_add_term2[9]), .Y(_48_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term1[9]), .B(_48_), .Y(_49_) );
OAI22X1 OAI22X1_3 ( .A(_43_), .B(_45_), .C(_47_), .D(_49_), .Y(_50_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_51_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_52_) );
NOR2X1 NOR2X1_20 ( .A(_51_), .B(_52_), .Y(_53_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_54_) );
NAND2X1 NAND2X1_5 ( .A(_53_), .B(_54_), .Y(_55_) );
NOR2X1 NOR2X1_21 ( .A(_50_), .B(_55_), .Y(_9_) );
INVX1 INVX1_15 ( .A(_7_), .Y(_56_) );
NAND2X1 NAND2X1_6 ( .A(1'b0), .B(_9_), .Y(_57_) );
OAI21X1 OAI21X1_3 ( .A(_9_), .B(_56_), .C(_57_), .Y(cskip3_inst_cin) );
INVX1 INVX1_16 ( .A(1'b0), .Y(_61_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_62_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_63_) );
NAND3X1 NAND3X1_1 ( .A(_61_), .B(_63_), .C(_62_), .Y(_64_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_58_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_59_) );
OAI21X1 OAI21X1_4 ( .A(_58_), .B(_59_), .C(1'b0), .Y(_60_) );
NAND2X1 NAND2X1_8 ( .A(_60_), .B(_64_), .Y(_0__0_) );
OAI21X1 OAI21X1_5 ( .A(_61_), .B(_58_), .C(_63_), .Y(_2__1_) );
INVX1 INVX1_17 ( .A(_2__1_), .Y(_68_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_69_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_70_) );
NAND3X1 NAND3X1_2 ( .A(_68_), .B(_70_), .C(_69_), .Y(_71_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_65_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_66_) );
OAI21X1 OAI21X1_6 ( .A(_65_), .B(_66_), .C(_2__1_), .Y(_67_) );
NAND2X1 NAND2X1_10 ( .A(_67_), .B(_71_), .Y(_0__1_) );
OAI21X1 OAI21X1_7 ( .A(_68_), .B(_65_), .C(_70_), .Y(_2__2_) );
INVX1 INVX1_18 ( .A(_2__2_), .Y(_75_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_76_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_77_) );
NAND3X1 NAND3X1_3 ( .A(_75_), .B(_77_), .C(_76_), .Y(_78_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_72_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_73_) );
OAI21X1 OAI21X1_8 ( .A(_72_), .B(_73_), .C(_2__2_), .Y(_74_) );
NAND2X1 NAND2X1_12 ( .A(_74_), .B(_78_), .Y(_0__2_) );
OAI21X1 OAI21X1_9 ( .A(_75_), .B(_72_), .C(_77_), .Y(_2__3_) );
INVX1 INVX1_19 ( .A(_2__3_), .Y(_82_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_83_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_84_) );
NAND3X1 NAND3X1_4 ( .A(_82_), .B(_84_), .C(_83_), .Y(_85_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_79_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_80_) );
OAI21X1 OAI21X1_10 ( .A(_79_), .B(_80_), .C(_2__3_), .Y(_81_) );
NAND2X1 NAND2X1_14 ( .A(_81_), .B(_85_), .Y(_0__3_) );
OAI21X1 OAI21X1_11 ( .A(_82_), .B(_79_), .C(_84_), .Y(_1_) );
INVX1 INVX1_20 ( .A(w_cout_1_), .Y(_89_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_90_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_91_) );
NAND3X1 NAND3X1_5 ( .A(_89_), .B(_91_), .C(_90_), .Y(_92_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_86_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_87_) );
OAI21X1 OAI21X1_12 ( .A(_86_), .B(_87_), .C(w_cout_1_), .Y(_88_) );
NAND2X1 NAND2X1_16 ( .A(_88_), .B(_92_), .Y(_0__4_) );
OAI21X1 OAI21X1_13 ( .A(_89_), .B(_86_), .C(_91_), .Y(_5__1_) );
INVX1 INVX1_21 ( .A(_5__1_), .Y(_96_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_97_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_98_) );
NAND3X1 NAND3X1_6 ( .A(_96_), .B(_98_), .C(_97_), .Y(_99_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_93_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_94_) );
OAI21X1 OAI21X1_14 ( .A(_93_), .B(_94_), .C(_5__1_), .Y(_95_) );
NAND2X1 NAND2X1_18 ( .A(_95_), .B(_99_), .Y(_0__5_) );
OAI21X1 OAI21X1_15 ( .A(_96_), .B(_93_), .C(_98_), .Y(_5__2_) );
INVX1 INVX1_22 ( .A(_5__2_), .Y(_103_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_104_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_105_) );
NAND3X1 NAND3X1_7 ( .A(_103_), .B(_105_), .C(_104_), .Y(_106_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_100_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_101_) );
OAI21X1 OAI21X1_16 ( .A(_100_), .B(_101_), .C(_5__2_), .Y(_102_) );
NAND2X1 NAND2X1_20 ( .A(_102_), .B(_106_), .Y(_0__6_) );
OAI21X1 OAI21X1_17 ( .A(_103_), .B(_100_), .C(_105_), .Y(_5__3_) );
INVX1 INVX1_23 ( .A(_5__3_), .Y(_110_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_111_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_112_) );
NAND3X1 NAND3X1_8 ( .A(_110_), .B(_112_), .C(_111_), .Y(_113_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_107_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_108_) );
OAI21X1 OAI21X1_18 ( .A(_107_), .B(_108_), .C(_5__3_), .Y(_109_) );
NAND2X1 NAND2X1_22 ( .A(_109_), .B(_113_), .Y(_0__7_) );
OAI21X1 OAI21X1_19 ( .A(_110_), .B(_107_), .C(_112_), .Y(_4_) );
INVX1 INVX1_24 ( .A(w_cout_2_), .Y(_117_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_118_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_119_) );
NAND3X1 NAND3X1_9 ( .A(_117_), .B(_119_), .C(_118_), .Y(_120_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_114_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_115_) );
OAI21X1 OAI21X1_20 ( .A(_114_), .B(_115_), .C(w_cout_2_), .Y(_116_) );
NAND2X1 NAND2X1_24 ( .A(_116_), .B(_120_), .Y(_0__8_) );
OAI21X1 OAI21X1_21 ( .A(_117_), .B(_114_), .C(_119_), .Y(_8__1_) );
INVX1 INVX1_25 ( .A(_8__1_), .Y(_124_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_125_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_126_) );
NAND3X1 NAND3X1_10 ( .A(_124_), .B(_126_), .C(_125_), .Y(_127_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_121_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_122_) );
OAI21X1 OAI21X1_22 ( .A(_121_), .B(_122_), .C(_8__1_), .Y(_123_) );
NAND2X1 NAND2X1_26 ( .A(_123_), .B(_127_), .Y(_0__9_) );
OAI21X1 OAI21X1_23 ( .A(_124_), .B(_121_), .C(_126_), .Y(_8__2_) );
INVX1 INVX1_26 ( .A(_8__2_), .Y(_131_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_132_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_133_) );
NAND3X1 NAND3X1_11 ( .A(_131_), .B(_133_), .C(_132_), .Y(_134_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_128_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_129_) );
OAI21X1 OAI21X1_24 ( .A(_128_), .B(_129_), .C(_8__2_), .Y(_130_) );
NAND2X1 NAND2X1_28 ( .A(_130_), .B(_134_), .Y(_0__10_) );
OAI21X1 OAI21X1_25 ( .A(_131_), .B(_128_), .C(_133_), .Y(_8__3_) );
INVX1 INVX1_27 ( .A(_8__3_), .Y(_138_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_139_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_140_) );
NAND3X1 NAND3X1_12 ( .A(_138_), .B(_140_), .C(_139_), .Y(_141_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_135_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_136_) );
OAI21X1 OAI21X1_26 ( .A(_135_), .B(_136_), .C(_8__3_), .Y(_137_) );
NAND2X1 NAND2X1_30 ( .A(_137_), .B(_141_), .Y(_0__11_) );
OAI21X1 OAI21X1_27 ( .A(_138_), .B(_135_), .C(_140_), .Y(_7_) );
INVX1 INVX1_28 ( .A(cskip3_inst_cin), .Y(_145_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_146_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_147_) );
NAND3X1 NAND3X1_13 ( .A(_145_), .B(_147_), .C(_146_), .Y(_148_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_142_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_143_) );
OAI21X1 OAI21X1_28 ( .A(_142_), .B(_143_), .C(cskip3_inst_cin), .Y(_144_) );
NAND2X1 NAND2X1_32 ( .A(_144_), .B(_148_), .Y(_0__12_) );
OAI21X1 OAI21X1_29 ( .A(_145_), .B(_142_), .C(_147_), .Y(cskip3_inst_rca0_w_CARRY_1_) );
INVX1 INVX1_29 ( .A(cskip3_inst_rca0_w_CARRY_1_), .Y(_152_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_153_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_154_) );
NAND3X1 NAND3X1_14 ( .A(_152_), .B(_154_), .C(_153_), .Y(_155_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_149_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_150_) );
OAI21X1 OAI21X1_30 ( .A(_149_), .B(_150_), .C(cskip3_inst_rca0_w_CARRY_1_), .Y(_151_) );
NAND2X1 NAND2X1_34 ( .A(_151_), .B(_155_), .Y(_0__13_) );
OAI21X1 OAI21X1_31 ( .A(_152_), .B(_149_), .C(_154_), .Y(cskip3_inst_rca0_w_CARRY_2_) );
INVX1 INVX1_30 ( .A(cskip3_inst_rca0_w_CARRY_2_), .Y(_159_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_160_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_161_) );
NAND3X1 NAND3X1_15 ( .A(_159_), .B(_161_), .C(_160_), .Y(_162_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_156_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_157_) );
OAI21X1 OAI21X1_32 ( .A(_156_), .B(_157_), .C(cskip3_inst_rca0_w_CARRY_2_), .Y(_158_) );
NAND2X1 NAND2X1_36 ( .A(_158_), .B(_162_), .Y(_0__14_) );
OAI21X1 OAI21X1_33 ( .A(_159_), .B(_156_), .C(_161_), .Y(cskip3_inst_rca0_w_CARRY_3_) );
INVX1 INVX1_31 ( .A(cskip3_inst_rca0_w_CARRY_3_), .Y(_164_) );
NAND2X1 NAND2X1_37 ( .A(1'b0), .B(1'b0), .Y(_165_) );
NOR2X1 NOR2X1_37 ( .A(1'b0), .B(1'b0), .Y(_163_) );
OAI21X1 OAI21X1_34 ( .A(_164_), .B(_163_), .C(_165_), .Y(cskip3_inst_cout0) );
OR2X2 OR2X2_16 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_169_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_170_) );
NAND2X1 NAND2X1_39 ( .A(_170_), .B(_169_), .Y(_166_) );
XNOR2X1 XNOR2X1_1 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_167_) );
XNOR2X1 XNOR2X1_2 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_168_) );
NOR3X1 NOR3X1_1 ( .A(_166_), .B(_167_), .C(_168_), .Y(cskip3_inst_skip0_P) );
INVX1 INVX1_32 ( .A(cskip3_inst_cout0), .Y(_171_) );
NAND2X1 NAND2X1_40 ( .A(1'b0), .B(cskip3_inst_skip0_P), .Y(_172_) );
OAI21X1 OAI21X1_35 ( .A(cskip3_inst_skip0_P), .B(_171_), .C(_172_), .Y(w_cout_4_) );
BUFX2 BUFX2_17 ( .A(1'b0), .Y(_2__0_) );
BUFX2 BUFX2_18 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_19 ( .A(w_cout_1_), .Y(_5__0_) );
BUFX2 BUFX2_20 ( .A(_4_), .Y(_5__4_) );
BUFX2 BUFX2_21 ( .A(w_cout_2_), .Y(_8__0_) );
BUFX2 BUFX2_22 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_23 ( .A(cskip3_inst_cin), .Y(cskip3_inst_rca0_w_CARRY_0_) );
BUFX2 BUFX2_24 ( .A(cskip3_inst_cout0), .Y(cskip3_inst_rca0_w_CARRY_4_) );
BUFX2 BUFX2_25 ( .A(1'b0), .Y(w_cout_0_) );
BUFX2 BUFX2_26 ( .A(cskip3_inst_cin), .Y(w_cout_3_) );
endmodule
