module cla_39bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [38:0] i_add1;
input [38:0] i_add2;
output [39:0] o_result;

NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_408_), .Y(_212__31_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(w_C_32_), .Y(_412_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_413_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_414_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_414_), .C(_413_), .Y(_415_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_409_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_410_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_410_), .C(w_C_32_), .Y(_411_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_415_), .Y(_212__32_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(w_C_33_), .Y(_419_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_420_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_421_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_421_), .C(_420_), .Y(_422_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_416_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_417_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_417_), .C(w_C_33_), .Y(_418_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_422_), .Y(_212__33_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(w_C_34_), .Y(_426_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_427_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_428_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_428_), .C(_427_), .Y(_429_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_423_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_424_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_424_), .C(w_C_34_), .Y(_425_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(_429_), .Y(_212__34_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(w_C_35_), .Y(_433_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_434_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_435_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_435_), .C(_434_), .Y(_436_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_430_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_431_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_431_), .C(w_C_35_), .Y(_432_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_432_), .B(_436_), .Y(_212__35_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(w_C_36_), .Y(_440_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_441_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_442_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_442_), .C(_441_), .Y(_443_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_437_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_438_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_438_), .C(w_C_36_), .Y(_439_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_443_), .Y(_212__36_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(w_C_37_), .Y(_447_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_448_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_449_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_449_), .C(_448_), .Y(_450_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_444_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_445_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_445_), .C(w_C_37_), .Y(_446_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(_450_), .Y(_212__37_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(w_C_38_), .Y(_454_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_455_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_456_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_454_), .B(_456_), .C(_455_), .Y(_457_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_451_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_452_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_452_), .C(w_C_38_), .Y(_453_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(_457_), .Y(_212__38_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_461_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_462_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_463_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_463_), .C(_462_), .Y(_464_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_458_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_459_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_459_), .C(gnd), .Y(_460_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_464_), .Y(_212__0_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_468_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_469_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_470_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_468_), .B(_470_), .C(_469_), .Y(_471_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_465_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_466_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_466_), .C(w_C_1_), .Y(_467_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_467_), .B(_471_), .Y(_212__1_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_475_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_476_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_477_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_477_), .C(_476_), .Y(_478_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_472_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_473_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_473_), .C(w_C_2_), .Y(_474_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_474_), .B(_478_), .Y(_212__2_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_482_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_483_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_484_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_482_), .B(_484_), .C(_483_), .Y(_485_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_479_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_480_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_480_), .C(w_C_3_), .Y(_481_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_485_), .Y(_212__3_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_7_), .Y(w_C_3_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_9_), .C(_7_), .Y(_10_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_8_), .Y(w_C_4_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_12_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_12_), .C(_10_), .Y(_13_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_13_), .Y(w_C_5_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_14_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_14_), .Y(_15_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_16_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_16_), .C(_13_), .Y(_17_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_15_), .Y(w_C_6_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .Y(_18_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add1[6]), .Y(_19_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_20_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_20_), .Y(_21_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_21_), .C(_17_), .Y(_22_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_19_), .C(_22_), .Y(w_C_7_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_23_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_23_), .Y(_24_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_19_), .Y(_25_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(_26_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_27_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(_28_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_28_), .C(_22_), .Y(_29_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_24_), .Y(w_C_8_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_30_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_31_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_32_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_32_), .Y(_33_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_33_), .C(_29_), .Y(_34_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_31_), .Y(_35_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_35_), .Y(w_C_9_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_36_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_36_), .Y(_37_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_38_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_35_), .C(_37_), .Y(w_C_10_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_39_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_39_), .Y(_40_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_38_), .Y(_41_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_37_), .C(_34_), .Y(_42_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_43_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(_44_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_44_), .C(_42_), .Y(_45_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_40_), .Y(_46_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_46_), .Y(w_C_11_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_47_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_47_), .Y(_48_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_49_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_46_), .C(_48_), .Y(w_C_12_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .Y(_50_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add1[12]), .Y(_51_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_49_), .Y(_52_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_48_), .C(_45_), .Y(_53_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_54_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_54_), .Y(_55_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_55_), .C(_53_), .Y(_56_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_51_), .C(_56_), .Y(w_C_13_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_51_), .Y(_57_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_57_), .Y(_58_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_59_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_59_), .Y(_60_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_60_), .C(_56_), .Y(_61_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .C(_61_), .Y(_62_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_62_), .Y(w_C_14_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .Y(_63_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add1[14]), .Y(_64_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_65_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_65_), .Y(_66_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_67_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_67_), .Y(_68_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_68_), .C(_61_), .Y(_69_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_64_), .C(_69_), .Y(w_C_15_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_64_), .Y(_70_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_70_), .Y(_71_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_72_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_72_), .Y(_73_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_73_), .C(_69_), .Y(_74_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .C(_74_), .Y(_75_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_75_), .Y(w_C_16_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .Y(_76_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add1[16]), .Y(_77_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_78_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_78_), .Y(_79_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_80_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_80_), .Y(_81_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_81_), .C(_74_), .Y(_82_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_77_), .C(_82_), .Y(w_C_17_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_77_), .Y(_83_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_83_), .Y(_84_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_85_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_85_), .Y(_86_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_86_), .C(_82_), .Y(_87_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .C(_87_), .Y(_88_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_88_), .Y(w_C_18_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .Y(_89_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add1[18]), .Y(_90_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_91_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_91_), .Y(_92_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_93_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_93_), .Y(_94_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_94_), .C(_87_), .Y(_95_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_90_), .C(_95_), .Y(w_C_19_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_90_), .Y(_96_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_96_), .Y(_97_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_98_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_98_), .Y(_99_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_99_), .C(_95_), .Y(_100_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .C(_100_), .Y(_101_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_101_), .Y(w_C_20_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .Y(_102_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add1[20]), .Y(_103_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_104_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_104_), .Y(_105_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_106_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_106_), .Y(_107_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_107_), .C(_100_), .Y(_108_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_103_), .C(_108_), .Y(w_C_21_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_103_), .Y(_109_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_109_), .Y(_110_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_111_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_111_), .Y(_112_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_112_), .C(_108_), .Y(_113_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .C(_113_), .Y(_114_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_114_), .Y(w_C_22_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .Y(_115_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add1[22]), .Y(_116_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_117_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_117_), .Y(_118_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_119_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_119_), .Y(_120_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_120_), .C(_113_), .Y(_121_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_116_), .C(_121_), .Y(w_C_23_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_116_), .Y(_122_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_122_), .Y(_123_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_124_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_124_), .Y(_125_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_123_), .B(_125_), .C(_121_), .Y(_126_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .C(_126_), .Y(_127_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(_127_), .Y(w_C_24_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .Y(_128_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add1[24]), .Y(_129_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_130_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_130_), .Y(_131_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_132_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_132_), .Y(_133_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_133_), .C(_126_), .Y(_134_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_129_), .C(_134_), .Y(w_C_25_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_129_), .Y(_135_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_135_), .Y(_136_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_137_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_137_), .Y(_138_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_138_), .C(_134_), .Y(_139_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .C(_139_), .Y(_140_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_140_), .Y(w_C_26_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .Y(_141_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add1[26]), .Y(_142_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_143_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_143_), .Y(_144_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_145_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_145_), .Y(_146_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_146_), .C(_139_), .Y(_147_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_142_), .C(_147_), .Y(w_C_27_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_142_), .Y(_148_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_148_), .Y(_149_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_150_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(_150_), .Y(_151_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_151_), .C(_147_), .Y(_152_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .C(_152_), .Y(_153_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_153_), .Y(w_C_28_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .Y(_154_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add1[28]), .Y(_155_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_156_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_157_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_158_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(_158_), .Y(_159_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_159_), .C(_152_), .Y(_160_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_155_), .C(_160_), .Y(w_C_29_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_155_), .Y(_161_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_161_), .Y(_162_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_163_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(_163_), .Y(_164_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_164_), .C(_160_), .Y(_165_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .C(_165_), .Y(_166_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(_166_), .Y(w_C_30_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .Y(_167_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add1[30]), .Y(_168_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_169_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_169_), .Y(_170_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_171_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(_171_), .Y(_172_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_172_), .C(_165_), .Y(_173_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_168_), .C(_173_), .Y(w_C_31_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_174_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(_174_), .Y(_175_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_168_), .Y(_176_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(_176_), .Y(_177_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_178_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_178_), .C(_173_), .Y(_179_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_175_), .Y(w_C_32_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .Y(_180_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add1[32]), .Y(_181_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_181_), .Y(_182_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_175_), .B(_182_), .C(_179_), .Y(_183_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_181_), .C(_183_), .Y(w_C_33_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .Y(_184_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add1[33]), .Y(_185_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_185_), .Y(_186_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_187_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_188_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(_188_), .C(_183_), .Y(_189_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_186_), .Y(w_C_34_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .Y(_190_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add1[34]), .Y(_191_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_191_), .Y(_192_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_192_), .C(_189_), .Y(_193_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_191_), .C(_193_), .Y(w_C_35_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_191_), .Y(_194_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_194_), .Y(_195_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_196_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_196_), .Y(_197_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_197_), .C(_193_), .Y(_198_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .C(_198_), .Y(_199_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_199_), .Y(w_C_36_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_200_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_201_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_199_), .C(_200_), .Y(w_C_37_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_202_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_203_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_203_), .Y(_204_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_201_), .Y(_205_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_205_), .C(_198_), .Y(_206_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_207_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_207_), .C(_206_), .Y(_208_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_202_), .Y(w_C_38_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_209_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_210_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_210_), .C(_208_), .Y(_211_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_211_), .Y(w_C_39_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_212__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_212__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_212__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_212__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_212__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_212__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_212__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_212__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_212__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_212__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_212__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_212__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_212__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_212__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_212__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_212__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_212__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_212__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_212__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_212__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_212__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_212__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_212__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_212__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_212__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_212__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_212__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_212__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_212__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_212__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_212__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_212__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_212__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_212__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_212__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_212__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_212__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_212__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_212__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(w_C_39_), .Y(o_result[39]) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_216_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_217_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_218_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_218_), .C(_217_), .Y(_219_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_213_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_214_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_214_), .C(w_C_4_), .Y(_215_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_219_), .Y(_212__4_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_223_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_224_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_225_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_225_), .C(_224_), .Y(_226_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_220_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_221_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_221_), .C(w_C_5_), .Y(_222_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_226_), .Y(_212__5_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_230_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_231_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_232_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_232_), .C(_231_), .Y(_233_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_227_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_228_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_228_), .C(w_C_6_), .Y(_229_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_233_), .Y(_212__6_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_237_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_238_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_239_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_239_), .C(_238_), .Y(_240_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_234_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_235_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_235_), .C(w_C_7_), .Y(_236_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_240_), .Y(_212__7_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_244_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_245_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_246_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_246_), .C(_245_), .Y(_247_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_241_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_242_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_242_), .C(w_C_8_), .Y(_243_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_247_), .Y(_212__8_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_251_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_252_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_253_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_253_), .C(_252_), .Y(_254_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_248_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_249_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_249_), .C(w_C_9_), .Y(_250_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_254_), .Y(_212__9_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_258_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_259_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_260_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_260_), .C(_259_), .Y(_261_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_255_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_256_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_256_), .C(w_C_10_), .Y(_257_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_261_), .Y(_212__10_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_265_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_266_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_267_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_267_), .C(_266_), .Y(_268_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_262_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_263_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_263_), .C(w_C_11_), .Y(_264_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_268_), .Y(_212__11_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(w_C_12_), .Y(_272_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_273_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_274_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_274_), .C(_273_), .Y(_275_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_269_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_270_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_270_), .C(w_C_12_), .Y(_271_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_275_), .Y(_212__12_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(w_C_13_), .Y(_279_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_280_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_281_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_279_), .B(_281_), .C(_280_), .Y(_282_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_276_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_277_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_277_), .C(w_C_13_), .Y(_278_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_282_), .Y(_212__13_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(w_C_14_), .Y(_286_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_287_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_288_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_288_), .C(_287_), .Y(_289_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_283_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_284_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_283_), .B(_284_), .C(w_C_14_), .Y(_285_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_289_), .Y(_212__14_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(_293_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_294_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_295_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_295_), .C(_294_), .Y(_296_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_290_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_291_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_291_), .C(w_C_15_), .Y(_292_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_292_), .B(_296_), .Y(_212__15_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(w_C_16_), .Y(_300_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_301_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_302_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_302_), .C(_301_), .Y(_303_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_297_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_298_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_298_), .C(w_C_16_), .Y(_299_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_303_), .Y(_212__16_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(w_C_17_), .Y(_307_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_308_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_309_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_309_), .C(_308_), .Y(_310_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_304_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_305_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_305_), .C(w_C_17_), .Y(_306_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_310_), .Y(_212__17_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(w_C_18_), .Y(_314_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_315_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_316_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_316_), .C(_315_), .Y(_317_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_311_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_312_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_312_), .C(w_C_18_), .Y(_313_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_317_), .Y(_212__18_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(w_C_19_), .Y(_321_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_322_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_323_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_323_), .C(_322_), .Y(_324_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_318_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_319_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_319_), .C(w_C_19_), .Y(_320_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_324_), .Y(_212__19_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(w_C_20_), .Y(_328_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_329_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_330_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_330_), .C(_329_), .Y(_331_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_325_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_326_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_326_), .C(w_C_20_), .Y(_327_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_331_), .Y(_212__20_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(w_C_21_), .Y(_335_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_336_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_337_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_335_), .B(_337_), .C(_336_), .Y(_338_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_332_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_333_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_333_), .C(w_C_21_), .Y(_334_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_338_), .Y(_212__21_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(w_C_22_), .Y(_342_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_343_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_344_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_344_), .C(_343_), .Y(_345_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_339_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_340_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_340_), .C(w_C_22_), .Y(_341_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_345_), .Y(_212__22_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(w_C_23_), .Y(_349_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_350_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_351_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_351_), .C(_350_), .Y(_352_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_346_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_347_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_347_), .C(w_C_23_), .Y(_348_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_352_), .Y(_212__23_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(w_C_24_), .Y(_356_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_357_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_358_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_358_), .C(_357_), .Y(_359_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_353_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_354_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_354_), .C(w_C_24_), .Y(_355_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_359_), .Y(_212__24_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(w_C_25_), .Y(_363_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_364_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_365_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_365_), .C(_364_), .Y(_366_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_360_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_361_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_361_), .C(w_C_25_), .Y(_362_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_366_), .Y(_212__25_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(w_C_26_), .Y(_370_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_371_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_372_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_372_), .C(_371_), .Y(_373_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_367_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_368_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_368_), .C(w_C_26_), .Y(_369_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_373_), .Y(_212__26_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(w_C_27_), .Y(_377_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_378_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_379_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_379_), .C(_378_), .Y(_380_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_374_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_375_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_375_), .C(w_C_27_), .Y(_376_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_380_), .Y(_212__27_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(w_C_28_), .Y(_384_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_385_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_386_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_386_), .C(_385_), .Y(_387_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_381_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_382_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_382_), .C(w_C_28_), .Y(_383_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_387_), .Y(_212__28_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(w_C_29_), .Y(_391_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_392_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_393_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_393_), .C(_392_), .Y(_394_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_388_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_389_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(_389_), .C(w_C_29_), .Y(_390_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_394_), .Y(_212__29_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(w_C_30_), .Y(_398_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_399_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_400_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_400_), .C(_399_), .Y(_401_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_395_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_396_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_396_), .C(w_C_30_), .Y(_397_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_401_), .Y(_212__30_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(w_C_31_), .Y(_405_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_406_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_407_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_407_), .C(_406_), .Y(_408_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_402_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_403_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_403_), .C(w_C_31_), .Y(_404_) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(w_C_39_), .Y(_212__39_) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
