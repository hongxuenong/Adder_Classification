module csa_38bit ( gnd, vdd, i_add_term1, i_add_term2, sum, cout);

input gnd, vdd;
output cout;
input [37:0] i_add_term1;
input [37:0] i_add_term2;
output [37:0] sum;

OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_296_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_297_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_297_), .C(_296_), .Y(_298_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_292_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_293_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_292_), .B(_293_), .C(_24__3_), .Y(_294_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_298_), .Y(_22__3_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_292_), .C(_297_), .Y(_20_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_24__1_), .Y(_302_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_303_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_304_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_304_), .C(_303_), .Y(_305_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_299_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_300_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_300_), .C(_24__1_), .Y(_301_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_305_), .Y(_22__1_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_299_), .C(_304_), .Y(_24__2_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_24__2_), .Y(_309_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_310_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_311_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_311_), .C(_310_), .Y(_312_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_306_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_307_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_307_), .C(_24__2_), .Y(_308_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_312_), .Y(_22__2_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_309_), .B(_306_), .C(_311_), .Y(_24__3_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(_313_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(w_cout_4_), .Y(_314_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_313_), .C(_314_), .Y(w_cout_5_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_27__0_), .Y(_315_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_28__0_), .B(w_cout_4_), .Y(_316_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_315_), .C(_316_), .Y(_0__20_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_27__1_), .Y(_317_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_28__1_), .Y(_318_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_317_), .C(_318_), .Y(_0__21_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_27__2_), .Y(_319_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_28__2_), .Y(_320_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_319_), .C(_320_), .Y(_0__22_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_27__3_), .Y(_321_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_28__3_), .Y(_322_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_321_), .C(_322_), .Y(_0__23_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_326_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_327_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_328_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_328_), .C(_327_), .Y(_329_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_323_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_324_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_324_), .C(gnd), .Y(_325_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_329_), .Y(_27__0_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_323_), .C(_328_), .Y(_29__1_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_29__3_), .Y(_333_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_334_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_335_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_335_), .C(_334_), .Y(_336_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_330_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_331_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_331_), .C(_29__3_), .Y(_332_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_336_), .Y(_27__3_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_330_), .C(_335_), .Y(_25_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_29__1_), .Y(_340_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_341_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_342_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_342_), .C(_341_), .Y(_343_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_337_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_338_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_338_), .C(_29__1_), .Y(_339_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_343_), .Y(_27__1_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_337_), .C(_342_), .Y(_29__2_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_29__2_), .Y(_347_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_348_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_349_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_349_), .C(_348_), .Y(_350_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_344_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_345_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_345_), .C(_29__2_), .Y(_346_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_350_), .Y(_27__2_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_344_), .C(_349_), .Y(_29__3_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_354_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_355_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_356_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_356_), .C(_355_), .Y(_357_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_351_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_352_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_352_), .C(vdd), .Y(_353_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_357_), .Y(_28__0_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_351_), .C(_356_), .Y(_30__1_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_30__3_), .Y(_361_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_362_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_363_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_363_), .C(_362_), .Y(_364_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_358_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_359_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_358_), .B(_359_), .C(_30__3_), .Y(_360_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_364_), .Y(_28__3_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_358_), .C(_363_), .Y(_26_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_30__1_), .Y(_368_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_369_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_370_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_370_), .C(_369_), .Y(_371_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_365_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_366_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_365_), .B(_366_), .C(_30__1_), .Y(_367_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_371_), .Y(_28__1_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_365_), .C(_370_), .Y(_30__2_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_30__2_), .Y(_375_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_376_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_377_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_377_), .C(_376_), .Y(_378_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_372_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_373_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_373_), .C(_30__2_), .Y(_374_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_378_), .Y(_28__2_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_372_), .C(_377_), .Y(_30__3_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_31_), .Y(_379_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(w_cout_5_), .Y(_380_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_379_), .C(_380_), .Y(w_cout_6_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_33__0_), .Y(_381_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_34__0_), .B(w_cout_5_), .Y(_382_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_381_), .C(_382_), .Y(_0__24_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_33__1_), .Y(_383_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_34__1_), .Y(_384_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_383_), .C(_384_), .Y(_0__25_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_33__2_), .Y(_385_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_34__2_), .Y(_386_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_385_), .C(_386_), .Y(_0__26_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_33__3_), .Y(_387_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_34__3_), .Y(_388_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_387_), .C(_388_), .Y(_0__27_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_392_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_393_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_394_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_392_), .B(_394_), .C(_393_), .Y(_395_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_389_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_390_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_390_), .C(gnd), .Y(_391_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_395_), .Y(_33__0_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_392_), .B(_389_), .C(_394_), .Y(_35__1_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_35__3_), .Y(_399_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_400_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_401_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_401_), .C(_400_), .Y(_402_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_396_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_397_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_397_), .C(_35__3_), .Y(_398_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_402_), .Y(_33__3_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_396_), .C(_401_), .Y(_31_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_35__1_), .Y(_406_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_407_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_408_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_406_), .B(_408_), .C(_407_), .Y(_409_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_403_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_404_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_404_), .C(_35__1_), .Y(_405_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_409_), .Y(_33__1_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_406_), .B(_403_), .C(_408_), .Y(_35__2_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_35__2_), .Y(_413_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_414_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_415_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_415_), .C(_414_), .Y(_416_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_410_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_411_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(_411_), .C(_35__2_), .Y(_412_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_416_), .Y(_33__2_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_410_), .C(_415_), .Y(_35__3_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_420_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_421_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_422_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_420_), .B(_422_), .C(_421_), .Y(_423_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_417_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_418_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_418_), .C(vdd), .Y(_419_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_423_), .Y(_34__0_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_420_), .B(_417_), .C(_422_), .Y(_36__1_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_36__3_), .Y(_427_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_428_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_429_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_427_), .B(_429_), .C(_428_), .Y(_430_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_424_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_425_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_425_), .C(_36__3_), .Y(_426_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_430_), .Y(_34__3_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_427_), .B(_424_), .C(_429_), .Y(_32_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_36__1_), .Y(_434_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_435_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_436_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_436_), .C(_435_), .Y(_437_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_431_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_432_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_432_), .C(_36__1_), .Y(_433_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_437_), .Y(_34__1_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_431_), .C(_436_), .Y(_36__2_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_36__2_), .Y(_441_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_442_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_443_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_443_), .C(_442_), .Y(_444_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_438_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_439_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_439_), .C(_36__2_), .Y(_440_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_444_), .Y(_34__2_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_438_), .C(_443_), .Y(_36__3_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_37_), .Y(_445_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(w_cout_6_), .Y(_446_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_445_), .C(_446_), .Y(w_cout_7_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_39__0_), .Y(_447_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_40__0_), .B(w_cout_6_), .Y(_448_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_447_), .C(_448_), .Y(_0__28_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_39__1_), .Y(_449_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_40__1_), .Y(_450_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_449_), .C(_450_), .Y(_0__29_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_39__2_), .Y(_451_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_40__2_), .Y(_452_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_451_), .C(_452_), .Y(_0__30_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_39__3_), .Y(_453_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_40__3_), .Y(_454_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_453_), .C(_454_), .Y(_0__31_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_458_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_459_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_460_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_460_), .C(_459_), .Y(_461_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_455_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_456_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_456_), .C(gnd), .Y(_457_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_461_), .Y(_39__0_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_455_), .C(_460_), .Y(_41__1_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_41__3_), .Y(_465_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_466_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_467_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_467_), .C(_466_), .Y(_468_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_462_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_463_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_462_), .B(_463_), .C(_41__3_), .Y(_464_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_468_), .Y(_39__3_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_462_), .C(_467_), .Y(_37_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_41__1_), .Y(_472_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_473_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_474_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_474_), .C(_473_), .Y(_475_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_469_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_470_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_470_), .C(_41__1_), .Y(_471_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_475_), .Y(_39__1_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_469_), .C(_474_), .Y(_41__2_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_41__2_), .Y(_479_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_480_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_481_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_481_), .C(_480_), .Y(_482_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_476_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_477_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_477_), .C(_41__2_), .Y(_478_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_482_), .Y(_39__2_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_476_), .C(_481_), .Y(_41__3_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_486_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_487_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_488_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_488_), .C(_487_), .Y(_489_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_483_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_484_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_483_), .B(_484_), .C(vdd), .Y(_485_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_489_), .Y(_40__0_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_483_), .C(_488_), .Y(_42__1_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_42__3_), .Y(_493_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_494_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_495_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_495_), .C(_494_), .Y(_496_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_490_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_491_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_490_), .B(_491_), .C(_42__3_), .Y(_492_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_492_), .B(_496_), .Y(_40__3_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_490_), .C(_495_), .Y(_38_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_42__1_), .Y(_500_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_501_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_502_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_502_), .C(_501_), .Y(_503_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_497_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_498_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_497_), .B(_498_), .C(_42__1_), .Y(_499_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_503_), .Y(_40__1_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_497_), .C(_502_), .Y(_42__2_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_42__2_), .Y(_507_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_508_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_509_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_509_), .C(_508_), .Y(_510_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_504_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_505_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_504_), .B(_505_), .C(_42__2_), .Y(_506_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_510_), .Y(_40__2_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_504_), .C(_509_), .Y(_42__3_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(_511_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(w_cout_7_), .Y(_512_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_511_), .C(_512_), .Y(csa_inst_cin) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_45__0_), .Y(_513_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_46__0_), .B(w_cout_7_), .Y(_514_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_513_), .C(_514_), .Y(_0__32_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_45__1_), .Y(_515_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_46__1_), .Y(_516_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_515_), .C(_516_), .Y(_0__33_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_45__2_), .Y(_517_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_46__2_), .Y(_518_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_517_), .C(_518_), .Y(_0__34_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_45__3_), .Y(_519_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_46__3_), .Y(_520_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_519_), .C(_520_), .Y(_0__35_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_524_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_525_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_526_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_526_), .C(_525_), .Y(_527_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_521_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_522_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_522_), .C(gnd), .Y(_523_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_527_), .Y(_45__0_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_521_), .C(_526_), .Y(_47__1_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_47__3_), .Y(_531_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_532_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_533_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_533_), .C(_532_), .Y(_534_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_528_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_529_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_529_), .C(_47__3_), .Y(_530_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_534_), .Y(_45__3_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_528_), .C(_533_), .Y(_43_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_47__1_), .Y(_538_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_539_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_540_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_540_), .C(_539_), .Y(_541_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_535_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_536_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_536_), .C(_47__1_), .Y(_537_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_541_), .Y(_45__1_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_535_), .C(_540_), .Y(_47__2_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_47__2_), .Y(_545_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_546_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_547_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_547_), .C(_546_), .Y(_548_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_542_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_543_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_542_), .B(_543_), .C(_47__2_), .Y(_544_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_548_), .Y(_45__2_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_542_), .C(_547_), .Y(_47__3_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_552_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_553_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_554_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_552_), .B(_554_), .C(_553_), .Y(_555_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_549_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_550_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(_550_), .C(vdd), .Y(_551_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_551_), .B(_555_), .Y(_46__0_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_552_), .B(_549_), .C(_554_), .Y(_48__1_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_48__3_), .Y(_559_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_560_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_561_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_561_), .C(_560_), .Y(_562_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_556_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_557_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_556_), .B(_557_), .C(_48__3_), .Y(_558_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_562_), .Y(_46__3_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_556_), .C(_561_), .Y(_44_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_48__1_), .Y(_566_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_567_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_568_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_568_), .C(_567_), .Y(_569_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_563_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_564_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(_564_), .C(_48__1_), .Y(_565_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_569_), .Y(_46__1_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_563_), .C(_568_), .Y(_48__2_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_48__2_), .Y(_573_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_574_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_575_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_575_), .C(_574_), .Y(_576_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_570_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_571_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_571_), .C(_48__2_), .Y(_572_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_576_), .Y(_46__2_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_570_), .C(_575_), .Y(_48__3_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cout0_0), .Y(_577_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cout0_1), .B(csa_inst_cin), .Y(_578_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .B(_577_), .C(_578_), .Y(w_cout_9_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_0_fa0_o_sum), .Y(_581_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_1_fa0_o_sum), .B(csa_inst_cin), .Y(_582_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .B(_581_), .C(_582_), .Y(_0__36_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_0_fa31_o_sum), .Y(_579_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .B(csa_inst_rca0_1_fa31_o_sum), .Y(_580_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .B(_579_), .C(_580_), .Y(_0__37_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_586_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_587_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_588_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_586_), .B(_588_), .C(_587_), .Y(_589_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_583_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_584_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_583_), .B(_584_), .C(gnd), .Y(_585_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_585_), .B(_589_), .Y(csa_inst_rca0_0_fa0_o_sum) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_586_), .B(_583_), .C(_588_), .Y(csa_inst_rca0_0_c) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_0_c), .Y(_593_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_594_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_595_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_595_), .C(_594_), .Y(_596_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_590_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_591_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_590_), .B(_591_), .C(csa_inst_rca0_0_c), .Y(_592_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_592_), .B(_596_), .Y(csa_inst_rca0_0_fa31_o_sum) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_590_), .C(_595_), .Y(csa_inst_cout0_0) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_600_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_601_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_602_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_602_), .C(_601_), .Y(_603_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_597_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_598_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_597_), .B(_598_), .C(vdd), .Y(_599_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_599_), .B(_603_), .Y(csa_inst_rca0_1_fa0_o_sum) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_597_), .C(_602_), .Y(csa_inst_rca0_1_c) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_1_c), .Y(_607_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_608_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_609_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_609_), .C(_608_), .Y(_610_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_604_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_605_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_604_), .B(_605_), .C(csa_inst_rca0_1_c), .Y(_606_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_610_), .Y(csa_inst_rca0_1_fa31_o_sum) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_604_), .C(_609_), .Y(csa_inst_cout0_1) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_614_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_615_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_616_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_616_), .C(_615_), .Y(_617_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_611_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_612_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_612_), .C(gnd), .Y(_613_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_613_), .B(_617_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_611_), .C(_616_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_i_carry), .Y(_621_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_622_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_623_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_623_), .C(_622_), .Y(_624_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_618_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_619_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_618_), .B(_619_), .C(rca_inst_fa3_i_carry), .Y(_620_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_624_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_618_), .C(_623_), .Y(rca_inst_cout) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_carry), .Y(_628_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_629_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_630_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_630_), .C(_629_), .Y(_631_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_625_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_626_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_625_), .B(_626_), .C(rca_inst_fa0_o_carry), .Y(_627_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(_631_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_625_), .C(_630_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_carry), .Y(_635_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_636_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_637_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_637_), .C(_636_), .Y(_638_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_632_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_633_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_632_), .B(_633_), .C(rca_inst_fa_1__o_carry), .Y(_634_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_634_), .B(_638_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_632_), .C(_637_), .Y(rca_inst_fa3_i_carry) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .Y(cout) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_0__37_), .Y(sum[37]) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_49_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(rca_inst_cout), .Y(_50_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_49_), .C(_50_), .Y(w_cout_1_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_3__0_), .Y(_51_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_4__0_), .B(rca_inst_cout), .Y(_52_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_51_), .C(_52_), .Y(_0__4_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_3__1_), .Y(_53_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_4__1_), .Y(_54_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_53_), .C(_54_), .Y(_0__5_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_3__2_), .Y(_55_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_4__2_), .Y(_56_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_55_), .C(_56_), .Y(_0__6_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_3__3_), .Y(_57_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_4__3_), .Y(_58_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_57_), .C(_58_), .Y(_0__7_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_62_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_63_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_64_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_64_), .C(_63_), .Y(_65_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_59_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_60_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_60_), .C(gnd), .Y(_61_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_65_), .Y(_3__0_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_59_), .C(_64_), .Y(_5__1_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_5__3_), .Y(_69_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_70_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_71_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_71_), .C(_70_), .Y(_72_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_66_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_67_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_67_), .C(_5__3_), .Y(_68_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_72_), .Y(_3__3_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_66_), .C(_71_), .Y(_1_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(_5__1_), .Y(_76_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_77_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_78_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_78_), .C(_77_), .Y(_79_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_73_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_74_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_74_), .C(_5__1_), .Y(_75_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_79_), .Y(_3__1_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_73_), .C(_78_), .Y(_5__2_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_5__2_), .Y(_83_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_84_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_85_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_85_), .C(_84_), .Y(_86_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_80_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_81_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_81_), .C(_5__2_), .Y(_82_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_86_), .Y(_3__2_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_80_), .C(_85_), .Y(_5__3_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_90_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_91_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_92_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_92_), .C(_91_), .Y(_93_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_87_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_88_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_88_), .C(vdd), .Y(_89_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_93_), .Y(_4__0_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_87_), .C(_92_), .Y(_6__1_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_6__3_), .Y(_97_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_98_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_99_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_99_), .C(_98_), .Y(_100_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_94_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_95_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_95_), .C(_6__3_), .Y(_96_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_100_), .Y(_4__3_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_94_), .C(_99_), .Y(_2_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_6__1_), .Y(_104_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_105_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_106_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_106_), .C(_105_), .Y(_107_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_101_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_102_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_102_), .C(_6__1_), .Y(_103_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_107_), .Y(_4__1_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_101_), .C(_106_), .Y(_6__2_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_6__2_), .Y(_111_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_112_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_113_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_113_), .C(_112_), .Y(_114_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_108_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_109_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_109_), .C(_6__2_), .Y(_110_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_114_), .Y(_4__2_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_108_), .C(_113_), .Y(_6__3_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_115_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(w_cout_1_), .Y(_116_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_115_), .C(_116_), .Y(w_cout_2_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_9__0_), .Y(_117_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_10__0_), .B(w_cout_1_), .Y(_118_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_117_), .C(_118_), .Y(_0__8_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_9__1_), .Y(_119_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_10__1_), .Y(_120_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_119_), .C(_120_), .Y(_0__9_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_9__2_), .Y(_121_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_10__2_), .Y(_122_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_121_), .C(_122_), .Y(_0__10_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_9__3_), .Y(_123_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_10__3_), .Y(_124_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_123_), .C(_124_), .Y(_0__11_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_128_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_129_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_130_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_130_), .C(_129_), .Y(_131_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_125_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_126_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_126_), .C(gnd), .Y(_127_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_131_), .Y(_9__0_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_125_), .C(_130_), .Y(_11__1_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_11__3_), .Y(_135_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_136_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_137_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_137_), .C(_136_), .Y(_138_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_132_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_133_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_133_), .C(_11__3_), .Y(_134_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_138_), .Y(_9__3_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_132_), .C(_137_), .Y(_7_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_11__1_), .Y(_142_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_143_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_144_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_144_), .C(_143_), .Y(_145_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_139_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_140_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_140_), .C(_11__1_), .Y(_141_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_145_), .Y(_9__1_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_139_), .C(_144_), .Y(_11__2_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(_11__2_), .Y(_149_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_150_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_151_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_151_), .C(_150_), .Y(_152_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_146_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_147_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_147_), .C(_11__2_), .Y(_148_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_152_), .Y(_9__2_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_146_), .C(_151_), .Y(_11__3_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_156_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_157_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_158_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_158_), .C(_157_), .Y(_159_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_153_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_154_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_154_), .C(vdd), .Y(_155_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_159_), .Y(_10__0_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_153_), .C(_158_), .Y(_12__1_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(_12__3_), .Y(_163_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_164_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_165_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_165_), .C(_164_), .Y(_166_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_160_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_161_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_161_), .C(_12__3_), .Y(_162_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_166_), .Y(_10__3_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_160_), .C(_165_), .Y(_8_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_12__1_), .Y(_170_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_171_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_172_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_172_), .C(_171_), .Y(_173_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_167_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_168_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_168_), .C(_12__1_), .Y(_169_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_173_), .Y(_10__1_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_167_), .C(_172_), .Y(_12__2_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(_12__2_), .Y(_177_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_178_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_179_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_179_), .C(_178_), .Y(_180_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_174_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_175_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_175_), .C(_12__2_), .Y(_176_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_180_), .Y(_10__2_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_174_), .C(_179_), .Y(_12__3_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_181_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(w_cout_2_), .Y(_182_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_181_), .C(_182_), .Y(w_cout_3_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(_15__0_), .Y(_183_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_16__0_), .B(w_cout_2_), .Y(_184_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_183_), .C(_184_), .Y(_0__12_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_15__1_), .Y(_185_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_16__1_), .Y(_186_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_185_), .C(_186_), .Y(_0__13_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_15__2_), .Y(_187_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_16__2_), .Y(_188_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_187_), .C(_188_), .Y(_0__14_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(_15__3_), .Y(_189_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_16__3_), .Y(_190_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_189_), .C(_190_), .Y(_0__15_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_194_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_195_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_196_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_196_), .C(_195_), .Y(_197_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_191_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_192_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_192_), .C(gnd), .Y(_193_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_197_), .Y(_15__0_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_191_), .C(_196_), .Y(_17__1_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(_17__3_), .Y(_201_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_202_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_203_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_203_), .C(_202_), .Y(_204_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_198_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_199_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_199_), .C(_17__3_), .Y(_200_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_204_), .Y(_15__3_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_198_), .C(_203_), .Y(_13_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(_17__1_), .Y(_208_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_209_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_210_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_210_), .C(_209_), .Y(_211_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_205_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_206_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_206_), .C(_17__1_), .Y(_207_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_211_), .Y(_15__1_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_205_), .C(_210_), .Y(_17__2_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(_17__2_), .Y(_215_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_216_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_217_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_217_), .C(_216_), .Y(_218_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_212_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_213_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_213_), .C(_17__2_), .Y(_214_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_218_), .Y(_15__2_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_212_), .C(_217_), .Y(_17__3_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_222_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_223_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_224_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_224_), .C(_223_), .Y(_225_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_219_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_220_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_220_), .C(vdd), .Y(_221_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_225_), .Y(_16__0_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_219_), .C(_224_), .Y(_18__1_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(_18__3_), .Y(_229_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_230_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_231_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_231_), .C(_230_), .Y(_232_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_226_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_227_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_227_), .C(_18__3_), .Y(_228_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_232_), .Y(_16__3_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_226_), .C(_231_), .Y(_14_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_18__1_), .Y(_236_) );
OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_237_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_238_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_238_), .C(_237_), .Y(_239_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_233_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_234_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_234_), .C(_18__1_), .Y(_235_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_239_), .Y(_16__1_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_233_), .C(_238_), .Y(_18__2_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(_18__2_), .Y(_243_) );
OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_244_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_245_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_245_), .C(_244_), .Y(_246_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_240_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_241_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_241_), .C(_18__2_), .Y(_242_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_246_), .Y(_16__2_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_240_), .C(_245_), .Y(_18__3_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_247_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(w_cout_3_), .Y(_248_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_247_), .C(_248_), .Y(w_cout_4_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_21__0_), .Y(_249_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_22__0_), .B(w_cout_3_), .Y(_250_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_249_), .C(_250_), .Y(_0__16_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_21__1_), .Y(_251_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_22__1_), .Y(_252_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_251_), .C(_252_), .Y(_0__17_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_21__2_), .Y(_253_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_22__2_), .Y(_254_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_253_), .C(_254_), .Y(_0__18_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_21__3_), .Y(_255_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_22__3_), .Y(_256_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_255_), .C(_256_), .Y(_0__19_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_260_) );
OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_261_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_262_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_262_), .C(_261_), .Y(_263_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_257_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_258_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_258_), .C(gnd), .Y(_259_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_263_), .Y(_21__0_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_257_), .C(_262_), .Y(_23__1_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_23__3_), .Y(_267_) );
OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_268_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_269_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_269_), .C(_268_), .Y(_270_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_264_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_265_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_265_), .C(_23__3_), .Y(_266_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_270_), .Y(_21__3_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_264_), .C(_269_), .Y(_19_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(_23__1_), .Y(_274_) );
OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_275_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_276_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_276_), .C(_275_), .Y(_277_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_271_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_272_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_272_), .C(_23__1_), .Y(_273_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_277_), .Y(_21__1_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_271_), .C(_276_), .Y(_23__2_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(_23__2_), .Y(_281_) );
OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_282_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_283_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_283_), .C(_282_), .Y(_284_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_278_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_279_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_279_), .C(_23__2_), .Y(_280_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_284_), .Y(_21__2_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_278_), .C(_283_), .Y(_23__3_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_288_) );
OR2X2 OR2X2_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_289_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_290_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_290_), .C(_289_), .Y(_291_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_285_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_286_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_286_), .C(vdd), .Y(_287_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_287_), .B(_291_), .Y(_22__0_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_285_), .C(_290_), .Y(_24__1_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(_24__3_), .Y(_295_) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .Y(w_cout_0_) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .Y(w_cout_8_) );
endmodule
