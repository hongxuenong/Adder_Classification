module carry_lookahead_adder_7bit (i_add1, i_add2, o_result);

input [6:0] i_add1;
input [6:0] i_add2;
output [7:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX2 BUFX2_1 ( .A(_21__1_), .Y(o_result[1]) );
BUFX2 BUFX2_2 ( .A(_21__2_), .Y(o_result[2]) );
BUFX2 BUFX2_3 ( .A(_21__3_), .Y(o_result[3]) );
BUFX2 BUFX2_4 ( .A(_21__4_), .Y(o_result[4]) );
BUFX2 BUFX2_5 ( .A(_21__5_), .Y(o_result[5]) );
BUFX2 BUFX2_6 ( .A(_21__6_), .Y(o_result[6]) );
BUFX2 BUFX2_7 ( .A(w_C_7_), .Y(o_result[7]) );
INVX1 INVX1_1 ( .A(w_C_4_), .Y(_25_) );
OR2X2 OR2X2_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_26_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_27_) );
NAND3X1 NAND3X1_1 ( .A(_25_), .B(_27_), .C(_26_), .Y(_28_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_22_) );
AND2X2 AND2X2_1 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_23_) );
OAI21X1 OAI21X1_1 ( .A(_22_), .B(_23_), .C(w_C_4_), .Y(_24_) );
NAND2X1 NAND2X1_2 ( .A(_24_), .B(_28_), .Y(_21__4_) );
INVX1 INVX1_2 ( .A(w_C_5_), .Y(_32_) );
OR2X2 OR2X2_2 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_33_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_34_) );
NAND3X1 NAND3X1_2 ( .A(_32_), .B(_34_), .C(_33_), .Y(_35_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_29_) );
AND2X2 AND2X2_2 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_30_) );
OAI21X1 OAI21X1_2 ( .A(_29_), .B(_30_), .C(w_C_5_), .Y(_31_) );
NAND2X1 NAND2X1_4 ( .A(_31_), .B(_35_), .Y(_21__5_) );
INVX1 INVX1_3 ( .A(w_C_6_), .Y(_39_) );
OR2X2 OR2X2_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_40_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_41_) );
NAND3X1 NAND3X1_3 ( .A(_39_), .B(_41_), .C(_40_), .Y(_42_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_36_) );
AND2X2 AND2X2_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_37_) );
OAI21X1 OAI21X1_3 ( .A(_36_), .B(_37_), .C(w_C_6_), .Y(_38_) );
NAND2X1 NAND2X1_6 ( .A(_38_), .B(_42_), .Y(_21__6_) );
INVX1 INVX1_4 ( .A(gnd), .Y(_46_) );
OR2X2 OR2X2_4 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_47_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_48_) );
NAND3X1 NAND3X1_4 ( .A(_46_), .B(_48_), .C(_47_), .Y(_49_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_43_) );
AND2X2 AND2X2_4 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_44_) );
OAI21X1 OAI21X1_4 ( .A(_43_), .B(_44_), .C(gnd), .Y(_45_) );
NAND2X1 NAND2X1_8 ( .A(_45_), .B(_49_), .Y(_21__0_) );
INVX1 INVX1_5 ( .A(w_C_1_), .Y(_53_) );
OR2X2 OR2X2_5 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_54_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_55_) );
NAND3X1 NAND3X1_5 ( .A(_53_), .B(_55_), .C(_54_), .Y(_56_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_50_) );
AND2X2 AND2X2_5 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_51_) );
OAI21X1 OAI21X1_5 ( .A(_50_), .B(_51_), .C(w_C_1_), .Y(_52_) );
NAND2X1 NAND2X1_10 ( .A(_52_), .B(_56_), .Y(_21__1_) );
INVX1 INVX1_6 ( .A(w_C_2_), .Y(_60_) );
OR2X2 OR2X2_6 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_61_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_62_) );
NAND3X1 NAND3X1_6 ( .A(_60_), .B(_62_), .C(_61_), .Y(_63_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_57_) );
AND2X2 AND2X2_6 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_58_) );
OAI21X1 OAI21X1_6 ( .A(_57_), .B(_58_), .C(w_C_2_), .Y(_59_) );
NAND2X1 NAND2X1_12 ( .A(_59_), .B(_63_), .Y(_21__2_) );
INVX1 INVX1_7 ( .A(w_C_3_), .Y(_67_) );
OR2X2 OR2X2_7 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_68_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_69_) );
NAND3X1 NAND3X1_7 ( .A(_67_), .B(_69_), .C(_68_), .Y(_70_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_64_) );
AND2X2 AND2X2_7 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_65_) );
OAI21X1 OAI21X1_7 ( .A(_64_), .B(_65_), .C(w_C_3_), .Y(_66_) );
NAND2X1 NAND2X1_14 ( .A(_66_), .B(_70_), .Y(_21__3_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_8 ( .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_17 ( .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_8 ( .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_9 ( .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_8 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_9 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_8 ( .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_19 ( .A(_4_), .B(_7_), .Y(w_C_3_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
NAND3X1 NAND3X1_9 ( .A(_4_), .B(_8_), .C(_7_), .Y(_9_) );
OAI21X1 OAI21X1_9 ( .A(i_add2[3]), .B(i_add1[3]), .C(_9_), .Y(_10_) );
INVX1 INVX1_10 ( .A(_10_), .Y(w_C_4_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
OR2X2 OR2X2_10 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_12_) );
OR2X2 OR2X2_11 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
NAND3X1 NAND3X1_10 ( .A(_12_), .B(_13_), .C(_9_), .Y(_14_) );
NAND2X1 NAND2X1_22 ( .A(_11_), .B(_14_), .Y(w_C_5_) );
OR2X2 OR2X2_12 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_15_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_16_) );
NAND3X1 NAND3X1_11 ( .A(_11_), .B(_16_), .C(_14_), .Y(_17_) );
AND2X2 AND2X2_8 ( .A(_17_), .B(_15_), .Y(w_C_6_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_18_) );
OR2X2 OR2X2_13 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_19_) );
NAND3X1 NAND3X1_12 ( .A(_15_), .B(_19_), .C(_17_), .Y(_20_) );
NAND2X1 NAND2X1_25 ( .A(_18_), .B(_20_), .Y(w_C_7_) );
BUFX2 BUFX2_8 ( .A(_21__0_), .Y(o_result[0]) );
BUFX2 BUFX2_9 ( .A(w_C_7_), .Y(_21__7_) );
BUFX2 BUFX2_10 ( .A(gnd), .Y(w_C_0_) );
endmodule
