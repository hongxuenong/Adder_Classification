module CSkipA_55bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [54:0] i_add_term1;
input [54:0] i_add_term2;
output [54:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

NAND2X1 NAND2X1_1 ( .A(_283_), .B(_287_), .Y(_0__22_) );
OAI21X1 OAI21X1_1 ( .A(_284_), .B(_281_), .C(_286_), .Y(_17__3_) );
INVX1 INVX1_1 ( .A(i_add_term1[20]), .Y(_288_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[20]), .B(_288_), .Y(_289_) );
INVX1 INVX1_2 ( .A(i_add_term2[20]), .Y(_290_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term1[20]), .B(_290_), .Y(_291_) );
INVX1 INVX1_3 ( .A(i_add_term1[21]), .Y(_292_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[21]), .B(_292_), .Y(_293_) );
INVX1 INVX1_4 ( .A(i_add_term2[21]), .Y(_294_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term1[21]), .B(_294_), .Y(_295_) );
OAI22X1 OAI22X1_1 ( .A(_289_), .B(_291_), .C(_293_), .D(_295_), .Y(_296_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_297_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_298_) );
NOR2X1 NOR2X1_6 ( .A(_297_), .B(_298_), .Y(_299_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_300_) );
NAND2X1 NAND2X1_2 ( .A(_299_), .B(_300_), .Y(_301_) );
NOR2X1 NOR2X1_7 ( .A(_296_), .B(_301_), .Y(_18_) );
INVX1 INVX1_5 ( .A(_16_), .Y(_302_) );
NAND2X1 NAND2X1_3 ( .A(gnd), .B(_18_), .Y(_303_) );
OAI21X1 OAI21X1_2 ( .A(_18_), .B(_302_), .C(_303_), .Y(w_cout_6_) );
INVX1 INVX1_6 ( .A(w_cout_6_), .Y(_307_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_308_) );
NAND2X1 NAND2X1_4 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_309_) );
NAND3X1 NAND3X1_1 ( .A(_307_), .B(_309_), .C(_308_), .Y(_310_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_304_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_305_) );
OAI21X1 OAI21X1_3 ( .A(_304_), .B(_305_), .C(w_cout_6_), .Y(_306_) );
NAND2X1 NAND2X1_5 ( .A(_306_), .B(_310_), .Y(_0__24_) );
OAI21X1 OAI21X1_4 ( .A(_307_), .B(_304_), .C(_309_), .Y(_20__1_) );
INVX1 INVX1_7 ( .A(_20__3_), .Y(_314_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_315_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_316_) );
NAND3X1 NAND3X1_2 ( .A(_314_), .B(_316_), .C(_315_), .Y(_317_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_311_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_312_) );
OAI21X1 OAI21X1_5 ( .A(_311_), .B(_312_), .C(_20__3_), .Y(_313_) );
NAND2X1 NAND2X1_7 ( .A(_313_), .B(_317_), .Y(_0__27_) );
OAI21X1 OAI21X1_6 ( .A(_314_), .B(_311_), .C(_316_), .Y(_19_) );
INVX1 INVX1_8 ( .A(_20__1_), .Y(_321_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_322_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_323_) );
NAND3X1 NAND3X1_3 ( .A(_321_), .B(_323_), .C(_322_), .Y(_324_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_318_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_319_) );
OAI21X1 OAI21X1_7 ( .A(_318_), .B(_319_), .C(_20__1_), .Y(_320_) );
NAND2X1 NAND2X1_9 ( .A(_320_), .B(_324_), .Y(_0__25_) );
OAI21X1 OAI21X1_8 ( .A(_321_), .B(_318_), .C(_323_), .Y(_20__2_) );
INVX1 INVX1_9 ( .A(_20__2_), .Y(_328_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_329_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_330_) );
NAND3X1 NAND3X1_4 ( .A(_328_), .B(_330_), .C(_329_), .Y(_331_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_325_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_326_) );
OAI21X1 OAI21X1_9 ( .A(_325_), .B(_326_), .C(_20__2_), .Y(_327_) );
NAND2X1 NAND2X1_11 ( .A(_327_), .B(_331_), .Y(_0__26_) );
OAI21X1 OAI21X1_10 ( .A(_328_), .B(_325_), .C(_330_), .Y(_20__3_) );
INVX1 INVX1_10 ( .A(i_add_term1[24]), .Y(_332_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[24]), .B(_332_), .Y(_333_) );
INVX1 INVX1_11 ( .A(i_add_term2[24]), .Y(_334_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term1[24]), .B(_334_), .Y(_335_) );
INVX1 INVX1_12 ( .A(i_add_term1[25]), .Y(_336_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[25]), .B(_336_), .Y(_337_) );
INVX1 INVX1_13 ( .A(i_add_term2[25]), .Y(_338_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term1[25]), .B(_338_), .Y(_339_) );
OAI22X1 OAI22X1_2 ( .A(_333_), .B(_335_), .C(_337_), .D(_339_), .Y(_340_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_341_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_342_) );
NOR2X1 NOR2X1_17 ( .A(_341_), .B(_342_), .Y(_343_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_344_) );
NAND2X1 NAND2X1_12 ( .A(_343_), .B(_344_), .Y(_345_) );
NOR2X1 NOR2X1_18 ( .A(_340_), .B(_345_), .Y(_21_) );
INVX1 INVX1_14 ( .A(_19_), .Y(_346_) );
NAND2X1 NAND2X1_13 ( .A(gnd), .B(_21_), .Y(_347_) );
OAI21X1 OAI21X1_11 ( .A(_21_), .B(_346_), .C(_347_), .Y(w_cout_7_) );
INVX1 INVX1_15 ( .A(w_cout_7_), .Y(_351_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_352_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_353_) );
NAND3X1 NAND3X1_5 ( .A(_351_), .B(_353_), .C(_352_), .Y(_354_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_348_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_349_) );
OAI21X1 OAI21X1_12 ( .A(_348_), .B(_349_), .C(w_cout_7_), .Y(_350_) );
NAND2X1 NAND2X1_15 ( .A(_350_), .B(_354_), .Y(_0__28_) );
OAI21X1 OAI21X1_13 ( .A(_351_), .B(_348_), .C(_353_), .Y(_23__1_) );
INVX1 INVX1_16 ( .A(_23__3_), .Y(_358_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_359_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_360_) );
NAND3X1 NAND3X1_6 ( .A(_358_), .B(_360_), .C(_359_), .Y(_361_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_355_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_356_) );
OAI21X1 OAI21X1_14 ( .A(_355_), .B(_356_), .C(_23__3_), .Y(_357_) );
NAND2X1 NAND2X1_17 ( .A(_357_), .B(_361_), .Y(_0__31_) );
OAI21X1 OAI21X1_15 ( .A(_358_), .B(_355_), .C(_360_), .Y(_22_) );
INVX1 INVX1_17 ( .A(_23__1_), .Y(_365_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_366_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_367_) );
NAND3X1 NAND3X1_7 ( .A(_365_), .B(_367_), .C(_366_), .Y(_368_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_362_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_363_) );
OAI21X1 OAI21X1_16 ( .A(_362_), .B(_363_), .C(_23__1_), .Y(_364_) );
NAND2X1 NAND2X1_19 ( .A(_364_), .B(_368_), .Y(_0__29_) );
OAI21X1 OAI21X1_17 ( .A(_365_), .B(_362_), .C(_367_), .Y(_23__2_) );
INVX1 INVX1_18 ( .A(_23__2_), .Y(_372_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_373_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_374_) );
NAND3X1 NAND3X1_8 ( .A(_372_), .B(_374_), .C(_373_), .Y(_375_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_369_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_370_) );
OAI21X1 OAI21X1_18 ( .A(_369_), .B(_370_), .C(_23__2_), .Y(_371_) );
NAND2X1 NAND2X1_21 ( .A(_371_), .B(_375_), .Y(_0__30_) );
OAI21X1 OAI21X1_19 ( .A(_372_), .B(_369_), .C(_374_), .Y(_23__3_) );
INVX1 INVX1_19 ( .A(i_add_term1[28]), .Y(_376_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[28]), .B(_376_), .Y(_377_) );
INVX1 INVX1_20 ( .A(i_add_term2[28]), .Y(_378_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term1[28]), .B(_378_), .Y(_379_) );
INVX1 INVX1_21 ( .A(i_add_term1[29]), .Y(_380_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[29]), .B(_380_), .Y(_381_) );
INVX1 INVX1_22 ( .A(i_add_term2[29]), .Y(_382_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term1[29]), .B(_382_), .Y(_383_) );
OAI22X1 OAI22X1_3 ( .A(_377_), .B(_379_), .C(_381_), .D(_383_), .Y(_384_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_385_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_386_) );
NOR2X1 NOR2X1_28 ( .A(_385_), .B(_386_), .Y(_387_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_388_) );
NAND2X1 NAND2X1_22 ( .A(_387_), .B(_388_), .Y(_389_) );
NOR2X1 NOR2X1_29 ( .A(_384_), .B(_389_), .Y(_24_) );
INVX1 INVX1_23 ( .A(_22_), .Y(_390_) );
NAND2X1 NAND2X1_23 ( .A(gnd), .B(_24_), .Y(_391_) );
OAI21X1 OAI21X1_20 ( .A(_24_), .B(_390_), .C(_391_), .Y(w_cout_8_) );
INVX1 INVX1_24 ( .A(w_cout_8_), .Y(_395_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_396_) );
NAND2X1 NAND2X1_24 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_397_) );
NAND3X1 NAND3X1_9 ( .A(_395_), .B(_397_), .C(_396_), .Y(_398_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_392_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_393_) );
OAI21X1 OAI21X1_21 ( .A(_392_), .B(_393_), .C(w_cout_8_), .Y(_394_) );
NAND2X1 NAND2X1_25 ( .A(_394_), .B(_398_), .Y(_0__32_) );
OAI21X1 OAI21X1_22 ( .A(_395_), .B(_392_), .C(_397_), .Y(_26__1_) );
INVX1 INVX1_25 ( .A(_26__3_), .Y(_402_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_403_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_404_) );
NAND3X1 NAND3X1_10 ( .A(_402_), .B(_404_), .C(_403_), .Y(_405_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_399_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_400_) );
OAI21X1 OAI21X1_23 ( .A(_399_), .B(_400_), .C(_26__3_), .Y(_401_) );
NAND2X1 NAND2X1_27 ( .A(_401_), .B(_405_), .Y(_0__35_) );
OAI21X1 OAI21X1_24 ( .A(_402_), .B(_399_), .C(_404_), .Y(_25_) );
INVX1 INVX1_26 ( .A(_26__1_), .Y(_409_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_410_) );
NAND2X1 NAND2X1_28 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_411_) );
NAND3X1 NAND3X1_11 ( .A(_409_), .B(_411_), .C(_410_), .Y(_412_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_406_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_407_) );
OAI21X1 OAI21X1_25 ( .A(_406_), .B(_407_), .C(_26__1_), .Y(_408_) );
NAND2X1 NAND2X1_29 ( .A(_408_), .B(_412_), .Y(_0__33_) );
OAI21X1 OAI21X1_26 ( .A(_409_), .B(_406_), .C(_411_), .Y(_26__2_) );
INVX1 INVX1_27 ( .A(_26__2_), .Y(_416_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_417_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_418_) );
NAND3X1 NAND3X1_12 ( .A(_416_), .B(_418_), .C(_417_), .Y(_419_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_413_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_414_) );
OAI21X1 OAI21X1_27 ( .A(_413_), .B(_414_), .C(_26__2_), .Y(_415_) );
NAND2X1 NAND2X1_31 ( .A(_415_), .B(_419_), .Y(_0__34_) );
OAI21X1 OAI21X1_28 ( .A(_416_), .B(_413_), .C(_418_), .Y(_26__3_) );
INVX1 INVX1_28 ( .A(i_add_term1[32]), .Y(_420_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[32]), .B(_420_), .Y(_421_) );
INVX1 INVX1_29 ( .A(i_add_term2[32]), .Y(_422_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term1[32]), .B(_422_), .Y(_423_) );
INVX1 INVX1_30 ( .A(i_add_term1[33]), .Y(_424_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[33]), .B(_424_), .Y(_425_) );
INVX1 INVX1_31 ( .A(i_add_term2[33]), .Y(_426_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term1[33]), .B(_426_), .Y(_427_) );
OAI22X1 OAI22X1_4 ( .A(_421_), .B(_423_), .C(_425_), .D(_427_), .Y(_428_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_429_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_430_) );
NOR2X1 NOR2X1_39 ( .A(_429_), .B(_430_), .Y(_431_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_432_) );
NAND2X1 NAND2X1_32 ( .A(_431_), .B(_432_), .Y(_433_) );
NOR2X1 NOR2X1_40 ( .A(_428_), .B(_433_), .Y(_27_) );
INVX1 INVX1_32 ( .A(_25_), .Y(_434_) );
NAND2X1 NAND2X1_33 ( .A(gnd), .B(_27_), .Y(_435_) );
OAI21X1 OAI21X1_29 ( .A(_27_), .B(_434_), .C(_435_), .Y(w_cout_9_) );
INVX1 INVX1_33 ( .A(w_cout_9_), .Y(_439_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_440_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_441_) );
NAND3X1 NAND3X1_13 ( .A(_439_), .B(_441_), .C(_440_), .Y(_442_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_436_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_437_) );
OAI21X1 OAI21X1_30 ( .A(_436_), .B(_437_), .C(w_cout_9_), .Y(_438_) );
NAND2X1 NAND2X1_35 ( .A(_438_), .B(_442_), .Y(_0__36_) );
OAI21X1 OAI21X1_31 ( .A(_439_), .B(_436_), .C(_441_), .Y(_29__1_) );
INVX1 INVX1_34 ( .A(_29__3_), .Y(_446_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_447_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_448_) );
NAND3X1 NAND3X1_14 ( .A(_446_), .B(_448_), .C(_447_), .Y(_449_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_443_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_444_) );
OAI21X1 OAI21X1_32 ( .A(_443_), .B(_444_), .C(_29__3_), .Y(_445_) );
NAND2X1 NAND2X1_37 ( .A(_445_), .B(_449_), .Y(_0__39_) );
OAI21X1 OAI21X1_33 ( .A(_446_), .B(_443_), .C(_448_), .Y(_28_) );
INVX1 INVX1_35 ( .A(_29__1_), .Y(_453_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_454_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_455_) );
NAND3X1 NAND3X1_15 ( .A(_453_), .B(_455_), .C(_454_), .Y(_456_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_450_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_451_) );
OAI21X1 OAI21X1_34 ( .A(_450_), .B(_451_), .C(_29__1_), .Y(_452_) );
NAND2X1 NAND2X1_39 ( .A(_452_), .B(_456_), .Y(_0__37_) );
OAI21X1 OAI21X1_35 ( .A(_453_), .B(_450_), .C(_455_), .Y(_29__2_) );
INVX1 INVX1_36 ( .A(_29__2_), .Y(_460_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_461_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_462_) );
NAND3X1 NAND3X1_16 ( .A(_460_), .B(_462_), .C(_461_), .Y(_463_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_457_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_458_) );
OAI21X1 OAI21X1_36 ( .A(_457_), .B(_458_), .C(_29__2_), .Y(_459_) );
NAND2X1 NAND2X1_41 ( .A(_459_), .B(_463_), .Y(_0__38_) );
OAI21X1 OAI21X1_37 ( .A(_460_), .B(_457_), .C(_462_), .Y(_29__3_) );
INVX1 INVX1_37 ( .A(i_add_term1[36]), .Y(_464_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[36]), .B(_464_), .Y(_465_) );
INVX1 INVX1_38 ( .A(i_add_term2[36]), .Y(_466_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term1[36]), .B(_466_), .Y(_467_) );
INVX1 INVX1_39 ( .A(i_add_term1[37]), .Y(_468_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[37]), .B(_468_), .Y(_469_) );
INVX1 INVX1_40 ( .A(i_add_term2[37]), .Y(_470_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term1[37]), .B(_470_), .Y(_471_) );
OAI22X1 OAI22X1_5 ( .A(_465_), .B(_467_), .C(_469_), .D(_471_), .Y(_472_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_473_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_474_) );
NOR2X1 NOR2X1_50 ( .A(_473_), .B(_474_), .Y(_475_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_476_) );
NAND2X1 NAND2X1_42 ( .A(_475_), .B(_476_), .Y(_477_) );
NOR2X1 NOR2X1_51 ( .A(_472_), .B(_477_), .Y(_30_) );
INVX1 INVX1_41 ( .A(_28_), .Y(_478_) );
NAND2X1 NAND2X1_43 ( .A(gnd), .B(_30_), .Y(_479_) );
OAI21X1 OAI21X1_38 ( .A(_30_), .B(_478_), .C(_479_), .Y(w_cout_10_) );
INVX1 INVX1_42 ( .A(w_cout_10_), .Y(_483_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_484_) );
NAND2X1 NAND2X1_44 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_485_) );
NAND3X1 NAND3X1_17 ( .A(_483_), .B(_485_), .C(_484_), .Y(_486_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_480_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_481_) );
OAI21X1 OAI21X1_39 ( .A(_480_), .B(_481_), .C(w_cout_10_), .Y(_482_) );
NAND2X1 NAND2X1_45 ( .A(_482_), .B(_486_), .Y(_0__40_) );
OAI21X1 OAI21X1_40 ( .A(_483_), .B(_480_), .C(_485_), .Y(_32__1_) );
INVX1 INVX1_43 ( .A(_32__3_), .Y(_490_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_491_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_492_) );
NAND3X1 NAND3X1_18 ( .A(_490_), .B(_492_), .C(_491_), .Y(_493_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_487_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_488_) );
OAI21X1 OAI21X1_41 ( .A(_487_), .B(_488_), .C(_32__3_), .Y(_489_) );
NAND2X1 NAND2X1_47 ( .A(_489_), .B(_493_), .Y(_0__43_) );
OAI21X1 OAI21X1_42 ( .A(_490_), .B(_487_), .C(_492_), .Y(_31_) );
INVX1 INVX1_44 ( .A(_32__1_), .Y(_497_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_498_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_499_) );
NAND3X1 NAND3X1_19 ( .A(_497_), .B(_499_), .C(_498_), .Y(_500_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_494_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_495_) );
OAI21X1 OAI21X1_43 ( .A(_494_), .B(_495_), .C(_32__1_), .Y(_496_) );
NAND2X1 NAND2X1_49 ( .A(_496_), .B(_500_), .Y(_0__41_) );
OAI21X1 OAI21X1_44 ( .A(_497_), .B(_494_), .C(_499_), .Y(_32__2_) );
INVX1 INVX1_45 ( .A(_32__2_), .Y(_504_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_505_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_506_) );
NAND3X1 NAND3X1_20 ( .A(_504_), .B(_506_), .C(_505_), .Y(_507_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_501_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_502_) );
OAI21X1 OAI21X1_45 ( .A(_501_), .B(_502_), .C(_32__2_), .Y(_503_) );
NAND2X1 NAND2X1_51 ( .A(_503_), .B(_507_), .Y(_0__42_) );
OAI21X1 OAI21X1_46 ( .A(_504_), .B(_501_), .C(_506_), .Y(_32__3_) );
INVX1 INVX1_46 ( .A(i_add_term1[40]), .Y(_508_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[40]), .B(_508_), .Y(_509_) );
INVX1 INVX1_47 ( .A(i_add_term2[40]), .Y(_510_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term1[40]), .B(_510_), .Y(_511_) );
INVX1 INVX1_48 ( .A(i_add_term1[41]), .Y(_512_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[41]), .B(_512_), .Y(_513_) );
INVX1 INVX1_49 ( .A(i_add_term2[41]), .Y(_514_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term1[41]), .B(_514_), .Y(_515_) );
OAI22X1 OAI22X1_6 ( .A(_509_), .B(_511_), .C(_513_), .D(_515_), .Y(_516_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_517_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_518_) );
NOR2X1 NOR2X1_61 ( .A(_517_), .B(_518_), .Y(_519_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_520_) );
NAND2X1 NAND2X1_52 ( .A(_519_), .B(_520_), .Y(_521_) );
NOR2X1 NOR2X1_62 ( .A(_516_), .B(_521_), .Y(_33_) );
INVX1 INVX1_50 ( .A(_31_), .Y(_522_) );
NAND2X1 NAND2X1_53 ( .A(gnd), .B(_33_), .Y(_523_) );
OAI21X1 OAI21X1_47 ( .A(_33_), .B(_522_), .C(_523_), .Y(w_cout_11_) );
INVX1 INVX1_51 ( .A(w_cout_11_), .Y(_527_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_528_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_529_) );
NAND3X1 NAND3X1_21 ( .A(_527_), .B(_529_), .C(_528_), .Y(_530_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_524_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_525_) );
OAI21X1 OAI21X1_48 ( .A(_524_), .B(_525_), .C(w_cout_11_), .Y(_526_) );
NAND2X1 NAND2X1_55 ( .A(_526_), .B(_530_), .Y(_0__44_) );
OAI21X1 OAI21X1_49 ( .A(_527_), .B(_524_), .C(_529_), .Y(_35__1_) );
INVX1 INVX1_52 ( .A(_35__3_), .Y(_534_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_535_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_536_) );
NAND3X1 NAND3X1_22 ( .A(_534_), .B(_536_), .C(_535_), .Y(_537_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_531_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_532_) );
OAI21X1 OAI21X1_50 ( .A(_531_), .B(_532_), .C(_35__3_), .Y(_533_) );
NAND2X1 NAND2X1_57 ( .A(_533_), .B(_537_), .Y(_0__47_) );
OAI21X1 OAI21X1_51 ( .A(_534_), .B(_531_), .C(_536_), .Y(_34_) );
INVX1 INVX1_53 ( .A(_35__1_), .Y(_541_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_542_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_543_) );
NAND3X1 NAND3X1_23 ( .A(_541_), .B(_543_), .C(_542_), .Y(_544_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_538_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_539_) );
OAI21X1 OAI21X1_52 ( .A(_538_), .B(_539_), .C(_35__1_), .Y(_540_) );
NAND2X1 NAND2X1_59 ( .A(_540_), .B(_544_), .Y(_0__45_) );
OAI21X1 OAI21X1_53 ( .A(_541_), .B(_538_), .C(_543_), .Y(_35__2_) );
INVX1 INVX1_54 ( .A(_35__2_), .Y(_548_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_549_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_550_) );
NAND3X1 NAND3X1_24 ( .A(_548_), .B(_550_), .C(_549_), .Y(_551_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_545_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_546_) );
OAI21X1 OAI21X1_54 ( .A(_545_), .B(_546_), .C(_35__2_), .Y(_547_) );
NAND2X1 NAND2X1_61 ( .A(_547_), .B(_551_), .Y(_0__46_) );
OAI21X1 OAI21X1_55 ( .A(_548_), .B(_545_), .C(_550_), .Y(_35__3_) );
INVX1 INVX1_55 ( .A(i_add_term1[44]), .Y(_552_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[44]), .B(_552_), .Y(_553_) );
INVX1 INVX1_56 ( .A(i_add_term2[44]), .Y(_554_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term1[44]), .B(_554_), .Y(_555_) );
INVX1 INVX1_57 ( .A(i_add_term1[45]), .Y(_556_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[45]), .B(_556_), .Y(_557_) );
INVX1 INVX1_58 ( .A(i_add_term2[45]), .Y(_558_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term1[45]), .B(_558_), .Y(_559_) );
OAI22X1 OAI22X1_7 ( .A(_553_), .B(_555_), .C(_557_), .D(_559_), .Y(_560_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_561_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_562_) );
NOR2X1 NOR2X1_72 ( .A(_561_), .B(_562_), .Y(_563_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_564_) );
NAND2X1 NAND2X1_62 ( .A(_563_), .B(_564_), .Y(_565_) );
NOR2X1 NOR2X1_73 ( .A(_560_), .B(_565_), .Y(_36_) );
INVX1 INVX1_59 ( .A(_34_), .Y(_566_) );
NAND2X1 NAND2X1_63 ( .A(gnd), .B(_36_), .Y(_567_) );
OAI21X1 OAI21X1_56 ( .A(_36_), .B(_566_), .C(_567_), .Y(w_cout_12_) );
INVX1 INVX1_60 ( .A(w_cout_12_), .Y(_571_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_572_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_573_) );
NAND3X1 NAND3X1_25 ( .A(_571_), .B(_573_), .C(_572_), .Y(_574_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_568_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_569_) );
OAI21X1 OAI21X1_57 ( .A(_568_), .B(_569_), .C(w_cout_12_), .Y(_570_) );
NAND2X1 NAND2X1_65 ( .A(_570_), .B(_574_), .Y(_0__48_) );
OAI21X1 OAI21X1_58 ( .A(_571_), .B(_568_), .C(_573_), .Y(_38__1_) );
INVX1 INVX1_61 ( .A(_38__3_), .Y(_578_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_579_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_580_) );
NAND3X1 NAND3X1_26 ( .A(_578_), .B(_580_), .C(_579_), .Y(_581_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_575_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_576_) );
OAI21X1 OAI21X1_59 ( .A(_575_), .B(_576_), .C(_38__3_), .Y(_577_) );
NAND2X1 NAND2X1_67 ( .A(_577_), .B(_581_), .Y(_0__51_) );
OAI21X1 OAI21X1_60 ( .A(_578_), .B(_575_), .C(_580_), .Y(_37_) );
INVX1 INVX1_62 ( .A(_38__1_), .Y(_585_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_586_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_587_) );
NAND3X1 NAND3X1_27 ( .A(_585_), .B(_587_), .C(_586_), .Y(_588_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_582_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_583_) );
OAI21X1 OAI21X1_61 ( .A(_582_), .B(_583_), .C(_38__1_), .Y(_584_) );
NAND2X1 NAND2X1_69 ( .A(_584_), .B(_588_), .Y(_0__49_) );
OAI21X1 OAI21X1_62 ( .A(_585_), .B(_582_), .C(_587_), .Y(_38__2_) );
INVX1 INVX1_63 ( .A(_38__2_), .Y(_592_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_593_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_594_) );
NAND3X1 NAND3X1_28 ( .A(_592_), .B(_594_), .C(_593_), .Y(_595_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_589_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_590_) );
OAI21X1 OAI21X1_63 ( .A(_589_), .B(_590_), .C(_38__2_), .Y(_591_) );
NAND2X1 NAND2X1_71 ( .A(_591_), .B(_595_), .Y(_0__50_) );
OAI21X1 OAI21X1_64 ( .A(_592_), .B(_589_), .C(_594_), .Y(_38__3_) );
INVX1 INVX1_64 ( .A(i_add_term1[48]), .Y(_596_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[48]), .B(_596_), .Y(_597_) );
INVX1 INVX1_65 ( .A(i_add_term2[48]), .Y(_598_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term1[48]), .B(_598_), .Y(_599_) );
INVX1 INVX1_66 ( .A(i_add_term1[49]), .Y(_600_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[49]), .B(_600_), .Y(_601_) );
INVX1 INVX1_67 ( .A(i_add_term2[49]), .Y(_602_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term1[49]), .B(_602_), .Y(_603_) );
OAI22X1 OAI22X1_8 ( .A(_597_), .B(_599_), .C(_601_), .D(_603_), .Y(_604_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_605_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_606_) );
NOR2X1 NOR2X1_83 ( .A(_605_), .B(_606_), .Y(_607_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_608_) );
NAND2X1 NAND2X1_72 ( .A(_607_), .B(_608_), .Y(_609_) );
NOR2X1 NOR2X1_84 ( .A(_604_), .B(_609_), .Y(_39_) );
INVX1 INVX1_68 ( .A(_37_), .Y(_610_) );
NAND2X1 NAND2X1_73 ( .A(gnd), .B(_39_), .Y(_611_) );
OAI21X1 OAI21X1_65 ( .A(_39_), .B(_610_), .C(_611_), .Y(cskip3_inst_cin) );
INVX1 INVX1_69 ( .A(cskip3_inst_cin), .Y(_615_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_616_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_617_) );
NAND3X1 NAND3X1_29 ( .A(_615_), .B(_617_), .C(_616_), .Y(_618_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_612_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_613_) );
OAI21X1 OAI21X1_66 ( .A(_612_), .B(_613_), .C(cskip3_inst_cin), .Y(_614_) );
NAND2X1 NAND2X1_75 ( .A(_614_), .B(_618_), .Y(cskip3_inst_rca0_fa0_o_sum) );
OAI21X1 OAI21X1_67 ( .A(_615_), .B(_612_), .C(_617_), .Y(cskip3_inst_rca0_fa0_o_carry) );
INVX1 INVX1_70 ( .A(cskip3_inst_rca0_fa0_o_carry), .Y(_622_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_623_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_624_) );
NAND3X1 NAND3X1_30 ( .A(_622_), .B(_624_), .C(_623_), .Y(_625_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_619_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_620_) );
OAI21X1 OAI21X1_68 ( .A(_619_), .B(_620_), .C(cskip3_inst_rca0_fa0_o_carry), .Y(_621_) );
NAND2X1 NAND2X1_77 ( .A(_621_), .B(_625_), .Y(cskip3_inst_rca0_fa1_o_sum) );
OAI21X1 OAI21X1_69 ( .A(_622_), .B(_619_), .C(_624_), .Y(cskip3_inst_rca0_fa1_o_carry) );
INVX1 INVX1_71 ( .A(cskip3_inst_rca0_fa1_o_carry), .Y(_629_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_630_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_631_) );
NAND3X1 NAND3X1_31 ( .A(_629_), .B(_631_), .C(_630_), .Y(_632_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_626_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_627_) );
OAI21X1 OAI21X1_70 ( .A(_626_), .B(_627_), .C(cskip3_inst_rca0_fa1_o_carry), .Y(_628_) );
NAND2X1 NAND2X1_79 ( .A(_628_), .B(_632_), .Y(cskip3_inst_rca0_fa2_o_sum) );
OAI21X1 OAI21X1_71 ( .A(_629_), .B(_626_), .C(_631_), .Y(cskip3_inst_cout0) );
OR2X2 OR2X2_32 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_636_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_637_) );
NAND2X1 NAND2X1_81 ( .A(_637_), .B(_636_), .Y(_633_) );
XNOR2X1 XNOR2X1_1 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_634_) );
XNOR2X1 XNOR2X1_2 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_635_) );
NOR3X1 NOR3X1_1 ( .A(_633_), .B(_634_), .C(_635_), .Y(cskip3_inst_skip0_P) );
INVX1 INVX1_72 ( .A(cskip3_inst_cout0), .Y(_638_) );
NAND2X1 NAND2X1_82 ( .A(gnd), .B(cskip3_inst_skip0_P), .Y(_639_) );
OAI21X1 OAI21X1_72 ( .A(cskip3_inst_skip0_P), .B(_638_), .C(_639_), .Y(w_cout_14_) );
BUFX2 BUFX2_1 ( .A(w_cout_14_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .A(cskip3_inst_rca0_fa0_o_sum), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .A(cskip3_inst_rca0_fa1_o_sum), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .A(cskip3_inst_rca0_fa2_o_sum), .Y(sum[54]) );
INVX1 INVX1_73 ( .A(gnd), .Y(_43_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_44_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_45_) );
NAND3X1 NAND3X1_32 ( .A(_43_), .B(_45_), .C(_44_), .Y(_46_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_40_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_41_) );
OAI21X1 OAI21X1_73 ( .A(_40_), .B(_41_), .C(gnd), .Y(_42_) );
NAND2X1 NAND2X1_84 ( .A(_42_), .B(_46_), .Y(_0__0_) );
OAI21X1 OAI21X1_74 ( .A(_43_), .B(_40_), .C(_45_), .Y(_2__1_) );
INVX1 INVX1_74 ( .A(_2__3_), .Y(_50_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_51_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_52_) );
NAND3X1 NAND3X1_33 ( .A(_50_), .B(_52_), .C(_51_), .Y(_53_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_47_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_48_) );
OAI21X1 OAI21X1_75 ( .A(_47_), .B(_48_), .C(_2__3_), .Y(_49_) );
NAND2X1 NAND2X1_86 ( .A(_49_), .B(_53_), .Y(_0__3_) );
OAI21X1 OAI21X1_76 ( .A(_50_), .B(_47_), .C(_52_), .Y(_1_) );
INVX1 INVX1_75 ( .A(_2__1_), .Y(_57_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_58_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_59_) );
NAND3X1 NAND3X1_34 ( .A(_57_), .B(_59_), .C(_58_), .Y(_60_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_54_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_55_) );
OAI21X1 OAI21X1_77 ( .A(_54_), .B(_55_), .C(_2__1_), .Y(_56_) );
NAND2X1 NAND2X1_88 ( .A(_56_), .B(_60_), .Y(_0__1_) );
OAI21X1 OAI21X1_78 ( .A(_57_), .B(_54_), .C(_59_), .Y(_2__2_) );
INVX1 INVX1_76 ( .A(_2__2_), .Y(_64_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_65_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_66_) );
NAND3X1 NAND3X1_35 ( .A(_64_), .B(_66_), .C(_65_), .Y(_67_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_61_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_62_) );
OAI21X1 OAI21X1_79 ( .A(_61_), .B(_62_), .C(_2__2_), .Y(_63_) );
NAND2X1 NAND2X1_90 ( .A(_63_), .B(_67_), .Y(_0__2_) );
OAI21X1 OAI21X1_80 ( .A(_64_), .B(_61_), .C(_66_), .Y(_2__3_) );
INVX1 INVX1_77 ( .A(i_add_term1[0]), .Y(_68_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[0]), .B(_68_), .Y(_69_) );
INVX1 INVX1_78 ( .A(i_add_term2[0]), .Y(_70_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term1[0]), .B(_70_), .Y(_71_) );
INVX1 INVX1_79 ( .A(i_add_term1[1]), .Y(_72_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[1]), .B(_72_), .Y(_73_) );
INVX1 INVX1_80 ( .A(i_add_term2[1]), .Y(_74_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term1[1]), .B(_74_), .Y(_75_) );
OAI22X1 OAI22X1_9 ( .A(_69_), .B(_71_), .C(_73_), .D(_75_), .Y(_76_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_77_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_78_) );
NOR2X1 NOR2X1_97 ( .A(_77_), .B(_78_), .Y(_79_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_80_) );
NAND2X1 NAND2X1_91 ( .A(_79_), .B(_80_), .Y(_81_) );
NOR2X1 NOR2X1_98 ( .A(_76_), .B(_81_), .Y(_3_) );
INVX1 INVX1_81 ( .A(_1_), .Y(_82_) );
NAND2X1 NAND2X1_92 ( .A(gnd), .B(_3_), .Y(_83_) );
OAI21X1 OAI21X1_81 ( .A(_3_), .B(_82_), .C(_83_), .Y(w_cout_1_) );
INVX1 INVX1_82 ( .A(w_cout_1_), .Y(_87_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_88_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_89_) );
NAND3X1 NAND3X1_36 ( .A(_87_), .B(_89_), .C(_88_), .Y(_90_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_84_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_85_) );
OAI21X1 OAI21X1_82 ( .A(_84_), .B(_85_), .C(w_cout_1_), .Y(_86_) );
NAND2X1 NAND2X1_94 ( .A(_86_), .B(_90_), .Y(_0__4_) );
OAI21X1 OAI21X1_83 ( .A(_87_), .B(_84_), .C(_89_), .Y(_5__1_) );
INVX1 INVX1_83 ( .A(_5__3_), .Y(_94_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_95_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_96_) );
NAND3X1 NAND3X1_37 ( .A(_94_), .B(_96_), .C(_95_), .Y(_97_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_91_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_92_) );
OAI21X1 OAI21X1_84 ( .A(_91_), .B(_92_), .C(_5__3_), .Y(_93_) );
NAND2X1 NAND2X1_96 ( .A(_93_), .B(_97_), .Y(_0__7_) );
OAI21X1 OAI21X1_85 ( .A(_94_), .B(_91_), .C(_96_), .Y(_4_) );
INVX1 INVX1_84 ( .A(_5__1_), .Y(_101_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_102_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_103_) );
NAND3X1 NAND3X1_38 ( .A(_101_), .B(_103_), .C(_102_), .Y(_104_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_98_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_99_) );
OAI21X1 OAI21X1_86 ( .A(_98_), .B(_99_), .C(_5__1_), .Y(_100_) );
NAND2X1 NAND2X1_98 ( .A(_100_), .B(_104_), .Y(_0__5_) );
OAI21X1 OAI21X1_87 ( .A(_101_), .B(_98_), .C(_103_), .Y(_5__2_) );
INVX1 INVX1_85 ( .A(_5__2_), .Y(_108_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_109_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_110_) );
NAND3X1 NAND3X1_39 ( .A(_108_), .B(_110_), .C(_109_), .Y(_111_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_105_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_106_) );
OAI21X1 OAI21X1_88 ( .A(_105_), .B(_106_), .C(_5__2_), .Y(_107_) );
NAND2X1 NAND2X1_100 ( .A(_107_), .B(_111_), .Y(_0__6_) );
OAI21X1 OAI21X1_89 ( .A(_108_), .B(_105_), .C(_110_), .Y(_5__3_) );
INVX1 INVX1_86 ( .A(i_add_term1[4]), .Y(_112_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[4]), .B(_112_), .Y(_113_) );
INVX1 INVX1_87 ( .A(i_add_term2[4]), .Y(_114_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term1[4]), .B(_114_), .Y(_115_) );
INVX1 INVX1_88 ( .A(i_add_term1[5]), .Y(_116_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[5]), .B(_116_), .Y(_117_) );
INVX1 INVX1_89 ( .A(i_add_term2[5]), .Y(_118_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term1[5]), .B(_118_), .Y(_119_) );
OAI22X1 OAI22X1_10 ( .A(_113_), .B(_115_), .C(_117_), .D(_119_), .Y(_120_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_121_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_122_) );
NOR2X1 NOR2X1_108 ( .A(_121_), .B(_122_), .Y(_123_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_124_) );
NAND2X1 NAND2X1_101 ( .A(_123_), .B(_124_), .Y(_125_) );
NOR2X1 NOR2X1_109 ( .A(_120_), .B(_125_), .Y(_6_) );
INVX1 INVX1_90 ( .A(_4_), .Y(_126_) );
NAND2X1 NAND2X1_102 ( .A(gnd), .B(_6_), .Y(_127_) );
OAI21X1 OAI21X1_90 ( .A(_6_), .B(_126_), .C(_127_), .Y(w_cout_2_) );
INVX1 INVX1_91 ( .A(w_cout_2_), .Y(_131_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_132_) );
NAND2X1 NAND2X1_103 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_133_) );
NAND3X1 NAND3X1_40 ( .A(_131_), .B(_133_), .C(_132_), .Y(_134_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_128_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_129_) );
OAI21X1 OAI21X1_91 ( .A(_128_), .B(_129_), .C(w_cout_2_), .Y(_130_) );
NAND2X1 NAND2X1_104 ( .A(_130_), .B(_134_), .Y(_0__8_) );
OAI21X1 OAI21X1_92 ( .A(_131_), .B(_128_), .C(_133_), .Y(_8__1_) );
INVX1 INVX1_92 ( .A(_8__3_), .Y(_138_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_139_) );
NAND2X1 NAND2X1_105 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_140_) );
NAND3X1 NAND3X1_41 ( .A(_138_), .B(_140_), .C(_139_), .Y(_141_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_135_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_136_) );
OAI21X1 OAI21X1_93 ( .A(_135_), .B(_136_), .C(_8__3_), .Y(_137_) );
NAND2X1 NAND2X1_106 ( .A(_137_), .B(_141_), .Y(_0__11_) );
OAI21X1 OAI21X1_94 ( .A(_138_), .B(_135_), .C(_140_), .Y(_7_) );
INVX1 INVX1_93 ( .A(_8__1_), .Y(_145_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_146_) );
NAND2X1 NAND2X1_107 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_147_) );
NAND3X1 NAND3X1_42 ( .A(_145_), .B(_147_), .C(_146_), .Y(_148_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_142_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_143_) );
OAI21X1 OAI21X1_95 ( .A(_142_), .B(_143_), .C(_8__1_), .Y(_144_) );
NAND2X1 NAND2X1_108 ( .A(_144_), .B(_148_), .Y(_0__9_) );
OAI21X1 OAI21X1_96 ( .A(_145_), .B(_142_), .C(_147_), .Y(_8__2_) );
INVX1 INVX1_94 ( .A(_8__2_), .Y(_152_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_153_) );
NAND2X1 NAND2X1_109 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_154_) );
NAND3X1 NAND3X1_43 ( .A(_152_), .B(_154_), .C(_153_), .Y(_155_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_149_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_150_) );
OAI21X1 OAI21X1_97 ( .A(_149_), .B(_150_), .C(_8__2_), .Y(_151_) );
NAND2X1 NAND2X1_110 ( .A(_151_), .B(_155_), .Y(_0__10_) );
OAI21X1 OAI21X1_98 ( .A(_152_), .B(_149_), .C(_154_), .Y(_8__3_) );
INVX1 INVX1_95 ( .A(i_add_term1[8]), .Y(_156_) );
NOR2X1 NOR2X1_114 ( .A(i_add_term2[8]), .B(_156_), .Y(_157_) );
INVX1 INVX1_96 ( .A(i_add_term2[8]), .Y(_158_) );
NOR2X1 NOR2X1_115 ( .A(i_add_term1[8]), .B(_158_), .Y(_159_) );
INVX1 INVX1_97 ( .A(i_add_term1[9]), .Y(_160_) );
NOR2X1 NOR2X1_116 ( .A(i_add_term2[9]), .B(_160_), .Y(_161_) );
INVX1 INVX1_98 ( .A(i_add_term2[9]), .Y(_162_) );
NOR2X1 NOR2X1_117 ( .A(i_add_term1[9]), .B(_162_), .Y(_163_) );
OAI22X1 OAI22X1_11 ( .A(_157_), .B(_159_), .C(_161_), .D(_163_), .Y(_164_) );
NOR2X1 NOR2X1_118 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_165_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_166_) );
NOR2X1 NOR2X1_119 ( .A(_165_), .B(_166_), .Y(_167_) );
XOR2X1 XOR2X1_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_168_) );
NAND2X1 NAND2X1_111 ( .A(_167_), .B(_168_), .Y(_169_) );
NOR2X1 NOR2X1_120 ( .A(_164_), .B(_169_), .Y(_9_) );
INVX1 INVX1_99 ( .A(_7_), .Y(_170_) );
NAND2X1 NAND2X1_112 ( .A(gnd), .B(_9_), .Y(_171_) );
OAI21X1 OAI21X1_99 ( .A(_9_), .B(_170_), .C(_171_), .Y(w_cout_3_) );
INVX1 INVX1_100 ( .A(w_cout_3_), .Y(_175_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_176_) );
NAND2X1 NAND2X1_113 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_177_) );
NAND3X1 NAND3X1_44 ( .A(_175_), .B(_177_), .C(_176_), .Y(_178_) );
NOR2X1 NOR2X1_121 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_172_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_173_) );
OAI21X1 OAI21X1_100 ( .A(_172_), .B(_173_), .C(w_cout_3_), .Y(_174_) );
NAND2X1 NAND2X1_114 ( .A(_174_), .B(_178_), .Y(_0__12_) );
OAI21X1 OAI21X1_101 ( .A(_175_), .B(_172_), .C(_177_), .Y(_11__1_) );
INVX1 INVX1_101 ( .A(_11__3_), .Y(_182_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_183_) );
NAND2X1 NAND2X1_115 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_184_) );
NAND3X1 NAND3X1_45 ( .A(_182_), .B(_184_), .C(_183_), .Y(_185_) );
NOR2X1 NOR2X1_122 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_179_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_180_) );
OAI21X1 OAI21X1_102 ( .A(_179_), .B(_180_), .C(_11__3_), .Y(_181_) );
NAND2X1 NAND2X1_116 ( .A(_181_), .B(_185_), .Y(_0__15_) );
OAI21X1 OAI21X1_103 ( .A(_182_), .B(_179_), .C(_184_), .Y(_10_) );
INVX1 INVX1_102 ( .A(_11__1_), .Y(_189_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_190_) );
NAND2X1 NAND2X1_117 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_191_) );
NAND3X1 NAND3X1_46 ( .A(_189_), .B(_191_), .C(_190_), .Y(_192_) );
NOR2X1 NOR2X1_123 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_186_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_187_) );
OAI21X1 OAI21X1_104 ( .A(_186_), .B(_187_), .C(_11__1_), .Y(_188_) );
NAND2X1 NAND2X1_118 ( .A(_188_), .B(_192_), .Y(_0__13_) );
OAI21X1 OAI21X1_105 ( .A(_189_), .B(_186_), .C(_191_), .Y(_11__2_) );
INVX1 INVX1_103 ( .A(_11__2_), .Y(_196_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_197_) );
NAND2X1 NAND2X1_119 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_198_) );
NAND3X1 NAND3X1_47 ( .A(_196_), .B(_198_), .C(_197_), .Y(_199_) );
NOR2X1 NOR2X1_124 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_193_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_194_) );
OAI21X1 OAI21X1_106 ( .A(_193_), .B(_194_), .C(_11__2_), .Y(_195_) );
NAND2X1 NAND2X1_120 ( .A(_195_), .B(_199_), .Y(_0__14_) );
OAI21X1 OAI21X1_107 ( .A(_196_), .B(_193_), .C(_198_), .Y(_11__3_) );
INVX1 INVX1_104 ( .A(i_add_term1[12]), .Y(_200_) );
NOR2X1 NOR2X1_125 ( .A(i_add_term2[12]), .B(_200_), .Y(_201_) );
INVX1 INVX1_105 ( .A(i_add_term2[12]), .Y(_202_) );
NOR2X1 NOR2X1_126 ( .A(i_add_term1[12]), .B(_202_), .Y(_203_) );
INVX1 INVX1_106 ( .A(i_add_term1[13]), .Y(_204_) );
NOR2X1 NOR2X1_127 ( .A(i_add_term2[13]), .B(_204_), .Y(_205_) );
INVX1 INVX1_107 ( .A(i_add_term2[13]), .Y(_206_) );
NOR2X1 NOR2X1_128 ( .A(i_add_term1[13]), .B(_206_), .Y(_207_) );
OAI22X1 OAI22X1_12 ( .A(_201_), .B(_203_), .C(_205_), .D(_207_), .Y(_208_) );
NOR2X1 NOR2X1_129 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_209_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_210_) );
NOR2X1 NOR2X1_130 ( .A(_209_), .B(_210_), .Y(_211_) );
XOR2X1 XOR2X1_12 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_212_) );
NAND2X1 NAND2X1_121 ( .A(_211_), .B(_212_), .Y(_213_) );
NOR2X1 NOR2X1_131 ( .A(_208_), .B(_213_), .Y(_12_) );
INVX1 INVX1_108 ( .A(_10_), .Y(_214_) );
NAND2X1 NAND2X1_122 ( .A(gnd), .B(_12_), .Y(_215_) );
OAI21X1 OAI21X1_108 ( .A(_12_), .B(_214_), .C(_215_), .Y(w_cout_4_) );
INVX1 INVX1_109 ( .A(w_cout_4_), .Y(_219_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_220_) );
NAND2X1 NAND2X1_123 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_221_) );
NAND3X1 NAND3X1_48 ( .A(_219_), .B(_221_), .C(_220_), .Y(_222_) );
NOR2X1 NOR2X1_132 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_216_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_217_) );
OAI21X1 OAI21X1_109 ( .A(_216_), .B(_217_), .C(w_cout_4_), .Y(_218_) );
NAND2X1 NAND2X1_124 ( .A(_218_), .B(_222_), .Y(_0__16_) );
OAI21X1 OAI21X1_110 ( .A(_219_), .B(_216_), .C(_221_), .Y(_14__1_) );
INVX1 INVX1_110 ( .A(_14__3_), .Y(_226_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_227_) );
NAND2X1 NAND2X1_125 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_228_) );
NAND3X1 NAND3X1_49 ( .A(_226_), .B(_228_), .C(_227_), .Y(_229_) );
NOR2X1 NOR2X1_133 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_223_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_224_) );
OAI21X1 OAI21X1_111 ( .A(_223_), .B(_224_), .C(_14__3_), .Y(_225_) );
NAND2X1 NAND2X1_126 ( .A(_225_), .B(_229_), .Y(_0__19_) );
OAI21X1 OAI21X1_112 ( .A(_226_), .B(_223_), .C(_228_), .Y(_13_) );
INVX1 INVX1_111 ( .A(_14__1_), .Y(_233_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_234_) );
NAND2X1 NAND2X1_127 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_235_) );
NAND3X1 NAND3X1_50 ( .A(_233_), .B(_235_), .C(_234_), .Y(_236_) );
NOR2X1 NOR2X1_134 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_230_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_231_) );
OAI21X1 OAI21X1_113 ( .A(_230_), .B(_231_), .C(_14__1_), .Y(_232_) );
NAND2X1 NAND2X1_128 ( .A(_232_), .B(_236_), .Y(_0__17_) );
OAI21X1 OAI21X1_114 ( .A(_233_), .B(_230_), .C(_235_), .Y(_14__2_) );
INVX1 INVX1_112 ( .A(_14__2_), .Y(_240_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_241_) );
NAND2X1 NAND2X1_129 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_242_) );
NAND3X1 NAND3X1_51 ( .A(_240_), .B(_242_), .C(_241_), .Y(_243_) );
NOR2X1 NOR2X1_135 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_237_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_238_) );
OAI21X1 OAI21X1_115 ( .A(_237_), .B(_238_), .C(_14__2_), .Y(_239_) );
NAND2X1 NAND2X1_130 ( .A(_239_), .B(_243_), .Y(_0__18_) );
OAI21X1 OAI21X1_116 ( .A(_240_), .B(_237_), .C(_242_), .Y(_14__3_) );
INVX1 INVX1_113 ( .A(i_add_term1[16]), .Y(_244_) );
NOR2X1 NOR2X1_136 ( .A(i_add_term2[16]), .B(_244_), .Y(_245_) );
INVX1 INVX1_114 ( .A(i_add_term2[16]), .Y(_246_) );
NOR2X1 NOR2X1_137 ( .A(i_add_term1[16]), .B(_246_), .Y(_247_) );
INVX1 INVX1_115 ( .A(i_add_term1[17]), .Y(_248_) );
NOR2X1 NOR2X1_138 ( .A(i_add_term2[17]), .B(_248_), .Y(_249_) );
INVX1 INVX1_116 ( .A(i_add_term2[17]), .Y(_250_) );
NOR2X1 NOR2X1_139 ( .A(i_add_term1[17]), .B(_250_), .Y(_251_) );
OAI22X1 OAI22X1_13 ( .A(_245_), .B(_247_), .C(_249_), .D(_251_), .Y(_252_) );
NOR2X1 NOR2X1_140 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_253_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_254_) );
NOR2X1 NOR2X1_141 ( .A(_253_), .B(_254_), .Y(_255_) );
XOR2X1 XOR2X1_13 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_256_) );
NAND2X1 NAND2X1_131 ( .A(_255_), .B(_256_), .Y(_257_) );
NOR2X1 NOR2X1_142 ( .A(_252_), .B(_257_), .Y(_15_) );
INVX1 INVX1_117 ( .A(_13_), .Y(_258_) );
NAND2X1 NAND2X1_132 ( .A(gnd), .B(_15_), .Y(_259_) );
OAI21X1 OAI21X1_117 ( .A(_15_), .B(_258_), .C(_259_), .Y(w_cout_5_) );
INVX1 INVX1_118 ( .A(w_cout_5_), .Y(_263_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_264_) );
NAND2X1 NAND2X1_133 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_265_) );
NAND3X1 NAND3X1_52 ( .A(_263_), .B(_265_), .C(_264_), .Y(_266_) );
NOR2X1 NOR2X1_143 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_260_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_261_) );
OAI21X1 OAI21X1_118 ( .A(_260_), .B(_261_), .C(w_cout_5_), .Y(_262_) );
NAND2X1 NAND2X1_134 ( .A(_262_), .B(_266_), .Y(_0__20_) );
OAI21X1 OAI21X1_119 ( .A(_263_), .B(_260_), .C(_265_), .Y(_17__1_) );
INVX1 INVX1_119 ( .A(_17__3_), .Y(_270_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_271_) );
NAND2X1 NAND2X1_135 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_272_) );
NAND3X1 NAND3X1_53 ( .A(_270_), .B(_272_), .C(_271_), .Y(_273_) );
NOR2X1 NOR2X1_144 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_267_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_268_) );
OAI21X1 OAI21X1_120 ( .A(_267_), .B(_268_), .C(_17__3_), .Y(_269_) );
NAND2X1 NAND2X1_136 ( .A(_269_), .B(_273_), .Y(_0__23_) );
OAI21X1 OAI21X1_121 ( .A(_270_), .B(_267_), .C(_272_), .Y(_16_) );
INVX1 INVX1_120 ( .A(_17__1_), .Y(_277_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_278_) );
NAND2X1 NAND2X1_137 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_279_) );
NAND3X1 NAND3X1_54 ( .A(_277_), .B(_279_), .C(_278_), .Y(_280_) );
NOR2X1 NOR2X1_145 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_274_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_275_) );
OAI21X1 OAI21X1_122 ( .A(_274_), .B(_275_), .C(_17__1_), .Y(_276_) );
NAND2X1 NAND2X1_138 ( .A(_276_), .B(_280_), .Y(_0__21_) );
OAI21X1 OAI21X1_123 ( .A(_277_), .B(_274_), .C(_279_), .Y(_17__2_) );
INVX1 INVX1_121 ( .A(_17__2_), .Y(_284_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_285_) );
NAND2X1 NAND2X1_139 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_286_) );
NAND3X1 NAND3X1_55 ( .A(_284_), .B(_286_), .C(_285_), .Y(_287_) );
NOR2X1 NOR2X1_146 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_281_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_282_) );
OAI21X1 OAI21X1_124 ( .A(_281_), .B(_282_), .C(_17__2_), .Y(_283_) );
BUFX2 BUFX2_57 ( .A(cskip3_inst_rca0_fa0_o_sum), .Y(_0__52_) );
BUFX2 BUFX2_58 ( .A(cskip3_inst_rca0_fa1_o_sum), .Y(_0__53_) );
BUFX2 BUFX2_59 ( .A(cskip3_inst_rca0_fa2_o_sum), .Y(_0__54_) );
BUFX2 BUFX2_60 ( .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_61 ( .A(cskip3_inst_cin), .Y(w_cout_13_) );
endmodule
