module CSkipA_5bit ( gnd, vdd, i_add_term1, i_add_term2, sum, cout);

input gnd, vdd;
output cout;
input [4:0] i_add_term1;
input [4:0] i_add_term2;
output [4:0] sum;

NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_27_), .Y(_1__0_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_21_), .C(_26_), .Y(_3__1_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_3__1_), .Y(_31_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_32_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_33_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_33_), .C(_32_), .Y(_34_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_28_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_29_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_29_), .C(_3__1_), .Y(_30_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_34_), .Y(_1__1_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_28_), .C(_33_), .Y(_3__2_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_3__2_), .Y(_38_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_39_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_40_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_40_), .C(_39_), .Y(_41_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_35_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_36_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_36_), .C(_3__2_), .Y(_37_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_41_), .Y(_1__2_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_35_), .C(_40_), .Y(_3__3_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_3__3_), .Y(_45_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_46_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_47_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_47_), .C(_46_), .Y(_48_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_42_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_43_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_43_), .C(_3__3_), .Y(_44_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_48_), .Y(_1__3_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_42_), .C(_47_), .Y(_2_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_cin), .Y(_52_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_53_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_54_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_54_), .C(_53_), .Y(_55_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_49_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_50_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_50_), .C(cskip1_inst_cin), .Y(_51_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_55_), .Y(cskip1_inst_sum) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_49_), .C(_54_), .Y(cskip1_inst_rca0_w_CARRY_1_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_rca0_w_CARRY_1_), .Y(_57_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_58_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_56_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_56_), .C(_58_), .Y(cskip1_inst_rca0_w_CARRY_2_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_rca0_w_CARRY_2_), .Y(_60_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_61_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_59_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_59_), .C(_61_), .Y(cskip1_inst_rca0_w_CARRY_3_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_rca0_w_CARRY_3_), .Y(_63_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_64_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_62_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_62_), .C(_64_), .Y(cskip1_inst_cout0) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_65_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_66_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_66_), .Y(cskip1_inst_skip0_P) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_cout0), .Y(_67_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(cskip1_inst_skip0_P), .Y(_68_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_skip0_P), .B(_67_), .C(_68_), .Y(_0_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(cout) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_1__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_1__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_1__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_1__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_sum), .Y(sum[4]) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .Y(_5_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(_5_), .Y(_6_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .Y(_7_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[0]), .B(_7_), .Y(_8_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .Y(_9_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(_9_), .Y(_10_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .Y(_11_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term1[1]), .B(_11_), .Y(_12_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_8_), .C(_10_), .D(_12_), .Y(_13_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_14_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_15_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_15_), .Y(_16_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_17_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_17_), .Y(_18_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_18_), .Y(_4_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_2_), .Y(_19_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_4_), .Y(_20_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_19_), .C(_20_), .Y(cskip1_inst_cin) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_24_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_25_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_26_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_26_), .C(_25_), .Y(_27_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_21_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_22_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_22_), .C(gnd), .Y(_23_) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_sum), .Y(_1__4_) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_3__0_) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_2_), .Y(_3__4_) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_cin), .Y(cskip1_inst_rca0_w_CARRY_0_) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(cskip1_inst_cout0), .Y(cskip1_inst_rca0_w_CARRY_4_) );
endmodule
