module cla_59bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [58:0] i_add1;
input [58:0] i_add2;
output [59:0] o_result;

OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .C(_276_), .Y(_277_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_277_), .Y(w_C_44_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .Y(_278_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add1[44]), .Y(_279_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_279_), .Y(_280_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_280_), .Y(_281_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_282_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_282_), .Y(_283_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_284_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_284_), .Y(_285_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_283_), .B(_285_), .C(_276_), .Y(_286_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_281_), .Y(_287_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_287_), .Y(w_C_45_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_288_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_288_), .Y(_289_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_289_), .C(_286_), .Y(_290_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .C(_290_), .Y(_291_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_291_), .Y(w_C_46_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .Y(_292_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add1[46]), .Y(_293_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_292_), .B(_293_), .Y(_294_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_294_), .Y(_295_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_296_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_296_), .Y(_297_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_298_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_298_), .Y(_299_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_299_), .C(_290_), .Y(_300_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_295_), .Y(_301_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_301_), .Y(w_C_47_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_302_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_302_), .Y(_303_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_303_), .C(_300_), .Y(_304_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .C(_304_), .Y(_305_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_305_), .Y(w_C_48_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_306_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_307_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_305_), .C(_306_), .Y(w_C_49_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_308_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_309_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_309_), .Y(_310_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_307_), .Y(_311_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_311_), .C(_304_), .Y(_312_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_313_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_313_), .C(_312_), .Y(_314_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_308_), .Y(w_C_50_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .Y(_315_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add1[50]), .Y(_316_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_316_), .Y(_317_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_317_), .C(_314_), .Y(_318_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_316_), .C(_318_), .Y(w_C_51_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .Y(_319_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add1[51]), .Y(_320_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_320_), .Y(_321_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_322_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_323_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_323_), .C(_318_), .Y(_324_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_321_), .Y(w_C_52_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .Y(_325_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add1[52]), .Y(_326_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_326_), .Y(_327_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_327_), .C(_324_), .Y(_328_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_326_), .C(_328_), .Y(w_C_53_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .Y(_329_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add1[53]), .Y(_330_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .C(w_C_53_), .Y(_331_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_330_), .C(_331_), .Y(w_C_54_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_330_), .Y(_332_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_332_), .Y(_333_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_334_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_334_), .Y(_335_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_335_), .C(_331_), .Y(_336_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .C(_336_), .Y(_337_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_337_), .Y(w_C_55_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_338_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_339_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_337_), .C(_338_), .Y(w_C_56_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_340_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_339_), .Y(_341_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_342_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_342_), .Y(_343_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_326_), .Y(_344_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_344_), .Y(_345_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_333_), .C(_328_), .Y(_346_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_347_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_347_), .Y(_348_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_348_), .C(_346_), .Y(_349_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_335_), .B(_338_), .C(_349_), .Y(_350_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_351_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_351_), .C(_350_), .Y(_352_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_352_), .Y(w_C_57_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_353_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_354_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_354_), .C(_352_), .Y(_355_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_353_), .Y(w_C_58_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_356_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_357_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_357_), .C(_355_), .Y(_358_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_358_), .Y(w_C_59_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_7_), .Y(w_C_3_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .Y(_8_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add1[3]), .Y(_9_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_9_), .Y(_10_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_11_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_11_), .C(_7_), .Y(_12_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_10_), .Y(w_C_4_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_14_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_14_), .C(_12_), .Y(_15_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_15_), .Y(w_C_5_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_16_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_17_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_18_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_18_), .C(_15_), .Y(_19_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_17_), .Y(w_C_6_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .Y(_20_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add1[6]), .Y(_21_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_23_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_23_), .C(_19_), .Y(_24_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .C(_24_), .Y(w_C_7_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_25_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(_26_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .Y(_27_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(_28_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .Y(_29_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add1[7]), .Y(_30_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_30_), .Y(_31_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_31_), .Y(_32_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_32_), .C(_24_), .Y(_33_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_26_), .Y(w_C_8_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .Y(_34_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add1[8]), .Y(_35_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_36_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_36_), .Y(_37_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_37_), .C(_33_), .Y(_38_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_35_), .C(_38_), .Y(w_C_9_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_35_), .Y(_39_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_39_), .Y(_40_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_41_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_41_), .Y(_42_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_42_), .C(_38_), .Y(_43_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .C(_43_), .Y(_44_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_44_), .Y(w_C_10_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .Y(_45_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add1[10]), .Y(_46_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_47_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_47_), .Y(_48_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_49_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_49_), .Y(_50_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_50_), .C(_43_), .Y(_51_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_46_), .C(_51_), .Y(w_C_11_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_46_), .Y(_52_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_52_), .Y(_53_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_54_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_54_), .Y(_55_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_55_), .C(_51_), .Y(_56_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .C(_56_), .Y(_57_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_57_), .Y(w_C_12_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .Y(_58_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add1[12]), .Y(_59_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_60_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_60_), .Y(_61_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_62_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_62_), .Y(_63_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_63_), .C(_56_), .Y(_64_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_59_), .C(_64_), .Y(w_C_13_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_59_), .Y(_65_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_65_), .Y(_66_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_67_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_67_), .Y(_68_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_68_), .C(_64_), .Y(_69_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .C(_69_), .Y(_70_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_70_), .Y(w_C_14_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .Y(_71_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add1[14]), .Y(_72_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_73_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_73_), .Y(_74_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_75_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(_75_), .Y(_76_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_76_), .C(_69_), .Y(_77_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_72_), .C(_77_), .Y(w_C_15_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_359__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_359__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_359__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_359__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_359__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_359__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_359__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_359__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_359__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_359__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_359__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_359__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_359__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_359__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_359__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_359__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_359__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_359__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_359__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_359__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_359__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_359__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_359__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_359__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_359__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_359__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_359__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_359__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_359__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_359__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_359__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_359__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_359__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_359__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_359__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_359__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_359__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_359__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_359__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_359__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_359__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_359__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_359__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_359__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_359__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_359__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_359__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_359__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_359__48_), .Y(o_result[48]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_359__49_), .Y(o_result[49]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_359__50_), .Y(o_result[50]) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_359__51_), .Y(o_result[51]) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(_359__52_), .Y(o_result[52]) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(_359__53_), .Y(o_result[53]) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(_359__54_), .Y(o_result[54]) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_359__55_), .Y(o_result[55]) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_359__56_), .Y(o_result[56]) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_359__57_), .Y(o_result[57]) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_359__58_), .Y(o_result[58]) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(w_C_59_), .Y(o_result[59]) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_363_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_364_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_365_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_365_), .C(_364_), .Y(_366_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_360_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_361_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_361_), .C(w_C_4_), .Y(_362_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_366_), .Y(_359__4_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_370_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_371_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_372_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_372_), .C(_371_), .Y(_373_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_367_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_368_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_368_), .C(w_C_5_), .Y(_369_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_373_), .Y(_359__5_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_377_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_378_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_379_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_379_), .C(_378_), .Y(_380_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_374_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_375_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_375_), .C(w_C_6_), .Y(_376_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_380_), .Y(_359__6_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_384_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_385_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_386_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_386_), .C(_385_), .Y(_387_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_381_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_382_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_382_), .C(w_C_7_), .Y(_383_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_387_), .Y(_359__7_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_391_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_392_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_393_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_393_), .C(_392_), .Y(_394_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_388_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_389_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(_389_), .C(w_C_8_), .Y(_390_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_394_), .Y(_359__8_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_398_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_399_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_400_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_400_), .C(_399_), .Y(_401_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_395_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_396_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_396_), .C(w_C_9_), .Y(_397_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_401_), .Y(_359__9_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_405_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_406_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_407_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_407_), .C(_406_), .Y(_408_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_402_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_403_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_403_), .C(w_C_10_), .Y(_404_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_408_), .Y(_359__10_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_412_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_413_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_414_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_414_), .C(_413_), .Y(_415_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_409_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_410_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_410_), .C(w_C_11_), .Y(_411_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_415_), .Y(_359__11_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(w_C_12_), .Y(_419_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_420_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_421_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_421_), .C(_420_), .Y(_422_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_416_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_417_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_417_), .C(w_C_12_), .Y(_418_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_422_), .Y(_359__12_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(w_C_13_), .Y(_426_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_427_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_428_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_428_), .C(_427_), .Y(_429_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_423_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_424_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_424_), .C(w_C_13_), .Y(_425_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(_429_), .Y(_359__13_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(w_C_14_), .Y(_433_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_434_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_435_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_435_), .C(_434_), .Y(_436_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_430_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_431_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_431_), .C(w_C_14_), .Y(_432_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_432_), .B(_436_), .Y(_359__14_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(_440_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_441_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_442_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_442_), .C(_441_), .Y(_443_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_437_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_438_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_438_), .C(w_C_15_), .Y(_439_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_443_), .Y(_359__15_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(w_C_16_), .Y(_447_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_448_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_449_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_449_), .C(_448_), .Y(_450_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_444_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_445_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_445_), .C(w_C_16_), .Y(_446_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(_450_), .Y(_359__16_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(w_C_17_), .Y(_454_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_455_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_456_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_454_), .B(_456_), .C(_455_), .Y(_457_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_451_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_452_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_452_), .C(w_C_17_), .Y(_453_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(_457_), .Y(_359__17_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(w_C_18_), .Y(_461_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_462_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_463_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_463_), .C(_462_), .Y(_464_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_458_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_459_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_459_), .C(w_C_18_), .Y(_460_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_464_), .Y(_359__18_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(w_C_19_), .Y(_468_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_469_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_470_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_468_), .B(_470_), .C(_469_), .Y(_471_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_465_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_466_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_466_), .C(w_C_19_), .Y(_467_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_467_), .B(_471_), .Y(_359__19_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(w_C_20_), .Y(_475_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_476_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_477_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_477_), .C(_476_), .Y(_478_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_472_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_473_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_473_), .C(w_C_20_), .Y(_474_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_474_), .B(_478_), .Y(_359__20_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(w_C_21_), .Y(_482_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_483_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_484_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_482_), .B(_484_), .C(_483_), .Y(_485_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_479_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_480_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_480_), .C(w_C_21_), .Y(_481_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_485_), .Y(_359__21_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(w_C_22_), .Y(_489_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_490_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_491_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_491_), .C(_490_), .Y(_492_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_486_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_487_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_487_), .C(w_C_22_), .Y(_488_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_492_), .Y(_359__22_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(w_C_23_), .Y(_496_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_497_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_498_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_498_), .C(_497_), .Y(_499_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_493_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_494_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_494_), .C(w_C_23_), .Y(_495_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_495_), .B(_499_), .Y(_359__23_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(w_C_24_), .Y(_503_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_504_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_505_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_505_), .C(_504_), .Y(_506_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_500_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_501_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_501_), .C(w_C_24_), .Y(_502_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_502_), .B(_506_), .Y(_359__24_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(w_C_25_), .Y(_510_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_511_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_512_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_512_), .C(_511_), .Y(_513_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_507_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_508_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_508_), .C(w_C_25_), .Y(_509_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_513_), .Y(_359__25_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(w_C_26_), .Y(_517_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_518_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_519_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_517_), .B(_519_), .C(_518_), .Y(_520_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_514_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_515_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_514_), .B(_515_), .C(w_C_26_), .Y(_516_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_520_), .Y(_359__26_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(w_C_27_), .Y(_524_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_525_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_526_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_526_), .C(_525_), .Y(_527_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_521_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_522_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_522_), .C(w_C_27_), .Y(_523_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_527_), .Y(_359__27_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(w_C_28_), .Y(_531_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_532_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_533_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_533_), .C(_532_), .Y(_534_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_528_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_529_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_529_), .C(w_C_28_), .Y(_530_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_534_), .Y(_359__28_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(w_C_29_), .Y(_538_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_539_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_540_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_538_), .B(_540_), .C(_539_), .Y(_541_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_535_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_536_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_536_), .C(w_C_29_), .Y(_537_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_541_), .Y(_359__29_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(w_C_30_), .Y(_545_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_546_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_547_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_545_), .B(_547_), .C(_546_), .Y(_548_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_542_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_543_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_542_), .B(_543_), .C(w_C_30_), .Y(_544_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_548_), .Y(_359__30_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(w_C_31_), .Y(_552_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_553_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_554_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_552_), .B(_554_), .C(_553_), .Y(_555_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_549_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_550_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(_550_), .C(w_C_31_), .Y(_551_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_551_), .B(_555_), .Y(_359__31_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(w_C_32_), .Y(_559_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_560_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_561_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_561_), .C(_560_), .Y(_562_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_556_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_557_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_556_), .B(_557_), .C(w_C_32_), .Y(_558_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_562_), .Y(_359__32_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(w_C_33_), .Y(_566_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_567_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_568_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_568_), .C(_567_), .Y(_569_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_563_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_564_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(_564_), .C(w_C_33_), .Y(_565_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_569_), .Y(_359__33_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(w_C_34_), .Y(_573_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_574_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_575_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_575_), .C(_574_), .Y(_576_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_570_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_571_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_571_), .C(w_C_34_), .Y(_572_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_576_), .Y(_359__34_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(w_C_35_), .Y(_580_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_581_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_582_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(_582_), .C(_581_), .Y(_583_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_577_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_578_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_578_), .C(w_C_35_), .Y(_579_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_583_), .Y(_359__35_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(w_C_36_), .Y(_587_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_588_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_589_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(_589_), .C(_588_), .Y(_590_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_584_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_585_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_585_), .C(w_C_36_), .Y(_586_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_586_), .B(_590_), .Y(_359__36_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(w_C_37_), .Y(_594_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_595_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_596_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_594_), .B(_596_), .C(_595_), .Y(_597_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_591_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_592_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_592_), .C(w_C_37_), .Y(_593_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_597_), .Y(_359__37_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(w_C_38_), .Y(_601_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_602_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_603_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_601_), .B(_603_), .C(_602_), .Y(_604_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_598_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_599_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_598_), .B(_599_), .C(w_C_38_), .Y(_600_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_604_), .Y(_359__38_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(w_C_39_), .Y(_608_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_609_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_610_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_608_), .B(_610_), .C(_609_), .Y(_611_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_605_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_606_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_606_), .C(w_C_39_), .Y(_607_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_611_), .Y(_359__39_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(w_C_40_), .Y(_615_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_616_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_617_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_615_), .B(_617_), .C(_616_), .Y(_618_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_612_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_613_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_612_), .B(_613_), .C(w_C_40_), .Y(_614_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_618_), .Y(_359__40_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(w_C_41_), .Y(_622_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_623_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_624_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_622_), .B(_624_), .C(_623_), .Y(_625_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_619_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_620_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_620_), .C(w_C_41_), .Y(_621_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_625_), .Y(_359__41_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(w_C_42_), .Y(_629_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_630_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_631_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_629_), .B(_631_), .C(_630_), .Y(_632_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_626_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_627_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_627_), .C(w_C_42_), .Y(_628_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_628_), .B(_632_), .Y(_359__42_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(w_C_43_), .Y(_636_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_637_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_638_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_636_), .B(_638_), .C(_637_), .Y(_639_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_633_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_634_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_634_), .C(w_C_43_), .Y(_635_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_639_), .Y(_359__43_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(w_C_44_), .Y(_643_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_644_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_645_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_645_), .C(_644_), .Y(_646_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_640_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[44]), .B(i_add1[44]), .Y(_641_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(_641_), .C(w_C_44_), .Y(_642_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_642_), .B(_646_), .Y(_359__44_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(w_C_45_), .Y(_650_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_651_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_652_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(_652_), .C(_651_), .Y(_653_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_647_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[45]), .B(i_add1[45]), .Y(_648_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_647_), .B(_648_), .C(w_C_45_), .Y(_649_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_653_), .Y(_359__45_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(w_C_46_), .Y(_657_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_658_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_659_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_657_), .B(_659_), .C(_658_), .Y(_660_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_654_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[46]), .B(i_add1[46]), .Y(_655_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_655_), .C(w_C_46_), .Y(_656_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_656_), .B(_660_), .Y(_359__46_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(w_C_47_), .Y(_664_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_665_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_666_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_664_), .B(_666_), .C(_665_), .Y(_667_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_661_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[47]), .B(i_add1[47]), .Y(_662_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_661_), .B(_662_), .C(w_C_47_), .Y(_663_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(_667_), .Y(_359__47_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(w_C_48_), .Y(_671_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_672_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_673_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_671_), .B(_673_), .C(_672_), .Y(_674_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_668_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[48]), .B(i_add1[48]), .Y(_669_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_669_), .C(w_C_48_), .Y(_670_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(_674_), .Y(_359__48_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(w_C_49_), .Y(_678_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_679_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_680_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_680_), .C(_679_), .Y(_681_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_675_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[49]), .B(i_add1[49]), .Y(_676_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_676_), .C(w_C_49_), .Y(_677_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_681_), .Y(_359__49_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(w_C_50_), .Y(_685_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_686_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_687_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_687_), .C(_686_), .Y(_688_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_682_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[50]), .B(i_add1[50]), .Y(_683_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_682_), .B(_683_), .C(w_C_50_), .Y(_684_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_684_), .B(_688_), .Y(_359__50_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(w_C_51_), .Y(_692_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_693_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_694_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_692_), .B(_694_), .C(_693_), .Y(_695_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_689_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[51]), .B(i_add1[51]), .Y(_690_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_690_), .C(w_C_51_), .Y(_691_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_691_), .B(_695_), .Y(_359__51_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(w_C_52_), .Y(_699_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_700_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_701_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_701_), .C(_700_), .Y(_702_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_696_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[52]), .B(i_add1[52]), .Y(_697_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_697_), .C(w_C_52_), .Y(_698_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_702_), .Y(_359__52_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(w_C_53_), .Y(_706_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_707_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_708_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_708_), .C(_707_), .Y(_709_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_703_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[53]), .B(i_add1[53]), .Y(_704_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_704_), .C(w_C_53_), .Y(_705_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_705_), .B(_709_), .Y(_359__53_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(w_C_54_), .Y(_713_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_714_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_715_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_715_), .C(_714_), .Y(_716_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_710_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[54]), .B(i_add1[54]), .Y(_711_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_710_), .B(_711_), .C(w_C_54_), .Y(_712_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_712_), .B(_716_), .Y(_359__54_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(w_C_55_), .Y(_720_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_721_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_722_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_720_), .B(_722_), .C(_721_), .Y(_723_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_717_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[55]), .B(i_add1[55]), .Y(_718_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_717_), .B(_718_), .C(w_C_55_), .Y(_719_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(_723_), .Y(_359__55_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(w_C_56_), .Y(_727_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_728_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_729_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_727_), .B(_729_), .C(_728_), .Y(_730_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_724_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[56]), .B(i_add1[56]), .Y(_725_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_724_), .B(_725_), .C(w_C_56_), .Y(_726_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_726_), .B(_730_), .Y(_359__56_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(w_C_57_), .Y(_734_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_735_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_736_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_734_), .B(_736_), .C(_735_), .Y(_737_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_731_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[57]), .B(i_add1[57]), .Y(_732_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_731_), .B(_732_), .C(w_C_57_), .Y(_733_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_733_), .B(_737_), .Y(_359__57_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(w_C_58_), .Y(_741_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_742_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_743_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_741_), .B(_743_), .C(_742_), .Y(_744_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_738_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[58]), .B(i_add1[58]), .Y(_739_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_738_), .B(_739_), .C(w_C_58_), .Y(_740_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_740_), .B(_744_), .Y(_359__58_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_748_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_749_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_750_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_748_), .B(_750_), .C(_749_), .Y(_751_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_745_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_746_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_745_), .B(_746_), .C(gnd), .Y(_747_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_747_), .B(_751_), .Y(_359__0_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_755_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_756_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_757_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_757_), .C(_756_), .Y(_758_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_752_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_753_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(_753_), .C(w_C_1_), .Y(_754_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_754_), .B(_758_), .Y(_359__1_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_762_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_763_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_764_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_762_), .B(_764_), .C(_763_), .Y(_765_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_759_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_760_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_759_), .B(_760_), .C(w_C_2_), .Y(_761_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_761_), .B(_765_), .Y(_359__2_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_769_) );
OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_770_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_771_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_769_), .B(_771_), .C(_770_), .Y(_772_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_766_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_767_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_766_), .B(_767_), .C(w_C_3_), .Y(_768_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_768_), .B(_772_), .Y(_359__3_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_72_), .Y(_78_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(_78_), .Y(_79_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_80_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(_80_), .Y(_81_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_81_), .C(_77_), .Y(_82_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .C(_82_), .Y(_83_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(_83_), .Y(w_C_16_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .Y(_84_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(i_add1[16]), .Y(_85_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_86_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(_86_), .Y(_87_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_88_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(_88_), .Y(_89_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_89_), .C(_82_), .Y(_90_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_85_), .C(_90_), .Y(w_C_17_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_85_), .Y(_91_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(_91_), .Y(_92_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_93_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(_93_), .Y(_94_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_94_), .C(_90_), .Y(_95_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .C(_95_), .Y(_96_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(_96_), .Y(w_C_18_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .Y(_97_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(i_add1[18]), .Y(_98_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_99_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(_99_), .Y(_100_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_101_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(_101_), .Y(_102_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_102_), .C(_95_), .Y(_103_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_98_), .C(_103_), .Y(w_C_19_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_98_), .Y(_104_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(_104_), .Y(_105_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_106_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(_106_), .Y(_107_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_107_), .C(_103_), .Y(_108_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .C(_108_), .Y(_109_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(_109_), .Y(w_C_20_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .Y(_110_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(i_add1[20]), .Y(_111_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_111_), .Y(_112_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(_112_), .Y(_113_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_114_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(_114_), .Y(_115_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_116_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(_116_), .Y(_117_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_117_), .C(_108_), .Y(_118_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_113_), .Y(_119_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(_119_), .Y(w_C_21_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_120_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(_120_), .Y(_121_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_121_), .C(_118_), .Y(_122_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .C(_122_), .Y(_123_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(_123_), .Y(w_C_22_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .Y(_124_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(i_add1[22]), .Y(_125_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_125_), .Y(_126_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(_126_), .Y(_127_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_128_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(_128_), .Y(_129_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_130_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(_130_), .Y(_131_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_129_), .B(_131_), .C(_122_), .Y(_132_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_127_), .Y(_133_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(_133_), .Y(w_C_23_) );
AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_134_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(_134_), .Y(_135_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_135_), .C(_132_), .Y(_136_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .C(_136_), .Y(_137_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(_137_), .Y(w_C_24_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .Y(_138_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(i_add1[24]), .Y(_139_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_139_), .Y(_140_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(_140_), .Y(_141_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_142_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(_142_), .Y(_143_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_144_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(_144_), .Y(_145_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_145_), .C(_136_), .Y(_146_) );
AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_141_), .Y(_147_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(_147_), .Y(w_C_25_) );
AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_148_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(_148_), .Y(_149_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_149_), .C(_146_), .Y(_150_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .C(_150_), .Y(_151_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(_151_), .Y(w_C_26_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .Y(_152_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(i_add1[26]), .Y(_153_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_153_), .Y(_154_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(_154_), .Y(_155_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_156_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_157_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_158_) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(_158_), .Y(_159_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_159_), .C(_150_), .Y(_160_) );
AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_155_), .Y(_161_) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(_161_), .Y(w_C_27_) );
AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_162_) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(_162_), .Y(_163_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_163_), .C(_160_), .Y(_164_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .C(_164_), .Y(_165_) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(_165_), .Y(w_C_28_) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .Y(_166_) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(i_add1[28]), .Y(_167_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_167_), .Y(_168_) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(_168_), .Y(_169_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_170_) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(_170_), .Y(_171_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_172_) );
INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(_172_), .Y(_173_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_173_), .C(_164_), .Y(_174_) );
AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_169_), .Y(_175_) );
INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(_175_), .Y(w_C_29_) );
AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_176_) );
INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(_176_), .Y(_177_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_177_), .C(_174_), .Y(_178_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .C(_178_), .Y(_179_) );
INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(_179_), .Y(w_C_30_) );
INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .Y(_180_) );
INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(i_add1[30]), .Y(_181_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_181_), .Y(_182_) );
INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(_182_), .Y(_183_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_184_) );
INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(_184_), .Y(_185_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_186_) );
INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(_186_), .Y(_187_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_187_), .C(_178_), .Y(_188_) );
AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_183_), .Y(_189_) );
INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(_189_), .Y(w_C_31_) );
AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_190_) );
INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(_190_), .Y(_191_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_191_), .C(_188_), .Y(_192_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .C(_192_), .Y(_193_) );
INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(_193_), .Y(w_C_32_) );
INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .Y(_194_) );
INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(i_add1[32]), .Y(_195_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_195_), .Y(_196_) );
INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(_196_), .Y(_197_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_198_) );
INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(_198_), .Y(_199_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_200_) );
INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(_200_), .Y(_201_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_201_), .C(_192_), .Y(_202_) );
AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_197_), .Y(_203_) );
INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(_203_), .Y(w_C_33_) );
AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_204_) );
INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(_204_), .Y(_205_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_205_), .C(_202_), .Y(_206_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .C(_206_), .Y(_207_) );
INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(_207_), .Y(w_C_34_) );
INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .Y(_208_) );
INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(i_add1[34]), .Y(_209_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_209_), .Y(_210_) );
INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(_210_), .Y(_211_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_212_) );
INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(_212_), .Y(_213_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_214_) );
INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(_214_), .Y(_215_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_215_), .C(_206_), .Y(_216_) );
AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_211_), .Y(_217_) );
INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(_217_), .Y(w_C_35_) );
AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_218_) );
INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(_218_), .Y(_219_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_219_), .C(_216_), .Y(_220_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .C(_220_), .Y(_221_) );
INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(_221_), .Y(w_C_36_) );
INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .Y(_222_) );
INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(i_add1[36]), .Y(_223_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_223_), .Y(_224_) );
INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(_224_), .Y(_225_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_226_) );
INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(_226_), .Y(_227_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_228_) );
INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(_228_), .Y(_229_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_229_), .C(_220_), .Y(_230_) );
AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_225_), .Y(_231_) );
INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(_231_), .Y(w_C_37_) );
AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_232_) );
INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(_232_), .Y(_233_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_233_), .C(_230_), .Y(_234_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .C(_234_), .Y(_235_) );
INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(_235_), .Y(w_C_38_) );
INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .Y(_236_) );
INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(i_add1[38]), .Y(_237_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_237_), .Y(_238_) );
INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(_238_), .Y(_239_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_240_) );
INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(_240_), .Y(_241_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_242_) );
INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(_242_), .Y(_243_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_243_), .C(_234_), .Y(_244_) );
AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_239_), .Y(_245_) );
INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(_245_), .Y(w_C_39_) );
AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_246_) );
INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(_246_), .Y(_247_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_247_), .C(_244_), .Y(_248_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .C(_248_), .Y(_249_) );
INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(_249_), .Y(w_C_40_) );
INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .Y(_250_) );
INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(i_add1[40]), .Y(_251_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_251_), .Y(_252_) );
INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(_252_), .Y(_253_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_254_) );
INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(_254_), .Y(_255_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_256_) );
INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(_256_), .Y(_257_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_257_), .C(_248_), .Y(_258_) );
AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_253_), .Y(_259_) );
INVX1 INVX1_233 ( .gnd(gnd), .vdd(vdd), .A(_259_), .Y(w_C_41_) );
AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_260_) );
INVX1 INVX1_234 ( .gnd(gnd), .vdd(vdd), .A(_260_), .Y(_261_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_253_), .B(_261_), .C(_258_), .Y(_262_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .C(_262_), .Y(_263_) );
INVX1 INVX1_235 ( .gnd(gnd), .vdd(vdd), .A(_263_), .Y(w_C_42_) );
INVX1 INVX1_236 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .Y(_264_) );
INVX1 INVX1_237 ( .gnd(gnd), .vdd(vdd), .A(i_add1[42]), .Y(_265_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_265_), .Y(_266_) );
INVX1 INVX1_238 ( .gnd(gnd), .vdd(vdd), .A(_266_), .Y(_267_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_268_) );
INVX1 INVX1_239 ( .gnd(gnd), .vdd(vdd), .A(_268_), .Y(_269_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_270_) );
INVX1 INVX1_240 ( .gnd(gnd), .vdd(vdd), .A(_270_), .Y(_271_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_271_), .C(_262_), .Y(_272_) );
AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_267_), .Y(_273_) );
INVX1 INVX1_241 ( .gnd(gnd), .vdd(vdd), .A(_273_), .Y(w_C_43_) );
AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_274_) );
INVX1 INVX1_242 ( .gnd(gnd), .vdd(vdd), .A(_274_), .Y(_275_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_275_), .C(_272_), .Y(_276_) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(w_C_59_), .Y(_359__59_) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
