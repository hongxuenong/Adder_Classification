module CSkipA_20bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [19:0] i_add_term1;
input [19:0] i_add_term2;
output [19:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX2 BUFX2_1 ( .A(w_cout_4_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
INVX1 INVX1_1 ( .A(skip0_cin_next), .Y(_16_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_17_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_18_) );
NAND3X1 NAND3X1_1 ( .A(_16_), .B(_18_), .C(_17_), .Y(_19_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_13_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_14_) );
OAI21X1 OAI21X1_1 ( .A(_13_), .B(_14_), .C(skip0_cin_next), .Y(_15_) );
NAND2X1 NAND2X1_2 ( .A(_15_), .B(_19_), .Y(_0__4_) );
OAI21X1 OAI21X1_2 ( .A(_16_), .B(_13_), .C(_18_), .Y(_2__1_) );
INVX1 INVX1_2 ( .A(_2__3_), .Y(_23_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_24_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_25_) );
NAND3X1 NAND3X1_2 ( .A(_23_), .B(_25_), .C(_24_), .Y(_26_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_20_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_21_) );
OAI21X1 OAI21X1_3 ( .A(_20_), .B(_21_), .C(_2__3_), .Y(_22_) );
NAND2X1 NAND2X1_4 ( .A(_22_), .B(_26_), .Y(_0__7_) );
OAI21X1 OAI21X1_4 ( .A(_23_), .B(_20_), .C(_25_), .Y(_1_) );
INVX1 INVX1_3 ( .A(_2__1_), .Y(_30_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_31_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_32_) );
NAND3X1 NAND3X1_3 ( .A(_30_), .B(_32_), .C(_31_), .Y(_33_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_27_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_28_) );
OAI21X1 OAI21X1_5 ( .A(_27_), .B(_28_), .C(_2__1_), .Y(_29_) );
NAND2X1 NAND2X1_6 ( .A(_29_), .B(_33_), .Y(_0__5_) );
OAI21X1 OAI21X1_6 ( .A(_30_), .B(_27_), .C(_32_), .Y(_2__2_) );
INVX1 INVX1_4 ( .A(_2__2_), .Y(_37_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_38_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_39_) );
NAND3X1 NAND3X1_4 ( .A(_37_), .B(_39_), .C(_38_), .Y(_40_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_34_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_35_) );
OAI21X1 OAI21X1_7 ( .A(_34_), .B(_35_), .C(_2__2_), .Y(_36_) );
NAND2X1 NAND2X1_8 ( .A(_36_), .B(_40_), .Y(_0__6_) );
OAI21X1 OAI21X1_8 ( .A(_37_), .B(_34_), .C(_39_), .Y(_2__3_) );
INVX1 INVX1_5 ( .A(i_add_term2[4]), .Y(_41_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term1[4]), .B(_41_), .Y(_42_) );
INVX1 INVX1_6 ( .A(i_add_term1[4]), .Y(_43_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[4]), .B(_43_), .Y(_44_) );
INVX1 INVX1_7 ( .A(i_add_term1[5]), .Y(_45_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[5]), .B(_45_), .Y(_46_) );
INVX1 INVX1_8 ( .A(i_add_term2[5]), .Y(_47_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term1[5]), .B(_47_), .Y(_48_) );
OAI22X1 OAI22X1_1 ( .A(_42_), .B(_44_), .C(_46_), .D(_48_), .Y(_49_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_50_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_51_) );
NOR2X1 NOR2X1_10 ( .A(_50_), .B(_51_), .Y(_52_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_53_) );
NAND2X1 NAND2X1_9 ( .A(_52_), .B(_53_), .Y(_54_) );
NOR2X1 NOR2X1_11 ( .A(_49_), .B(_54_), .Y(_3_) );
INVX1 INVX1_9 ( .A(_1_), .Y(_55_) );
NAND2X1 NAND2X1_10 ( .A(gnd), .B(_3_), .Y(_56_) );
OAI21X1 OAI21X1_9 ( .A(_3_), .B(_55_), .C(_56_), .Y(w_cout_1_) );
INVX1 INVX1_10 ( .A(w_cout_1_), .Y(_60_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_61_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_62_) );
NAND3X1 NAND3X1_5 ( .A(_60_), .B(_62_), .C(_61_), .Y(_63_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_57_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_58_) );
OAI21X1 OAI21X1_10 ( .A(_57_), .B(_58_), .C(w_cout_1_), .Y(_59_) );
NAND2X1 NAND2X1_12 ( .A(_59_), .B(_63_), .Y(_0__8_) );
OAI21X1 OAI21X1_11 ( .A(_60_), .B(_57_), .C(_62_), .Y(_5__1_) );
INVX1 INVX1_11 ( .A(_5__3_), .Y(_67_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_68_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_69_) );
NAND3X1 NAND3X1_6 ( .A(_67_), .B(_69_), .C(_68_), .Y(_70_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_64_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_65_) );
OAI21X1 OAI21X1_12 ( .A(_64_), .B(_65_), .C(_5__3_), .Y(_66_) );
NAND2X1 NAND2X1_14 ( .A(_66_), .B(_70_), .Y(_0__11_) );
OAI21X1 OAI21X1_13 ( .A(_67_), .B(_64_), .C(_69_), .Y(_4_) );
INVX1 INVX1_12 ( .A(_5__1_), .Y(_74_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_75_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_76_) );
NAND3X1 NAND3X1_7 ( .A(_74_), .B(_76_), .C(_75_), .Y(_77_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_71_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_72_) );
OAI21X1 OAI21X1_14 ( .A(_71_), .B(_72_), .C(_5__1_), .Y(_73_) );
NAND2X1 NAND2X1_16 ( .A(_73_), .B(_77_), .Y(_0__9_) );
OAI21X1 OAI21X1_15 ( .A(_74_), .B(_71_), .C(_76_), .Y(_5__2_) );
INVX1 INVX1_13 ( .A(_5__2_), .Y(_81_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_82_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_83_) );
NAND3X1 NAND3X1_8 ( .A(_81_), .B(_83_), .C(_82_), .Y(_84_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_78_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_79_) );
OAI21X1 OAI21X1_16 ( .A(_78_), .B(_79_), .C(_5__2_), .Y(_80_) );
NAND2X1 NAND2X1_18 ( .A(_80_), .B(_84_), .Y(_0__10_) );
OAI21X1 OAI21X1_17 ( .A(_81_), .B(_78_), .C(_83_), .Y(_5__3_) );
INVX1 INVX1_14 ( .A(i_add_term2[8]), .Y(_85_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term1[8]), .B(_85_), .Y(_86_) );
INVX1 INVX1_15 ( .A(i_add_term1[8]), .Y(_87_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[8]), .B(_87_), .Y(_88_) );
INVX1 INVX1_16 ( .A(i_add_term1[9]), .Y(_89_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[9]), .B(_89_), .Y(_90_) );
INVX1 INVX1_17 ( .A(i_add_term2[9]), .Y(_91_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term1[9]), .B(_91_), .Y(_92_) );
OAI22X1 OAI22X1_2 ( .A(_86_), .B(_88_), .C(_90_), .D(_92_), .Y(_93_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_94_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_95_) );
NOR2X1 NOR2X1_21 ( .A(_94_), .B(_95_), .Y(_96_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_97_) );
NAND2X1 NAND2X1_19 ( .A(_96_), .B(_97_), .Y(_98_) );
NOR2X1 NOR2X1_22 ( .A(_93_), .B(_98_), .Y(_6_) );
INVX1 INVX1_18 ( .A(_4_), .Y(_99_) );
NAND2X1 NAND2X1_20 ( .A(gnd), .B(_6_), .Y(_100_) );
OAI21X1 OAI21X1_18 ( .A(_6_), .B(_99_), .C(_100_), .Y(w_cout_2_) );
INVX1 INVX1_19 ( .A(w_cout_2_), .Y(_104_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_105_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_106_) );
NAND3X1 NAND3X1_9 ( .A(_104_), .B(_106_), .C(_105_), .Y(_107_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_101_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_102_) );
OAI21X1 OAI21X1_19 ( .A(_101_), .B(_102_), .C(w_cout_2_), .Y(_103_) );
NAND2X1 NAND2X1_22 ( .A(_103_), .B(_107_), .Y(_0__12_) );
OAI21X1 OAI21X1_20 ( .A(_104_), .B(_101_), .C(_106_), .Y(_8__1_) );
INVX1 INVX1_20 ( .A(_8__3_), .Y(_111_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_112_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_113_) );
NAND3X1 NAND3X1_10 ( .A(_111_), .B(_113_), .C(_112_), .Y(_114_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_108_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_109_) );
OAI21X1 OAI21X1_21 ( .A(_108_), .B(_109_), .C(_8__3_), .Y(_110_) );
NAND2X1 NAND2X1_24 ( .A(_110_), .B(_114_), .Y(_0__15_) );
OAI21X1 OAI21X1_22 ( .A(_111_), .B(_108_), .C(_113_), .Y(_7_) );
INVX1 INVX1_21 ( .A(_8__1_), .Y(_118_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_119_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_120_) );
NAND3X1 NAND3X1_11 ( .A(_118_), .B(_120_), .C(_119_), .Y(_121_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_115_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_116_) );
OAI21X1 OAI21X1_23 ( .A(_115_), .B(_116_), .C(_8__1_), .Y(_117_) );
NAND2X1 NAND2X1_26 ( .A(_117_), .B(_121_), .Y(_0__13_) );
OAI21X1 OAI21X1_24 ( .A(_118_), .B(_115_), .C(_120_), .Y(_8__2_) );
INVX1 INVX1_22 ( .A(_8__2_), .Y(_125_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_126_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_127_) );
NAND3X1 NAND3X1_12 ( .A(_125_), .B(_127_), .C(_126_), .Y(_128_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_122_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_123_) );
OAI21X1 OAI21X1_25 ( .A(_122_), .B(_123_), .C(_8__2_), .Y(_124_) );
NAND2X1 NAND2X1_28 ( .A(_124_), .B(_128_), .Y(_0__14_) );
OAI21X1 OAI21X1_26 ( .A(_125_), .B(_122_), .C(_127_), .Y(_8__3_) );
INVX1 INVX1_23 ( .A(i_add_term2[12]), .Y(_129_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term1[12]), .B(_129_), .Y(_130_) );
INVX1 INVX1_24 ( .A(i_add_term1[12]), .Y(_131_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[12]), .B(_131_), .Y(_132_) );
INVX1 INVX1_25 ( .A(i_add_term1[13]), .Y(_133_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[13]), .B(_133_), .Y(_134_) );
INVX1 INVX1_26 ( .A(i_add_term2[13]), .Y(_135_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term1[13]), .B(_135_), .Y(_136_) );
OAI22X1 OAI22X1_3 ( .A(_130_), .B(_132_), .C(_134_), .D(_136_), .Y(_137_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_138_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_139_) );
NOR2X1 NOR2X1_32 ( .A(_138_), .B(_139_), .Y(_140_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_141_) );
NAND2X1 NAND2X1_29 ( .A(_140_), .B(_141_), .Y(_142_) );
NOR2X1 NOR2X1_33 ( .A(_137_), .B(_142_), .Y(_9_) );
INVX1 INVX1_27 ( .A(_7_), .Y(_143_) );
NAND2X1 NAND2X1_30 ( .A(gnd), .B(_9_), .Y(_144_) );
OAI21X1 OAI21X1_27 ( .A(_9_), .B(_143_), .C(_144_), .Y(w_cout_3_) );
INVX1 INVX1_28 ( .A(w_cout_3_), .Y(_148_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_149_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_150_) );
NAND3X1 NAND3X1_13 ( .A(_148_), .B(_150_), .C(_149_), .Y(_151_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_145_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_146_) );
OAI21X1 OAI21X1_28 ( .A(_145_), .B(_146_), .C(w_cout_3_), .Y(_147_) );
NAND2X1 NAND2X1_32 ( .A(_147_), .B(_151_), .Y(_0__16_) );
OAI21X1 OAI21X1_29 ( .A(_148_), .B(_145_), .C(_150_), .Y(_11__1_) );
INVX1 INVX1_29 ( .A(_11__3_), .Y(_155_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_156_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_157_) );
NAND3X1 NAND3X1_14 ( .A(_155_), .B(_157_), .C(_156_), .Y(_158_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_152_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_153_) );
OAI21X1 OAI21X1_30 ( .A(_152_), .B(_153_), .C(_11__3_), .Y(_154_) );
NAND2X1 NAND2X1_34 ( .A(_154_), .B(_158_), .Y(_0__19_) );
OAI21X1 OAI21X1_31 ( .A(_155_), .B(_152_), .C(_157_), .Y(_10_) );
INVX1 INVX1_30 ( .A(_11__1_), .Y(_162_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_163_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_164_) );
NAND3X1 NAND3X1_15 ( .A(_162_), .B(_164_), .C(_163_), .Y(_165_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_159_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_160_) );
OAI21X1 OAI21X1_32 ( .A(_159_), .B(_160_), .C(_11__1_), .Y(_161_) );
NAND2X1 NAND2X1_36 ( .A(_161_), .B(_165_), .Y(_0__17_) );
OAI21X1 OAI21X1_33 ( .A(_162_), .B(_159_), .C(_164_), .Y(_11__2_) );
INVX1 INVX1_31 ( .A(_11__2_), .Y(_169_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_170_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_171_) );
NAND3X1 NAND3X1_16 ( .A(_169_), .B(_171_), .C(_170_), .Y(_172_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_166_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_167_) );
OAI21X1 OAI21X1_34 ( .A(_166_), .B(_167_), .C(_11__2_), .Y(_168_) );
NAND2X1 NAND2X1_38 ( .A(_168_), .B(_172_), .Y(_0__18_) );
OAI21X1 OAI21X1_35 ( .A(_169_), .B(_166_), .C(_171_), .Y(_11__3_) );
INVX1 INVX1_32 ( .A(i_add_term2[16]), .Y(_173_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term1[16]), .B(_173_), .Y(_174_) );
INVX1 INVX1_33 ( .A(i_add_term1[16]), .Y(_175_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[16]), .B(_175_), .Y(_176_) );
INVX1 INVX1_34 ( .A(i_add_term1[17]), .Y(_177_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[17]), .B(_177_), .Y(_178_) );
INVX1 INVX1_35 ( .A(i_add_term2[17]), .Y(_179_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term1[17]), .B(_179_), .Y(_180_) );
OAI22X1 OAI22X1_4 ( .A(_174_), .B(_176_), .C(_178_), .D(_180_), .Y(_181_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_182_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_183_) );
NOR2X1 NOR2X1_43 ( .A(_182_), .B(_183_), .Y(_184_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_185_) );
NAND2X1 NAND2X1_39 ( .A(_184_), .B(_185_), .Y(_186_) );
NOR2X1 NOR2X1_44 ( .A(_181_), .B(_186_), .Y(_12_) );
INVX1 INVX1_36 ( .A(_10_), .Y(_187_) );
NAND2X1 NAND2X1_40 ( .A(gnd), .B(_12_), .Y(_188_) );
OAI21X1 OAI21X1_36 ( .A(_12_), .B(_187_), .C(_188_), .Y(w_cout_4_) );
INVX1 INVX1_37 ( .A(gnd), .Y(_192_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_193_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_194_) );
NAND3X1 NAND3X1_17 ( .A(_192_), .B(_194_), .C(_193_), .Y(_195_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_189_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_190_) );
OAI21X1 OAI21X1_37 ( .A(_189_), .B(_190_), .C(gnd), .Y(_191_) );
NAND2X1 NAND2X1_42 ( .A(_191_), .B(_195_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_38 ( .A(_192_), .B(_189_), .C(_194_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_38 ( .A(rca_inst_fa3_i_carry), .Y(_199_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_200_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_201_) );
NAND3X1 NAND3X1_18 ( .A(_199_), .B(_201_), .C(_200_), .Y(_202_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_196_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_197_) );
OAI21X1 OAI21X1_39 ( .A(_196_), .B(_197_), .C(rca_inst_fa3_i_carry), .Y(_198_) );
NAND2X1 NAND2X1_44 ( .A(_198_), .B(_202_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_40 ( .A(_199_), .B(_196_), .C(_201_), .Y(cout0) );
INVX1 INVX1_39 ( .A(rca_inst_fa0_o_carry), .Y(_206_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_207_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_208_) );
NAND3X1 NAND3X1_19 ( .A(_206_), .B(_208_), .C(_207_), .Y(_209_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_203_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_204_) );
OAI21X1 OAI21X1_41 ( .A(_203_), .B(_204_), .C(rca_inst_fa0_o_carry), .Y(_205_) );
NAND2X1 NAND2X1_46 ( .A(_205_), .B(_209_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_42 ( .A(_206_), .B(_203_), .C(_208_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_40 ( .A(rca_inst_fa_1__o_carry), .Y(_213_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_214_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_215_) );
NAND3X1 NAND3X1_20 ( .A(_213_), .B(_215_), .C(_214_), .Y(_216_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_210_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_211_) );
OAI21X1 OAI21X1_43 ( .A(_210_), .B(_211_), .C(rca_inst_fa_1__o_carry), .Y(_212_) );
NAND2X1 NAND2X1_48 ( .A(_212_), .B(_216_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_44 ( .A(_213_), .B(_210_), .C(_215_), .Y(rca_inst_fa3_i_carry) );
INVX1 INVX1_41 ( .A(i_add_term2[0]), .Y(_217_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term1[0]), .B(_217_), .Y(_218_) );
INVX1 INVX1_42 ( .A(i_add_term1[0]), .Y(_219_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[0]), .B(_219_), .Y(_220_) );
INVX1 INVX1_43 ( .A(i_add_term1[1]), .Y(_221_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[1]), .B(_221_), .Y(_222_) );
INVX1 INVX1_44 ( .A(i_add_term2[1]), .Y(_223_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term1[1]), .B(_223_), .Y(_224_) );
OAI22X1 OAI22X1_5 ( .A(_218_), .B(_220_), .C(_222_), .D(_224_), .Y(_225_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_226_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_227_) );
NOR2X1 NOR2X1_54 ( .A(_226_), .B(_227_), .Y(_228_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_229_) );
NAND2X1 NAND2X1_49 ( .A(_228_), .B(_229_), .Y(_230_) );
NOR2X1 NOR2X1_55 ( .A(_225_), .B(_230_), .Y(skip0_P) );
INVX1 INVX1_45 ( .A(cout0), .Y(_231_) );
NAND2X1 NAND2X1_50 ( .A(gnd), .B(skip0_P), .Y(_232_) );
OAI21X1 OAI21X1_45 ( .A(skip0_P), .B(_231_), .C(_232_), .Y(skip0_cin_next) );
BUFX2 BUFX2_22 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_23 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_24 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_25 ( .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_26 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
