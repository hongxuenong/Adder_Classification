module csa_41bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output cout;

OAI21X1 OAI21X1_1 ( .A(_220_), .B(_217_), .C(_222_), .Y(_11__1_) );
INVX1 INVX1_1 ( .A(_11__1_), .Y(_227_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_228_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_229_) );
NAND3X1 NAND3X1_1 ( .A(_227_), .B(_229_), .C(_228_), .Y(_230_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_224_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_225_) );
OAI21X1 OAI21X1_2 ( .A(_224_), .B(_225_), .C(_11__1_), .Y(_226_) );
NAND2X1 NAND2X1_2 ( .A(_226_), .B(_230_), .Y(_9__1_) );
OAI21X1 OAI21X1_3 ( .A(_227_), .B(_224_), .C(_229_), .Y(_11__2_) );
INVX1 INVX1_2 ( .A(_11__2_), .Y(_234_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_235_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_236_) );
NAND3X1 NAND3X1_2 ( .A(_234_), .B(_236_), .C(_235_), .Y(_237_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_231_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_232_) );
OAI21X1 OAI21X1_4 ( .A(_231_), .B(_232_), .C(_11__2_), .Y(_233_) );
NAND2X1 NAND2X1_4 ( .A(_233_), .B(_237_), .Y(_9__2_) );
OAI21X1 OAI21X1_5 ( .A(_234_), .B(_231_), .C(_236_), .Y(_11__3_) );
INVX1 INVX1_3 ( .A(_11__3_), .Y(_241_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_242_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_243_) );
NAND3X1 NAND3X1_3 ( .A(_241_), .B(_243_), .C(_242_), .Y(_244_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_238_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_239_) );
OAI21X1 OAI21X1_6 ( .A(_238_), .B(_239_), .C(_11__3_), .Y(_240_) );
NAND2X1 NAND2X1_6 ( .A(_240_), .B(_244_), .Y(_9__3_) );
OAI21X1 OAI21X1_7 ( .A(_241_), .B(_238_), .C(_243_), .Y(_7_) );
INVX1 INVX1_4 ( .A(1'b1), .Y(_248_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_249_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_250_) );
NAND3X1 NAND3X1_4 ( .A(_248_), .B(_250_), .C(_249_), .Y(_251_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_245_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_246_) );
OAI21X1 OAI21X1_8 ( .A(_245_), .B(_246_), .C(1'b1), .Y(_247_) );
NAND2X1 NAND2X1_8 ( .A(_247_), .B(_251_), .Y(_10__0_) );
OAI21X1 OAI21X1_9 ( .A(_248_), .B(_245_), .C(_250_), .Y(_12__1_) );
INVX1 INVX1_5 ( .A(_12__1_), .Y(_255_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_256_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_257_) );
NAND3X1 NAND3X1_5 ( .A(_255_), .B(_257_), .C(_256_), .Y(_258_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_252_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_253_) );
OAI21X1 OAI21X1_10 ( .A(_252_), .B(_253_), .C(_12__1_), .Y(_254_) );
NAND2X1 NAND2X1_10 ( .A(_254_), .B(_258_), .Y(_10__1_) );
OAI21X1 OAI21X1_11 ( .A(_255_), .B(_252_), .C(_257_), .Y(_12__2_) );
INVX1 INVX1_6 ( .A(_12__2_), .Y(_262_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_263_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_264_) );
NAND3X1 NAND3X1_6 ( .A(_262_), .B(_264_), .C(_263_), .Y(_265_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_259_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_260_) );
OAI21X1 OAI21X1_12 ( .A(_259_), .B(_260_), .C(_12__2_), .Y(_261_) );
NAND2X1 NAND2X1_12 ( .A(_261_), .B(_265_), .Y(_10__2_) );
OAI21X1 OAI21X1_13 ( .A(_262_), .B(_259_), .C(_264_), .Y(_12__3_) );
INVX1 INVX1_7 ( .A(_12__3_), .Y(_269_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_270_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_271_) );
NAND3X1 NAND3X1_7 ( .A(_269_), .B(_271_), .C(_270_), .Y(_272_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_266_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_267_) );
OAI21X1 OAI21X1_14 ( .A(_266_), .B(_267_), .C(_12__3_), .Y(_268_) );
NAND2X1 NAND2X1_14 ( .A(_268_), .B(_272_), .Y(_10__3_) );
OAI21X1 OAI21X1_15 ( .A(_269_), .B(_266_), .C(_271_), .Y(_8_) );
INVX1 INVX1_8 ( .A(1'b0), .Y(_276_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_277_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_278_) );
NAND3X1 NAND3X1_8 ( .A(_276_), .B(_278_), .C(_277_), .Y(_279_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_273_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_274_) );
OAI21X1 OAI21X1_16 ( .A(_273_), .B(_274_), .C(1'b0), .Y(_275_) );
NAND2X1 NAND2X1_16 ( .A(_275_), .B(_279_), .Y(_15__0_) );
OAI21X1 OAI21X1_17 ( .A(_276_), .B(_273_), .C(_278_), .Y(_17__1_) );
INVX1 INVX1_9 ( .A(_17__1_), .Y(_283_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_284_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_285_) );
NAND3X1 NAND3X1_9 ( .A(_283_), .B(_285_), .C(_284_), .Y(_286_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_280_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_281_) );
OAI21X1 OAI21X1_18 ( .A(_280_), .B(_281_), .C(_17__1_), .Y(_282_) );
NAND2X1 NAND2X1_18 ( .A(_282_), .B(_286_), .Y(_15__1_) );
OAI21X1 OAI21X1_19 ( .A(_283_), .B(_280_), .C(_285_), .Y(_17__2_) );
INVX1 INVX1_10 ( .A(_17__2_), .Y(_290_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_291_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_292_) );
NAND3X1 NAND3X1_10 ( .A(_290_), .B(_292_), .C(_291_), .Y(_293_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_287_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_288_) );
OAI21X1 OAI21X1_20 ( .A(_287_), .B(_288_), .C(_17__2_), .Y(_289_) );
NAND2X1 NAND2X1_20 ( .A(_289_), .B(_293_), .Y(_15__2_) );
OAI21X1 OAI21X1_21 ( .A(_290_), .B(_287_), .C(_292_), .Y(_17__3_) );
INVX1 INVX1_11 ( .A(_17__3_), .Y(_297_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_298_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_299_) );
NAND3X1 NAND3X1_11 ( .A(_297_), .B(_299_), .C(_298_), .Y(_300_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_294_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_295_) );
OAI21X1 OAI21X1_22 ( .A(_294_), .B(_295_), .C(_17__3_), .Y(_296_) );
NAND2X1 NAND2X1_22 ( .A(_296_), .B(_300_), .Y(_15__3_) );
OAI21X1 OAI21X1_23 ( .A(_297_), .B(_294_), .C(_299_), .Y(_13_) );
INVX1 INVX1_12 ( .A(1'b1), .Y(_304_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_305_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_306_) );
NAND3X1 NAND3X1_12 ( .A(_304_), .B(_306_), .C(_305_), .Y(_307_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_301_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_302_) );
OAI21X1 OAI21X1_24 ( .A(_301_), .B(_302_), .C(1'b1), .Y(_303_) );
NAND2X1 NAND2X1_24 ( .A(_303_), .B(_307_), .Y(_16__0_) );
OAI21X1 OAI21X1_25 ( .A(_304_), .B(_301_), .C(_306_), .Y(_18__1_) );
INVX1 INVX1_13 ( .A(_18__1_), .Y(_311_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_312_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_313_) );
NAND3X1 NAND3X1_13 ( .A(_311_), .B(_313_), .C(_312_), .Y(_314_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_308_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_309_) );
OAI21X1 OAI21X1_26 ( .A(_308_), .B(_309_), .C(_18__1_), .Y(_310_) );
NAND2X1 NAND2X1_26 ( .A(_310_), .B(_314_), .Y(_16__1_) );
OAI21X1 OAI21X1_27 ( .A(_311_), .B(_308_), .C(_313_), .Y(_18__2_) );
INVX1 INVX1_14 ( .A(_18__2_), .Y(_318_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_319_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_320_) );
NAND3X1 NAND3X1_14 ( .A(_318_), .B(_320_), .C(_319_), .Y(_321_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_315_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_316_) );
OAI21X1 OAI21X1_28 ( .A(_315_), .B(_316_), .C(_18__2_), .Y(_317_) );
NAND2X1 NAND2X1_28 ( .A(_317_), .B(_321_), .Y(_16__2_) );
OAI21X1 OAI21X1_29 ( .A(_318_), .B(_315_), .C(_320_), .Y(_18__3_) );
INVX1 INVX1_15 ( .A(_18__3_), .Y(_325_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_326_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_327_) );
NAND3X1 NAND3X1_15 ( .A(_325_), .B(_327_), .C(_326_), .Y(_328_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_322_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_323_) );
OAI21X1 OAI21X1_30 ( .A(_322_), .B(_323_), .C(_18__3_), .Y(_324_) );
NAND2X1 NAND2X1_30 ( .A(_324_), .B(_328_), .Y(_16__3_) );
OAI21X1 OAI21X1_31 ( .A(_325_), .B(_322_), .C(_327_), .Y(_14_) );
INVX1 INVX1_16 ( .A(1'b0), .Y(_332_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_333_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_334_) );
NAND3X1 NAND3X1_16 ( .A(_332_), .B(_334_), .C(_333_), .Y(_335_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_329_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_330_) );
OAI21X1 OAI21X1_32 ( .A(_329_), .B(_330_), .C(1'b0), .Y(_331_) );
NAND2X1 NAND2X1_32 ( .A(_331_), .B(_335_), .Y(_21__0_) );
OAI21X1 OAI21X1_33 ( .A(_332_), .B(_329_), .C(_334_), .Y(_23__1_) );
INVX1 INVX1_17 ( .A(_23__1_), .Y(_339_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_340_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_341_) );
NAND3X1 NAND3X1_17 ( .A(_339_), .B(_341_), .C(_340_), .Y(_342_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_336_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_337_) );
OAI21X1 OAI21X1_34 ( .A(_336_), .B(_337_), .C(_23__1_), .Y(_338_) );
NAND2X1 NAND2X1_34 ( .A(_338_), .B(_342_), .Y(_21__1_) );
OAI21X1 OAI21X1_35 ( .A(_339_), .B(_336_), .C(_341_), .Y(_23__2_) );
INVX1 INVX1_18 ( .A(_23__2_), .Y(_346_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_347_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_348_) );
NAND3X1 NAND3X1_18 ( .A(_346_), .B(_348_), .C(_347_), .Y(_349_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_343_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_344_) );
OAI21X1 OAI21X1_36 ( .A(_343_), .B(_344_), .C(_23__2_), .Y(_345_) );
NAND2X1 NAND2X1_36 ( .A(_345_), .B(_349_), .Y(_21__2_) );
OAI21X1 OAI21X1_37 ( .A(_346_), .B(_343_), .C(_348_), .Y(_23__3_) );
INVX1 INVX1_19 ( .A(_23__3_), .Y(_353_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_354_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_355_) );
NAND3X1 NAND3X1_19 ( .A(_353_), .B(_355_), .C(_354_), .Y(_356_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_350_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_351_) );
OAI21X1 OAI21X1_38 ( .A(_350_), .B(_351_), .C(_23__3_), .Y(_352_) );
NAND2X1 NAND2X1_38 ( .A(_352_), .B(_356_), .Y(_21__3_) );
OAI21X1 OAI21X1_39 ( .A(_353_), .B(_350_), .C(_355_), .Y(_19_) );
INVX1 INVX1_20 ( .A(1'b1), .Y(_360_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_361_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_362_) );
NAND3X1 NAND3X1_20 ( .A(_360_), .B(_362_), .C(_361_), .Y(_363_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_357_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_358_) );
OAI21X1 OAI21X1_40 ( .A(_357_), .B(_358_), .C(1'b1), .Y(_359_) );
NAND2X1 NAND2X1_40 ( .A(_359_), .B(_363_), .Y(_22__0_) );
OAI21X1 OAI21X1_41 ( .A(_360_), .B(_357_), .C(_362_), .Y(_24__1_) );
INVX1 INVX1_21 ( .A(_24__1_), .Y(_367_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_368_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_369_) );
NAND3X1 NAND3X1_21 ( .A(_367_), .B(_369_), .C(_368_), .Y(_370_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_364_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_365_) );
OAI21X1 OAI21X1_42 ( .A(_364_), .B(_365_), .C(_24__1_), .Y(_366_) );
NAND2X1 NAND2X1_42 ( .A(_366_), .B(_370_), .Y(_22__1_) );
OAI21X1 OAI21X1_43 ( .A(_367_), .B(_364_), .C(_369_), .Y(_24__2_) );
INVX1 INVX1_22 ( .A(_24__2_), .Y(_374_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_375_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_376_) );
NAND3X1 NAND3X1_22 ( .A(_374_), .B(_376_), .C(_375_), .Y(_377_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_371_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_372_) );
OAI21X1 OAI21X1_44 ( .A(_371_), .B(_372_), .C(_24__2_), .Y(_373_) );
NAND2X1 NAND2X1_44 ( .A(_373_), .B(_377_), .Y(_22__2_) );
OAI21X1 OAI21X1_45 ( .A(_374_), .B(_371_), .C(_376_), .Y(_24__3_) );
INVX1 INVX1_23 ( .A(_24__3_), .Y(_381_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_382_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_383_) );
NAND3X1 NAND3X1_23 ( .A(_381_), .B(_383_), .C(_382_), .Y(_384_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_378_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_379_) );
OAI21X1 OAI21X1_46 ( .A(_378_), .B(_379_), .C(_24__3_), .Y(_380_) );
NAND2X1 NAND2X1_46 ( .A(_380_), .B(_384_), .Y(_22__3_) );
OAI21X1 OAI21X1_47 ( .A(_381_), .B(_378_), .C(_383_), .Y(_20_) );
INVX1 INVX1_24 ( .A(1'b0), .Y(_388_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_389_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_390_) );
NAND3X1 NAND3X1_24 ( .A(_388_), .B(_390_), .C(_389_), .Y(_391_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_385_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_386_) );
OAI21X1 OAI21X1_48 ( .A(_385_), .B(_386_), .C(1'b0), .Y(_387_) );
NAND2X1 NAND2X1_48 ( .A(_387_), .B(_391_), .Y(_27__0_) );
OAI21X1 OAI21X1_49 ( .A(_388_), .B(_385_), .C(_390_), .Y(_29__1_) );
INVX1 INVX1_25 ( .A(_29__1_), .Y(_395_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_396_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_397_) );
NAND3X1 NAND3X1_25 ( .A(_395_), .B(_397_), .C(_396_), .Y(_398_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_392_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_393_) );
OAI21X1 OAI21X1_50 ( .A(_392_), .B(_393_), .C(_29__1_), .Y(_394_) );
NAND2X1 NAND2X1_50 ( .A(_394_), .B(_398_), .Y(_27__1_) );
OAI21X1 OAI21X1_51 ( .A(_395_), .B(_392_), .C(_397_), .Y(_29__2_) );
INVX1 INVX1_26 ( .A(_29__2_), .Y(_402_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_403_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_404_) );
NAND3X1 NAND3X1_26 ( .A(_402_), .B(_404_), .C(_403_), .Y(_405_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_399_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_400_) );
OAI21X1 OAI21X1_52 ( .A(_399_), .B(_400_), .C(_29__2_), .Y(_401_) );
NAND2X1 NAND2X1_52 ( .A(_401_), .B(_405_), .Y(_27__2_) );
OAI21X1 OAI21X1_53 ( .A(_402_), .B(_399_), .C(_404_), .Y(_29__3_) );
INVX1 INVX1_27 ( .A(_29__3_), .Y(_409_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_410_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_411_) );
NAND3X1 NAND3X1_27 ( .A(_409_), .B(_411_), .C(_410_), .Y(_412_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_406_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_407_) );
OAI21X1 OAI21X1_54 ( .A(_406_), .B(_407_), .C(_29__3_), .Y(_408_) );
NAND2X1 NAND2X1_54 ( .A(_408_), .B(_412_), .Y(_27__3_) );
OAI21X1 OAI21X1_55 ( .A(_409_), .B(_406_), .C(_411_), .Y(_25_) );
INVX1 INVX1_28 ( .A(1'b1), .Y(_416_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_417_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_418_) );
NAND3X1 NAND3X1_28 ( .A(_416_), .B(_418_), .C(_417_), .Y(_419_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_413_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_414_) );
OAI21X1 OAI21X1_56 ( .A(_413_), .B(_414_), .C(1'b1), .Y(_415_) );
NAND2X1 NAND2X1_56 ( .A(_415_), .B(_419_), .Y(_28__0_) );
OAI21X1 OAI21X1_57 ( .A(_416_), .B(_413_), .C(_418_), .Y(_30__1_) );
INVX1 INVX1_29 ( .A(_30__1_), .Y(_423_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_424_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_425_) );
NAND3X1 NAND3X1_29 ( .A(_423_), .B(_425_), .C(_424_), .Y(_426_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_420_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_421_) );
OAI21X1 OAI21X1_58 ( .A(_420_), .B(_421_), .C(_30__1_), .Y(_422_) );
NAND2X1 NAND2X1_58 ( .A(_422_), .B(_426_), .Y(_28__1_) );
OAI21X1 OAI21X1_59 ( .A(_423_), .B(_420_), .C(_425_), .Y(_30__2_) );
INVX1 INVX1_30 ( .A(_30__2_), .Y(_430_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_431_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_432_) );
NAND3X1 NAND3X1_30 ( .A(_430_), .B(_432_), .C(_431_), .Y(_433_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_427_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_428_) );
OAI21X1 OAI21X1_60 ( .A(_427_), .B(_428_), .C(_30__2_), .Y(_429_) );
NAND2X1 NAND2X1_60 ( .A(_429_), .B(_433_), .Y(_28__2_) );
OAI21X1 OAI21X1_61 ( .A(_430_), .B(_427_), .C(_432_), .Y(_30__3_) );
INVX1 INVX1_31 ( .A(_30__3_), .Y(_437_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_438_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_439_) );
NAND3X1 NAND3X1_31 ( .A(_437_), .B(_439_), .C(_438_), .Y(_440_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_434_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_435_) );
OAI21X1 OAI21X1_62 ( .A(_434_), .B(_435_), .C(_30__3_), .Y(_436_) );
NAND2X1 NAND2X1_62 ( .A(_436_), .B(_440_), .Y(_28__3_) );
OAI21X1 OAI21X1_63 ( .A(_437_), .B(_434_), .C(_439_), .Y(_26_) );
INVX1 INVX1_32 ( .A(1'b0), .Y(_444_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_445_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_446_) );
NAND3X1 NAND3X1_32 ( .A(_444_), .B(_446_), .C(_445_), .Y(_447_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_441_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_442_) );
OAI21X1 OAI21X1_64 ( .A(_441_), .B(_442_), .C(1'b0), .Y(_443_) );
NAND2X1 NAND2X1_64 ( .A(_443_), .B(_447_), .Y(_33__0_) );
OAI21X1 OAI21X1_65 ( .A(_444_), .B(_441_), .C(_446_), .Y(_35__1_) );
INVX1 INVX1_33 ( .A(_35__1_), .Y(_451_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_452_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_453_) );
NAND3X1 NAND3X1_33 ( .A(_451_), .B(_453_), .C(_452_), .Y(_454_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_448_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_449_) );
OAI21X1 OAI21X1_66 ( .A(_448_), .B(_449_), .C(_35__1_), .Y(_450_) );
NAND2X1 NAND2X1_66 ( .A(_450_), .B(_454_), .Y(_33__1_) );
OAI21X1 OAI21X1_67 ( .A(_451_), .B(_448_), .C(_453_), .Y(_35__2_) );
INVX1 INVX1_34 ( .A(_35__2_), .Y(_458_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_459_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_460_) );
NAND3X1 NAND3X1_34 ( .A(_458_), .B(_460_), .C(_459_), .Y(_461_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_455_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_456_) );
OAI21X1 OAI21X1_68 ( .A(_455_), .B(_456_), .C(_35__2_), .Y(_457_) );
NAND2X1 NAND2X1_68 ( .A(_457_), .B(_461_), .Y(_33__2_) );
OAI21X1 OAI21X1_69 ( .A(_458_), .B(_455_), .C(_460_), .Y(_35__3_) );
INVX1 INVX1_35 ( .A(_35__3_), .Y(_465_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_466_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_467_) );
NAND3X1 NAND3X1_35 ( .A(_465_), .B(_467_), .C(_466_), .Y(_468_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_462_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_463_) );
OAI21X1 OAI21X1_70 ( .A(_462_), .B(_463_), .C(_35__3_), .Y(_464_) );
NAND2X1 NAND2X1_70 ( .A(_464_), .B(_468_), .Y(_33__3_) );
OAI21X1 OAI21X1_71 ( .A(_465_), .B(_462_), .C(_467_), .Y(_31_) );
INVX1 INVX1_36 ( .A(1'b1), .Y(_472_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_473_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_474_) );
NAND3X1 NAND3X1_36 ( .A(_472_), .B(_474_), .C(_473_), .Y(_475_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_469_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_470_) );
OAI21X1 OAI21X1_72 ( .A(_469_), .B(_470_), .C(1'b1), .Y(_471_) );
NAND2X1 NAND2X1_72 ( .A(_471_), .B(_475_), .Y(_34__0_) );
OAI21X1 OAI21X1_73 ( .A(_472_), .B(_469_), .C(_474_), .Y(_36__1_) );
INVX1 INVX1_37 ( .A(_36__1_), .Y(_479_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_480_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_481_) );
NAND3X1 NAND3X1_37 ( .A(_479_), .B(_481_), .C(_480_), .Y(_482_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_476_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_477_) );
OAI21X1 OAI21X1_74 ( .A(_476_), .B(_477_), .C(_36__1_), .Y(_478_) );
NAND2X1 NAND2X1_74 ( .A(_478_), .B(_482_), .Y(_34__1_) );
OAI21X1 OAI21X1_75 ( .A(_479_), .B(_476_), .C(_481_), .Y(_36__2_) );
INVX1 INVX1_38 ( .A(_36__2_), .Y(_486_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_487_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_488_) );
NAND3X1 NAND3X1_38 ( .A(_486_), .B(_488_), .C(_487_), .Y(_489_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_483_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_484_) );
OAI21X1 OAI21X1_76 ( .A(_483_), .B(_484_), .C(_36__2_), .Y(_485_) );
NAND2X1 NAND2X1_76 ( .A(_485_), .B(_489_), .Y(_34__2_) );
OAI21X1 OAI21X1_77 ( .A(_486_), .B(_483_), .C(_488_), .Y(_36__3_) );
INVX1 INVX1_39 ( .A(_36__3_), .Y(_493_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_494_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_495_) );
NAND3X1 NAND3X1_39 ( .A(_493_), .B(_495_), .C(_494_), .Y(_496_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_490_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_491_) );
OAI21X1 OAI21X1_78 ( .A(_490_), .B(_491_), .C(_36__3_), .Y(_492_) );
NAND2X1 NAND2X1_78 ( .A(_492_), .B(_496_), .Y(_34__3_) );
OAI21X1 OAI21X1_79 ( .A(_493_), .B(_490_), .C(_495_), .Y(_32_) );
INVX1 INVX1_40 ( .A(1'b0), .Y(_500_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_501_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_502_) );
NAND3X1 NAND3X1_40 ( .A(_500_), .B(_502_), .C(_501_), .Y(_503_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_497_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_498_) );
OAI21X1 OAI21X1_80 ( .A(_497_), .B(_498_), .C(1'b0), .Y(_499_) );
NAND2X1 NAND2X1_80 ( .A(_499_), .B(_503_), .Y(_39__0_) );
OAI21X1 OAI21X1_81 ( .A(_500_), .B(_497_), .C(_502_), .Y(_41__1_) );
INVX1 INVX1_41 ( .A(_41__1_), .Y(_507_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_508_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_509_) );
NAND3X1 NAND3X1_41 ( .A(_507_), .B(_509_), .C(_508_), .Y(_510_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_504_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_505_) );
OAI21X1 OAI21X1_82 ( .A(_504_), .B(_505_), .C(_41__1_), .Y(_506_) );
NAND2X1 NAND2X1_82 ( .A(_506_), .B(_510_), .Y(_39__1_) );
OAI21X1 OAI21X1_83 ( .A(_507_), .B(_504_), .C(_509_), .Y(_41__2_) );
INVX1 INVX1_42 ( .A(_41__2_), .Y(_514_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_515_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_516_) );
NAND3X1 NAND3X1_42 ( .A(_514_), .B(_516_), .C(_515_), .Y(_517_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_511_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_512_) );
OAI21X1 OAI21X1_84 ( .A(_511_), .B(_512_), .C(_41__2_), .Y(_513_) );
NAND2X1 NAND2X1_84 ( .A(_513_), .B(_517_), .Y(_39__2_) );
OAI21X1 OAI21X1_85 ( .A(_514_), .B(_511_), .C(_516_), .Y(_41__3_) );
INVX1 INVX1_43 ( .A(_41__3_), .Y(_521_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_522_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_523_) );
NAND3X1 NAND3X1_43 ( .A(_521_), .B(_523_), .C(_522_), .Y(_524_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_518_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_519_) );
OAI21X1 OAI21X1_86 ( .A(_518_), .B(_519_), .C(_41__3_), .Y(_520_) );
NAND2X1 NAND2X1_86 ( .A(_520_), .B(_524_), .Y(_39__3_) );
OAI21X1 OAI21X1_87 ( .A(_521_), .B(_518_), .C(_523_), .Y(_37_) );
INVX1 INVX1_44 ( .A(1'b1), .Y(_528_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_529_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_530_) );
NAND3X1 NAND3X1_44 ( .A(_528_), .B(_530_), .C(_529_), .Y(_531_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_525_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_526_) );
OAI21X1 OAI21X1_88 ( .A(_525_), .B(_526_), .C(1'b1), .Y(_527_) );
NAND2X1 NAND2X1_88 ( .A(_527_), .B(_531_), .Y(_40__0_) );
OAI21X1 OAI21X1_89 ( .A(_528_), .B(_525_), .C(_530_), .Y(_42__1_) );
INVX1 INVX1_45 ( .A(_42__1_), .Y(_535_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_536_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_537_) );
NAND3X1 NAND3X1_45 ( .A(_535_), .B(_537_), .C(_536_), .Y(_538_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_532_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_533_) );
OAI21X1 OAI21X1_90 ( .A(_532_), .B(_533_), .C(_42__1_), .Y(_534_) );
NAND2X1 NAND2X1_90 ( .A(_534_), .B(_538_), .Y(_40__1_) );
OAI21X1 OAI21X1_91 ( .A(_535_), .B(_532_), .C(_537_), .Y(_42__2_) );
INVX1 INVX1_46 ( .A(_42__2_), .Y(_542_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_543_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_544_) );
NAND3X1 NAND3X1_46 ( .A(_542_), .B(_544_), .C(_543_), .Y(_545_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_539_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_540_) );
OAI21X1 OAI21X1_92 ( .A(_539_), .B(_540_), .C(_42__2_), .Y(_541_) );
NAND2X1 NAND2X1_92 ( .A(_541_), .B(_545_), .Y(_40__2_) );
OAI21X1 OAI21X1_93 ( .A(_542_), .B(_539_), .C(_544_), .Y(_42__3_) );
INVX1 INVX1_47 ( .A(_42__3_), .Y(_549_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_550_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_551_) );
NAND3X1 NAND3X1_47 ( .A(_549_), .B(_551_), .C(_550_), .Y(_552_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_546_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_547_) );
OAI21X1 OAI21X1_94 ( .A(_546_), .B(_547_), .C(_42__3_), .Y(_548_) );
NAND2X1 NAND2X1_94 ( .A(_548_), .B(_552_), .Y(_40__3_) );
OAI21X1 OAI21X1_95 ( .A(_549_), .B(_546_), .C(_551_), .Y(_38_) );
INVX1 INVX1_48 ( .A(1'b0), .Y(_556_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_557_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_558_) );
NAND3X1 NAND3X1_48 ( .A(_556_), .B(_558_), .C(_557_), .Y(_559_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_553_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_554_) );
OAI21X1 OAI21X1_96 ( .A(_553_), .B(_554_), .C(1'b0), .Y(_555_) );
NAND2X1 NAND2X1_96 ( .A(_555_), .B(_559_), .Y(_45__0_) );
OAI21X1 OAI21X1_97 ( .A(_556_), .B(_553_), .C(_558_), .Y(_47__1_) );
INVX1 INVX1_49 ( .A(_47__1_), .Y(_563_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_564_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_565_) );
NAND3X1 NAND3X1_49 ( .A(_563_), .B(_565_), .C(_564_), .Y(_566_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_560_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_561_) );
OAI21X1 OAI21X1_98 ( .A(_560_), .B(_561_), .C(_47__1_), .Y(_562_) );
NAND2X1 NAND2X1_98 ( .A(_562_), .B(_566_), .Y(_45__1_) );
OAI21X1 OAI21X1_99 ( .A(_563_), .B(_560_), .C(_565_), .Y(_47__2_) );
INVX1 INVX1_50 ( .A(_47__2_), .Y(_570_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_571_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_572_) );
NAND3X1 NAND3X1_50 ( .A(_570_), .B(_572_), .C(_571_), .Y(_573_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_567_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_568_) );
OAI21X1 OAI21X1_100 ( .A(_567_), .B(_568_), .C(_47__2_), .Y(_569_) );
NAND2X1 NAND2X1_100 ( .A(_569_), .B(_573_), .Y(_45__2_) );
OAI21X1 OAI21X1_101 ( .A(_570_), .B(_567_), .C(_572_), .Y(_47__3_) );
INVX1 INVX1_51 ( .A(_47__3_), .Y(_577_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_578_) );
NAND2X1 NAND2X1_101 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_579_) );
NAND3X1 NAND3X1_51 ( .A(_577_), .B(_579_), .C(_578_), .Y(_580_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_574_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_575_) );
OAI21X1 OAI21X1_102 ( .A(_574_), .B(_575_), .C(_47__3_), .Y(_576_) );
NAND2X1 NAND2X1_102 ( .A(_576_), .B(_580_), .Y(_45__3_) );
OAI21X1 OAI21X1_103 ( .A(_577_), .B(_574_), .C(_579_), .Y(_43_) );
INVX1 INVX1_52 ( .A(1'b1), .Y(_584_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_585_) );
NAND2X1 NAND2X1_103 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_586_) );
NAND3X1 NAND3X1_52 ( .A(_584_), .B(_586_), .C(_585_), .Y(_587_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_581_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_582_) );
OAI21X1 OAI21X1_104 ( .A(_581_), .B(_582_), .C(1'b1), .Y(_583_) );
NAND2X1 NAND2X1_104 ( .A(_583_), .B(_587_), .Y(_46__0_) );
OAI21X1 OAI21X1_105 ( .A(_584_), .B(_581_), .C(_586_), .Y(_48__1_) );
INVX1 INVX1_53 ( .A(_48__1_), .Y(_591_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_592_) );
NAND2X1 NAND2X1_105 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_593_) );
NAND3X1 NAND3X1_53 ( .A(_591_), .B(_593_), .C(_592_), .Y(_594_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_588_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_589_) );
OAI21X1 OAI21X1_106 ( .A(_588_), .B(_589_), .C(_48__1_), .Y(_590_) );
NAND2X1 NAND2X1_106 ( .A(_590_), .B(_594_), .Y(_46__1_) );
OAI21X1 OAI21X1_107 ( .A(_591_), .B(_588_), .C(_593_), .Y(_48__2_) );
INVX1 INVX1_54 ( .A(_48__2_), .Y(_598_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_599_) );
NAND2X1 NAND2X1_107 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_600_) );
NAND3X1 NAND3X1_54 ( .A(_598_), .B(_600_), .C(_599_), .Y(_601_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_595_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_596_) );
OAI21X1 OAI21X1_108 ( .A(_595_), .B(_596_), .C(_48__2_), .Y(_597_) );
NAND2X1 NAND2X1_108 ( .A(_597_), .B(_601_), .Y(_46__2_) );
OAI21X1 OAI21X1_109 ( .A(_598_), .B(_595_), .C(_600_), .Y(_48__3_) );
INVX1 INVX1_55 ( .A(_48__3_), .Y(_605_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_606_) );
NAND2X1 NAND2X1_109 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_607_) );
NAND3X1 NAND3X1_55 ( .A(_605_), .B(_607_), .C(_606_), .Y(_608_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_602_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_603_) );
OAI21X1 OAI21X1_110 ( .A(_602_), .B(_603_), .C(_48__3_), .Y(_604_) );
NAND2X1 NAND2X1_110 ( .A(_604_), .B(_608_), .Y(_46__3_) );
OAI21X1 OAI21X1_111 ( .A(_605_), .B(_602_), .C(_607_), .Y(_44_) );
INVX1 INVX1_56 ( .A(1'b0), .Y(_612_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_613_) );
NAND2X1 NAND2X1_111 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_614_) );
NAND3X1 NAND3X1_56 ( .A(_612_), .B(_614_), .C(_613_), .Y(_615_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_609_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_610_) );
OAI21X1 OAI21X1_112 ( .A(_609_), .B(_610_), .C(1'b0), .Y(_611_) );
NAND2X1 NAND2X1_112 ( .A(_611_), .B(_615_), .Y(_51__0_) );
OAI21X1 OAI21X1_113 ( .A(_612_), .B(_609_), .C(_614_), .Y(_53__1_) );
INVX1 INVX1_57 ( .A(_53__1_), .Y(_619_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_620_) );
NAND2X1 NAND2X1_113 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_621_) );
NAND3X1 NAND3X1_57 ( .A(_619_), .B(_621_), .C(_620_), .Y(_622_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_616_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_617_) );
OAI21X1 OAI21X1_114 ( .A(_616_), .B(_617_), .C(_53__1_), .Y(_618_) );
NAND2X1 NAND2X1_114 ( .A(_618_), .B(_622_), .Y(_51__1_) );
OAI21X1 OAI21X1_115 ( .A(_619_), .B(_616_), .C(_621_), .Y(_53__2_) );
INVX1 INVX1_58 ( .A(_53__2_), .Y(_626_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_627_) );
NAND2X1 NAND2X1_115 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_628_) );
NAND3X1 NAND3X1_58 ( .A(_626_), .B(_628_), .C(_627_), .Y(_629_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_623_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_624_) );
OAI21X1 OAI21X1_116 ( .A(_623_), .B(_624_), .C(_53__2_), .Y(_625_) );
NAND2X1 NAND2X1_116 ( .A(_625_), .B(_629_), .Y(_51__2_) );
OAI21X1 OAI21X1_117 ( .A(_626_), .B(_623_), .C(_628_), .Y(_53__3_) );
INVX1 INVX1_59 ( .A(_53__3_), .Y(_633_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_634_) );
NAND2X1 NAND2X1_117 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_635_) );
NAND3X1 NAND3X1_59 ( .A(_633_), .B(_635_), .C(_634_), .Y(_636_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_630_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_631_) );
OAI21X1 OAI21X1_118 ( .A(_630_), .B(_631_), .C(_53__3_), .Y(_632_) );
NAND2X1 NAND2X1_118 ( .A(_632_), .B(_636_), .Y(_51__3_) );
OAI21X1 OAI21X1_119 ( .A(_633_), .B(_630_), .C(_635_), .Y(_49_) );
INVX1 INVX1_60 ( .A(1'b1), .Y(_640_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_641_) );
NAND2X1 NAND2X1_119 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_642_) );
NAND3X1 NAND3X1_60 ( .A(_640_), .B(_642_), .C(_641_), .Y(_643_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_637_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_638_) );
OAI21X1 OAI21X1_120 ( .A(_637_), .B(_638_), .C(1'b1), .Y(_639_) );
NAND2X1 NAND2X1_120 ( .A(_639_), .B(_643_), .Y(_52__0_) );
OAI21X1 OAI21X1_121 ( .A(_640_), .B(_637_), .C(_642_), .Y(_54__1_) );
INVX1 INVX1_61 ( .A(_54__1_), .Y(_647_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_648_) );
NAND2X1 NAND2X1_121 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_649_) );
NAND3X1 NAND3X1_61 ( .A(_647_), .B(_649_), .C(_648_), .Y(_650_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_644_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_645_) );
OAI21X1 OAI21X1_122 ( .A(_644_), .B(_645_), .C(_54__1_), .Y(_646_) );
NAND2X1 NAND2X1_122 ( .A(_646_), .B(_650_), .Y(_52__1_) );
OAI21X1 OAI21X1_123 ( .A(_647_), .B(_644_), .C(_649_), .Y(_54__2_) );
INVX1 INVX1_62 ( .A(_54__2_), .Y(_654_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_655_) );
NAND2X1 NAND2X1_123 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_656_) );
NAND3X1 NAND3X1_62 ( .A(_654_), .B(_656_), .C(_655_), .Y(_657_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_651_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_652_) );
OAI21X1 OAI21X1_124 ( .A(_651_), .B(_652_), .C(_54__2_), .Y(_653_) );
NAND2X1 NAND2X1_124 ( .A(_653_), .B(_657_), .Y(_52__2_) );
OAI21X1 OAI21X1_125 ( .A(_654_), .B(_651_), .C(_656_), .Y(_54__3_) );
INVX1 INVX1_63 ( .A(_54__3_), .Y(_661_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_662_) );
NAND2X1 NAND2X1_125 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_663_) );
NAND3X1 NAND3X1_63 ( .A(_661_), .B(_663_), .C(_662_), .Y(_664_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_658_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_659_) );
OAI21X1 OAI21X1_126 ( .A(_658_), .B(_659_), .C(_54__3_), .Y(_660_) );
NAND2X1 NAND2X1_126 ( .A(_660_), .B(_664_), .Y(_52__3_) );
OAI21X1 OAI21X1_127 ( .A(_661_), .B(_658_), .C(_663_), .Y(_50_) );
INVX1 INVX1_64 ( .A(1'b0), .Y(_668_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_669_) );
NAND2X1 NAND2X1_127 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_670_) );
NAND3X1 NAND3X1_64 ( .A(_668_), .B(_670_), .C(_669_), .Y(_671_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_665_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_666_) );
OAI21X1 OAI21X1_128 ( .A(_665_), .B(_666_), .C(1'b0), .Y(_667_) );
NAND2X1 NAND2X1_128 ( .A(_667_), .B(_671_), .Y(_57__0_) );
OAI21X1 OAI21X1_129 ( .A(_668_), .B(_665_), .C(_670_), .Y(_59__1_) );
INVX1 INVX1_65 ( .A(_59__1_), .Y(_675_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_676_) );
NAND2X1 NAND2X1_129 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_677_) );
NAND3X1 NAND3X1_65 ( .A(_675_), .B(_677_), .C(_676_), .Y(_678_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_672_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_673_) );
OAI21X1 OAI21X1_130 ( .A(_672_), .B(_673_), .C(_59__1_), .Y(_674_) );
NAND2X1 NAND2X1_130 ( .A(_674_), .B(_678_), .Y(_57__1_) );
OAI21X1 OAI21X1_131 ( .A(_675_), .B(_672_), .C(_677_), .Y(_59__2_) );
INVX1 INVX1_66 ( .A(_59__2_), .Y(_682_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_683_) );
NAND2X1 NAND2X1_131 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_684_) );
NAND3X1 NAND3X1_66 ( .A(_682_), .B(_684_), .C(_683_), .Y(_685_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_679_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_680_) );
OAI21X1 OAI21X1_132 ( .A(_679_), .B(_680_), .C(_59__2_), .Y(_681_) );
NAND2X1 NAND2X1_132 ( .A(_681_), .B(_685_), .Y(_57__2_) );
OAI21X1 OAI21X1_133 ( .A(_682_), .B(_679_), .C(_684_), .Y(_59__3_) );
INVX1 INVX1_67 ( .A(_59__3_), .Y(_689_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_690_) );
NAND2X1 NAND2X1_133 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_691_) );
NAND3X1 NAND3X1_67 ( .A(_689_), .B(_691_), .C(_690_), .Y(_692_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_686_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_687_) );
OAI21X1 OAI21X1_134 ( .A(_686_), .B(_687_), .C(_59__3_), .Y(_688_) );
NAND2X1 NAND2X1_134 ( .A(_688_), .B(_692_), .Y(_57__3_) );
OAI21X1 OAI21X1_135 ( .A(_689_), .B(_686_), .C(_691_), .Y(_55_) );
INVX1 INVX1_68 ( .A(1'b1), .Y(_696_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_697_) );
NAND2X1 NAND2X1_135 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_698_) );
NAND3X1 NAND3X1_68 ( .A(_696_), .B(_698_), .C(_697_), .Y(_699_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_693_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_694_) );
OAI21X1 OAI21X1_136 ( .A(_693_), .B(_694_), .C(1'b1), .Y(_695_) );
NAND2X1 NAND2X1_136 ( .A(_695_), .B(_699_), .Y(_58__0_) );
OAI21X1 OAI21X1_137 ( .A(_696_), .B(_693_), .C(_698_), .Y(_60__1_) );
INVX1 INVX1_69 ( .A(_60__1_), .Y(_703_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_704_) );
NAND2X1 NAND2X1_137 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_705_) );
NAND3X1 NAND3X1_69 ( .A(_703_), .B(_705_), .C(_704_), .Y(_706_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_700_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_701_) );
OAI21X1 OAI21X1_138 ( .A(_700_), .B(_701_), .C(_60__1_), .Y(_702_) );
NAND2X1 NAND2X1_138 ( .A(_702_), .B(_706_), .Y(_58__1_) );
OAI21X1 OAI21X1_139 ( .A(_703_), .B(_700_), .C(_705_), .Y(_60__2_) );
INVX1 INVX1_70 ( .A(_60__2_), .Y(_710_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_711_) );
NAND2X1 NAND2X1_139 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_712_) );
NAND3X1 NAND3X1_70 ( .A(_710_), .B(_712_), .C(_711_), .Y(_713_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_707_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_708_) );
OAI21X1 OAI21X1_140 ( .A(_707_), .B(_708_), .C(_60__2_), .Y(_709_) );
NAND2X1 NAND2X1_140 ( .A(_709_), .B(_713_), .Y(_58__2_) );
OAI21X1 OAI21X1_141 ( .A(_710_), .B(_707_), .C(_712_), .Y(_60__3_) );
INVX1 INVX1_71 ( .A(_60__3_), .Y(_717_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_718_) );
NAND2X1 NAND2X1_141 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_719_) );
NAND3X1 NAND3X1_71 ( .A(_717_), .B(_719_), .C(_718_), .Y(_720_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_714_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_715_) );
OAI21X1 OAI21X1_142 ( .A(_714_), .B(_715_), .C(_60__3_), .Y(_716_) );
NAND2X1 NAND2X1_142 ( .A(_716_), .B(_720_), .Y(_58__3_) );
OAI21X1 OAI21X1_143 ( .A(_717_), .B(_714_), .C(_719_), .Y(_56_) );
INVX1 INVX1_72 ( .A(1'b0), .Y(_724_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_725_) );
NAND2X1 NAND2X1_143 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_726_) );
NAND3X1 NAND3X1_72 ( .A(_724_), .B(_726_), .C(_725_), .Y(_727_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_721_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_722_) );
OAI21X1 OAI21X1_144 ( .A(_721_), .B(_722_), .C(1'b0), .Y(_723_) );
NAND2X1 NAND2X1_144 ( .A(_723_), .B(_727_), .Y(rca_inst_w_SUM) );
BUFX2 BUFX2_1 ( .A(w_cout_10_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_w_SUM), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
INVX1 INVX1_73 ( .A(_1_), .Y(_61_) );
NAND2X1 NAND2X1_145 ( .A(_2_), .B(1'b0), .Y(_62_) );
OAI21X1 OAI21X1_145 ( .A(1'b0), .B(_61_), .C(_62_), .Y(w_cout_1_) );
INVX1 INVX1_74 ( .A(_3__0_), .Y(_63_) );
NAND2X1 NAND2X1_146 ( .A(_4__0_), .B(1'b0), .Y(_64_) );
OAI21X1 OAI21X1_146 ( .A(1'b0), .B(_63_), .C(_64_), .Y(_0__1_) );
INVX1 INVX1_75 ( .A(_3__1_), .Y(_65_) );
NAND2X1 NAND2X1_147 ( .A(1'b0), .B(_4__1_), .Y(_66_) );
OAI21X1 OAI21X1_147 ( .A(1'b0), .B(_65_), .C(_66_), .Y(_0__2_) );
INVX1 INVX1_76 ( .A(_3__2_), .Y(_67_) );
NAND2X1 NAND2X1_148 ( .A(1'b0), .B(_4__2_), .Y(_68_) );
OAI21X1 OAI21X1_148 ( .A(1'b0), .B(_67_), .C(_68_), .Y(_0__3_) );
INVX1 INVX1_77 ( .A(_3__3_), .Y(_69_) );
NAND2X1 NAND2X1_149 ( .A(1'b0), .B(_4__3_), .Y(_70_) );
OAI21X1 OAI21X1_149 ( .A(1'b0), .B(_69_), .C(_70_), .Y(_0__4_) );
INVX1 INVX1_78 ( .A(_7_), .Y(_71_) );
NAND2X1 NAND2X1_150 ( .A(_8_), .B(w_cout_1_), .Y(_72_) );
OAI21X1 OAI21X1_150 ( .A(w_cout_1_), .B(_71_), .C(_72_), .Y(w_cout_2_) );
INVX1 INVX1_79 ( .A(_9__0_), .Y(_73_) );
NAND2X1 NAND2X1_151 ( .A(_10__0_), .B(w_cout_1_), .Y(_74_) );
OAI21X1 OAI21X1_151 ( .A(w_cout_1_), .B(_73_), .C(_74_), .Y(_0__5_) );
INVX1 INVX1_80 ( .A(_9__1_), .Y(_75_) );
NAND2X1 NAND2X1_152 ( .A(w_cout_1_), .B(_10__1_), .Y(_76_) );
OAI21X1 OAI21X1_152 ( .A(w_cout_1_), .B(_75_), .C(_76_), .Y(_0__6_) );
INVX1 INVX1_81 ( .A(_9__2_), .Y(_77_) );
NAND2X1 NAND2X1_153 ( .A(w_cout_1_), .B(_10__2_), .Y(_78_) );
OAI21X1 OAI21X1_153 ( .A(w_cout_1_), .B(_77_), .C(_78_), .Y(_0__7_) );
INVX1 INVX1_82 ( .A(_9__3_), .Y(_79_) );
NAND2X1 NAND2X1_154 ( .A(w_cout_1_), .B(_10__3_), .Y(_80_) );
OAI21X1 OAI21X1_154 ( .A(w_cout_1_), .B(_79_), .C(_80_), .Y(_0__8_) );
INVX1 INVX1_83 ( .A(_13_), .Y(_81_) );
NAND2X1 NAND2X1_155 ( .A(_14_), .B(w_cout_2_), .Y(_82_) );
OAI21X1 OAI21X1_155 ( .A(w_cout_2_), .B(_81_), .C(_82_), .Y(w_cout_3_) );
INVX1 INVX1_84 ( .A(_15__0_), .Y(_83_) );
NAND2X1 NAND2X1_156 ( .A(_16__0_), .B(w_cout_2_), .Y(_84_) );
OAI21X1 OAI21X1_156 ( .A(w_cout_2_), .B(_83_), .C(_84_), .Y(_0__9_) );
INVX1 INVX1_85 ( .A(_15__1_), .Y(_85_) );
NAND2X1 NAND2X1_157 ( .A(w_cout_2_), .B(_16__1_), .Y(_86_) );
OAI21X1 OAI21X1_157 ( .A(w_cout_2_), .B(_85_), .C(_86_), .Y(_0__10_) );
INVX1 INVX1_86 ( .A(_15__2_), .Y(_87_) );
NAND2X1 NAND2X1_158 ( .A(w_cout_2_), .B(_16__2_), .Y(_88_) );
OAI21X1 OAI21X1_158 ( .A(w_cout_2_), .B(_87_), .C(_88_), .Y(_0__11_) );
INVX1 INVX1_87 ( .A(_15__3_), .Y(_89_) );
NAND2X1 NAND2X1_159 ( .A(w_cout_2_), .B(_16__3_), .Y(_90_) );
OAI21X1 OAI21X1_159 ( .A(w_cout_2_), .B(_89_), .C(_90_), .Y(_0__12_) );
INVX1 INVX1_88 ( .A(_19_), .Y(_91_) );
NAND2X1 NAND2X1_160 ( .A(_20_), .B(w_cout_3_), .Y(_92_) );
OAI21X1 OAI21X1_160 ( .A(w_cout_3_), .B(_91_), .C(_92_), .Y(w_cout_4_) );
INVX1 INVX1_89 ( .A(_21__0_), .Y(_93_) );
NAND2X1 NAND2X1_161 ( .A(_22__0_), .B(w_cout_3_), .Y(_94_) );
OAI21X1 OAI21X1_161 ( .A(w_cout_3_), .B(_93_), .C(_94_), .Y(_0__13_) );
INVX1 INVX1_90 ( .A(_21__1_), .Y(_95_) );
NAND2X1 NAND2X1_162 ( .A(w_cout_3_), .B(_22__1_), .Y(_96_) );
OAI21X1 OAI21X1_162 ( .A(w_cout_3_), .B(_95_), .C(_96_), .Y(_0__14_) );
INVX1 INVX1_91 ( .A(_21__2_), .Y(_97_) );
NAND2X1 NAND2X1_163 ( .A(w_cout_3_), .B(_22__2_), .Y(_98_) );
OAI21X1 OAI21X1_163 ( .A(w_cout_3_), .B(_97_), .C(_98_), .Y(_0__15_) );
INVX1 INVX1_92 ( .A(_21__3_), .Y(_99_) );
NAND2X1 NAND2X1_164 ( .A(w_cout_3_), .B(_22__3_), .Y(_100_) );
OAI21X1 OAI21X1_164 ( .A(w_cout_3_), .B(_99_), .C(_100_), .Y(_0__16_) );
INVX1 INVX1_93 ( .A(_25_), .Y(_101_) );
NAND2X1 NAND2X1_165 ( .A(_26_), .B(w_cout_4_), .Y(_102_) );
OAI21X1 OAI21X1_165 ( .A(w_cout_4_), .B(_101_), .C(_102_), .Y(w_cout_5_) );
INVX1 INVX1_94 ( .A(_27__0_), .Y(_103_) );
NAND2X1 NAND2X1_166 ( .A(_28__0_), .B(w_cout_4_), .Y(_104_) );
OAI21X1 OAI21X1_166 ( .A(w_cout_4_), .B(_103_), .C(_104_), .Y(_0__17_) );
INVX1 INVX1_95 ( .A(_27__1_), .Y(_105_) );
NAND2X1 NAND2X1_167 ( .A(w_cout_4_), .B(_28__1_), .Y(_106_) );
OAI21X1 OAI21X1_167 ( .A(w_cout_4_), .B(_105_), .C(_106_), .Y(_0__18_) );
INVX1 INVX1_96 ( .A(_27__2_), .Y(_107_) );
NAND2X1 NAND2X1_168 ( .A(w_cout_4_), .B(_28__2_), .Y(_108_) );
OAI21X1 OAI21X1_168 ( .A(w_cout_4_), .B(_107_), .C(_108_), .Y(_0__19_) );
INVX1 INVX1_97 ( .A(_27__3_), .Y(_109_) );
NAND2X1 NAND2X1_169 ( .A(w_cout_4_), .B(_28__3_), .Y(_110_) );
OAI21X1 OAI21X1_169 ( .A(w_cout_4_), .B(_109_), .C(_110_), .Y(_0__20_) );
INVX1 INVX1_98 ( .A(_31_), .Y(_111_) );
NAND2X1 NAND2X1_170 ( .A(_32_), .B(w_cout_5_), .Y(_112_) );
OAI21X1 OAI21X1_170 ( .A(w_cout_5_), .B(_111_), .C(_112_), .Y(w_cout_6_) );
INVX1 INVX1_99 ( .A(_33__0_), .Y(_113_) );
NAND2X1 NAND2X1_171 ( .A(_34__0_), .B(w_cout_5_), .Y(_114_) );
OAI21X1 OAI21X1_171 ( .A(w_cout_5_), .B(_113_), .C(_114_), .Y(_0__21_) );
INVX1 INVX1_100 ( .A(_33__1_), .Y(_115_) );
NAND2X1 NAND2X1_172 ( .A(w_cout_5_), .B(_34__1_), .Y(_116_) );
OAI21X1 OAI21X1_172 ( .A(w_cout_5_), .B(_115_), .C(_116_), .Y(_0__22_) );
INVX1 INVX1_101 ( .A(_33__2_), .Y(_117_) );
NAND2X1 NAND2X1_173 ( .A(w_cout_5_), .B(_34__2_), .Y(_118_) );
OAI21X1 OAI21X1_173 ( .A(w_cout_5_), .B(_117_), .C(_118_), .Y(_0__23_) );
INVX1 INVX1_102 ( .A(_33__3_), .Y(_119_) );
NAND2X1 NAND2X1_174 ( .A(w_cout_5_), .B(_34__3_), .Y(_120_) );
OAI21X1 OAI21X1_174 ( .A(w_cout_5_), .B(_119_), .C(_120_), .Y(_0__24_) );
INVX1 INVX1_103 ( .A(_37_), .Y(_121_) );
NAND2X1 NAND2X1_175 ( .A(_38_), .B(w_cout_6_), .Y(_122_) );
OAI21X1 OAI21X1_175 ( .A(w_cout_6_), .B(_121_), .C(_122_), .Y(w_cout_7_) );
INVX1 INVX1_104 ( .A(_39__0_), .Y(_123_) );
NAND2X1 NAND2X1_176 ( .A(_40__0_), .B(w_cout_6_), .Y(_124_) );
OAI21X1 OAI21X1_176 ( .A(w_cout_6_), .B(_123_), .C(_124_), .Y(_0__25_) );
INVX1 INVX1_105 ( .A(_39__1_), .Y(_125_) );
NAND2X1 NAND2X1_177 ( .A(w_cout_6_), .B(_40__1_), .Y(_126_) );
OAI21X1 OAI21X1_177 ( .A(w_cout_6_), .B(_125_), .C(_126_), .Y(_0__26_) );
INVX1 INVX1_106 ( .A(_39__2_), .Y(_127_) );
NAND2X1 NAND2X1_178 ( .A(w_cout_6_), .B(_40__2_), .Y(_128_) );
OAI21X1 OAI21X1_178 ( .A(w_cout_6_), .B(_127_), .C(_128_), .Y(_0__27_) );
INVX1 INVX1_107 ( .A(_39__3_), .Y(_129_) );
NAND2X1 NAND2X1_179 ( .A(w_cout_6_), .B(_40__3_), .Y(_130_) );
OAI21X1 OAI21X1_179 ( .A(w_cout_6_), .B(_129_), .C(_130_), .Y(_0__28_) );
INVX1 INVX1_108 ( .A(_43_), .Y(_131_) );
NAND2X1 NAND2X1_180 ( .A(_44_), .B(w_cout_7_), .Y(_132_) );
OAI21X1 OAI21X1_180 ( .A(w_cout_7_), .B(_131_), .C(_132_), .Y(w_cout_8_) );
INVX1 INVX1_109 ( .A(_45__0_), .Y(_133_) );
NAND2X1 NAND2X1_181 ( .A(_46__0_), .B(w_cout_7_), .Y(_134_) );
OAI21X1 OAI21X1_181 ( .A(w_cout_7_), .B(_133_), .C(_134_), .Y(_0__29_) );
INVX1 INVX1_110 ( .A(_45__1_), .Y(_135_) );
NAND2X1 NAND2X1_182 ( .A(w_cout_7_), .B(_46__1_), .Y(_136_) );
OAI21X1 OAI21X1_182 ( .A(w_cout_7_), .B(_135_), .C(_136_), .Y(_0__30_) );
INVX1 INVX1_111 ( .A(_45__2_), .Y(_137_) );
NAND2X1 NAND2X1_183 ( .A(w_cout_7_), .B(_46__2_), .Y(_138_) );
OAI21X1 OAI21X1_183 ( .A(w_cout_7_), .B(_137_), .C(_138_), .Y(_0__31_) );
INVX1 INVX1_112 ( .A(_45__3_), .Y(_139_) );
NAND2X1 NAND2X1_184 ( .A(w_cout_7_), .B(_46__3_), .Y(_140_) );
OAI21X1 OAI21X1_184 ( .A(w_cout_7_), .B(_139_), .C(_140_), .Y(_0__32_) );
INVX1 INVX1_113 ( .A(_49_), .Y(_141_) );
NAND2X1 NAND2X1_185 ( .A(_50_), .B(w_cout_8_), .Y(_142_) );
OAI21X1 OAI21X1_185 ( .A(w_cout_8_), .B(_141_), .C(_142_), .Y(w_cout_9_) );
INVX1 INVX1_114 ( .A(_51__0_), .Y(_143_) );
NAND2X1 NAND2X1_186 ( .A(_52__0_), .B(w_cout_8_), .Y(_144_) );
OAI21X1 OAI21X1_186 ( .A(w_cout_8_), .B(_143_), .C(_144_), .Y(_0__33_) );
INVX1 INVX1_115 ( .A(_51__1_), .Y(_145_) );
NAND2X1 NAND2X1_187 ( .A(w_cout_8_), .B(_52__1_), .Y(_146_) );
OAI21X1 OAI21X1_187 ( .A(w_cout_8_), .B(_145_), .C(_146_), .Y(_0__34_) );
INVX1 INVX1_116 ( .A(_51__2_), .Y(_147_) );
NAND2X1 NAND2X1_188 ( .A(w_cout_8_), .B(_52__2_), .Y(_148_) );
OAI21X1 OAI21X1_188 ( .A(w_cout_8_), .B(_147_), .C(_148_), .Y(_0__35_) );
INVX1 INVX1_117 ( .A(_51__3_), .Y(_149_) );
NAND2X1 NAND2X1_189 ( .A(w_cout_8_), .B(_52__3_), .Y(_150_) );
OAI21X1 OAI21X1_189 ( .A(w_cout_8_), .B(_149_), .C(_150_), .Y(_0__36_) );
INVX1 INVX1_118 ( .A(_55_), .Y(_151_) );
NAND2X1 NAND2X1_190 ( .A(_56_), .B(w_cout_9_), .Y(_152_) );
OAI21X1 OAI21X1_190 ( .A(w_cout_9_), .B(_151_), .C(_152_), .Y(w_cout_10_) );
INVX1 INVX1_119 ( .A(_57__0_), .Y(_153_) );
NAND2X1 NAND2X1_191 ( .A(_58__0_), .B(w_cout_9_), .Y(_154_) );
OAI21X1 OAI21X1_191 ( .A(w_cout_9_), .B(_153_), .C(_154_), .Y(_0__37_) );
INVX1 INVX1_120 ( .A(_57__1_), .Y(_155_) );
NAND2X1 NAND2X1_192 ( .A(w_cout_9_), .B(_58__1_), .Y(_156_) );
OAI21X1 OAI21X1_192 ( .A(w_cout_9_), .B(_155_), .C(_156_), .Y(_0__38_) );
INVX1 INVX1_121 ( .A(_57__2_), .Y(_157_) );
NAND2X1 NAND2X1_193 ( .A(w_cout_9_), .B(_58__2_), .Y(_158_) );
OAI21X1 OAI21X1_193 ( .A(w_cout_9_), .B(_157_), .C(_158_), .Y(_0__39_) );
INVX1 INVX1_122 ( .A(_57__3_), .Y(_159_) );
NAND2X1 NAND2X1_194 ( .A(w_cout_9_), .B(_58__3_), .Y(_160_) );
OAI21X1 OAI21X1_194 ( .A(w_cout_9_), .B(_159_), .C(_160_), .Y(_0__40_) );
INVX1 INVX1_123 ( .A(1'b0), .Y(_164_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_165_) );
NAND2X1 NAND2X1_195 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_166_) );
NAND3X1 NAND3X1_73 ( .A(_164_), .B(_166_), .C(_165_), .Y(_167_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_161_) );
AND2X2 AND2X2_73 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_162_) );
OAI21X1 OAI21X1_195 ( .A(_161_), .B(_162_), .C(1'b0), .Y(_163_) );
NAND2X1 NAND2X1_196 ( .A(_163_), .B(_167_), .Y(_3__0_) );
OAI21X1 OAI21X1_196 ( .A(_164_), .B(_161_), .C(_166_), .Y(_5__1_) );
INVX1 INVX1_124 ( .A(_5__1_), .Y(_171_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_172_) );
NAND2X1 NAND2X1_197 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_173_) );
NAND3X1 NAND3X1_74 ( .A(_171_), .B(_173_), .C(_172_), .Y(_174_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_168_) );
AND2X2 AND2X2_74 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_169_) );
OAI21X1 OAI21X1_197 ( .A(_168_), .B(_169_), .C(_5__1_), .Y(_170_) );
NAND2X1 NAND2X1_198 ( .A(_170_), .B(_174_), .Y(_3__1_) );
OAI21X1 OAI21X1_198 ( .A(_171_), .B(_168_), .C(_173_), .Y(_5__2_) );
INVX1 INVX1_125 ( .A(_5__2_), .Y(_178_) );
OR2X2 OR2X2_75 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_179_) );
NAND2X1 NAND2X1_199 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_180_) );
NAND3X1 NAND3X1_75 ( .A(_178_), .B(_180_), .C(_179_), .Y(_181_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_175_) );
AND2X2 AND2X2_75 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_176_) );
OAI21X1 OAI21X1_199 ( .A(_175_), .B(_176_), .C(_5__2_), .Y(_177_) );
NAND2X1 NAND2X1_200 ( .A(_177_), .B(_181_), .Y(_3__2_) );
OAI21X1 OAI21X1_200 ( .A(_178_), .B(_175_), .C(_180_), .Y(_5__3_) );
INVX1 INVX1_126 ( .A(_5__3_), .Y(_185_) );
OR2X2 OR2X2_76 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_186_) );
NAND2X1 NAND2X1_201 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_187_) );
NAND3X1 NAND3X1_76 ( .A(_185_), .B(_187_), .C(_186_), .Y(_188_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_182_) );
AND2X2 AND2X2_76 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_183_) );
OAI21X1 OAI21X1_201 ( .A(_182_), .B(_183_), .C(_5__3_), .Y(_184_) );
NAND2X1 NAND2X1_202 ( .A(_184_), .B(_188_), .Y(_3__3_) );
OAI21X1 OAI21X1_202 ( .A(_185_), .B(_182_), .C(_187_), .Y(_1_) );
INVX1 INVX1_127 ( .A(1'b1), .Y(_192_) );
OR2X2 OR2X2_77 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_193_) );
NAND2X1 NAND2X1_203 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_194_) );
NAND3X1 NAND3X1_77 ( .A(_192_), .B(_194_), .C(_193_), .Y(_195_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_189_) );
AND2X2 AND2X2_77 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_190_) );
OAI21X1 OAI21X1_203 ( .A(_189_), .B(_190_), .C(1'b1), .Y(_191_) );
NAND2X1 NAND2X1_204 ( .A(_191_), .B(_195_), .Y(_4__0_) );
OAI21X1 OAI21X1_204 ( .A(_192_), .B(_189_), .C(_194_), .Y(_6__1_) );
INVX1 INVX1_128 ( .A(_6__1_), .Y(_199_) );
OR2X2 OR2X2_78 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_200_) );
NAND2X1 NAND2X1_205 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_201_) );
NAND3X1 NAND3X1_78 ( .A(_199_), .B(_201_), .C(_200_), .Y(_202_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_196_) );
AND2X2 AND2X2_78 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_197_) );
OAI21X1 OAI21X1_205 ( .A(_196_), .B(_197_), .C(_6__1_), .Y(_198_) );
NAND2X1 NAND2X1_206 ( .A(_198_), .B(_202_), .Y(_4__1_) );
OAI21X1 OAI21X1_206 ( .A(_199_), .B(_196_), .C(_201_), .Y(_6__2_) );
INVX1 INVX1_129 ( .A(_6__2_), .Y(_206_) );
OR2X2 OR2X2_79 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_207_) );
NAND2X1 NAND2X1_207 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_208_) );
NAND3X1 NAND3X1_79 ( .A(_206_), .B(_208_), .C(_207_), .Y(_209_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_203_) );
AND2X2 AND2X2_79 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_204_) );
OAI21X1 OAI21X1_207 ( .A(_203_), .B(_204_), .C(_6__2_), .Y(_205_) );
NAND2X1 NAND2X1_208 ( .A(_205_), .B(_209_), .Y(_4__2_) );
OAI21X1 OAI21X1_208 ( .A(_206_), .B(_203_), .C(_208_), .Y(_6__3_) );
INVX1 INVX1_130 ( .A(_6__3_), .Y(_213_) );
OR2X2 OR2X2_80 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_214_) );
NAND2X1 NAND2X1_209 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_215_) );
NAND3X1 NAND3X1_80 ( .A(_213_), .B(_215_), .C(_214_), .Y(_216_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_210_) );
AND2X2 AND2X2_80 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_211_) );
OAI21X1 OAI21X1_209 ( .A(_210_), .B(_211_), .C(_6__3_), .Y(_212_) );
NAND2X1 NAND2X1_210 ( .A(_212_), .B(_216_), .Y(_4__3_) );
OAI21X1 OAI21X1_210 ( .A(_213_), .B(_210_), .C(_215_), .Y(_2_) );
INVX1 INVX1_131 ( .A(1'b0), .Y(_220_) );
OR2X2 OR2X2_81 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_221_) );
NAND2X1 NAND2X1_211 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_222_) );
NAND3X1 NAND3X1_81 ( .A(_220_), .B(_222_), .C(_221_), .Y(_223_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_217_) );
AND2X2 AND2X2_81 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_218_) );
OAI21X1 OAI21X1_211 ( .A(_217_), .B(_218_), .C(1'b0), .Y(_219_) );
NAND2X1 NAND2X1_212 ( .A(_219_), .B(_223_), .Y(_9__0_) );
BUFX2 BUFX2_43 ( .A(rca_inst_w_SUM), .Y(_0__0_) );
BUFX2 BUFX2_44 ( .A(1'b0), .Y(_5__0_) );
BUFX2 BUFX2_45 ( .A(_1_), .Y(_5__4_) );
BUFX2 BUFX2_46 ( .A(1'b1), .Y(_6__0_) );
BUFX2 BUFX2_47 ( .A(_2_), .Y(_6__4_) );
BUFX2 BUFX2_48 ( .A(1'b0), .Y(_11__0_) );
BUFX2 BUFX2_49 ( .A(_7_), .Y(_11__4_) );
BUFX2 BUFX2_50 ( .A(1'b1), .Y(_12__0_) );
BUFX2 BUFX2_51 ( .A(_8_), .Y(_12__4_) );
BUFX2 BUFX2_52 ( .A(1'b0), .Y(_17__0_) );
BUFX2 BUFX2_53 ( .A(_13_), .Y(_17__4_) );
BUFX2 BUFX2_54 ( .A(1'b1), .Y(_18__0_) );
BUFX2 BUFX2_55 ( .A(_14_), .Y(_18__4_) );
BUFX2 BUFX2_56 ( .A(1'b0), .Y(_23__0_) );
BUFX2 BUFX2_57 ( .A(_19_), .Y(_23__4_) );
BUFX2 BUFX2_58 ( .A(1'b1), .Y(_24__0_) );
BUFX2 BUFX2_59 ( .A(_20_), .Y(_24__4_) );
BUFX2 BUFX2_60 ( .A(1'b0), .Y(_29__0_) );
BUFX2 BUFX2_61 ( .A(_25_), .Y(_29__4_) );
BUFX2 BUFX2_62 ( .A(1'b1), .Y(_30__0_) );
BUFX2 BUFX2_63 ( .A(_26_), .Y(_30__4_) );
BUFX2 BUFX2_64 ( .A(1'b0), .Y(_35__0_) );
BUFX2 BUFX2_65 ( .A(_31_), .Y(_35__4_) );
BUFX2 BUFX2_66 ( .A(1'b1), .Y(_36__0_) );
BUFX2 BUFX2_67 ( .A(_32_), .Y(_36__4_) );
BUFX2 BUFX2_68 ( .A(1'b0), .Y(_41__0_) );
BUFX2 BUFX2_69 ( .A(_37_), .Y(_41__4_) );
BUFX2 BUFX2_70 ( .A(1'b1), .Y(_42__0_) );
BUFX2 BUFX2_71 ( .A(_38_), .Y(_42__4_) );
BUFX2 BUFX2_72 ( .A(1'b0), .Y(_47__0_) );
BUFX2 BUFX2_73 ( .A(_43_), .Y(_47__4_) );
BUFX2 BUFX2_74 ( .A(1'b1), .Y(_48__0_) );
BUFX2 BUFX2_75 ( .A(_44_), .Y(_48__4_) );
BUFX2 BUFX2_76 ( .A(1'b0), .Y(_53__0_) );
BUFX2 BUFX2_77 ( .A(_49_), .Y(_53__4_) );
BUFX2 BUFX2_78 ( .A(1'b1), .Y(_54__0_) );
BUFX2 BUFX2_79 ( .A(_50_), .Y(_54__4_) );
BUFX2 BUFX2_80 ( .A(1'b0), .Y(_59__0_) );
BUFX2 BUFX2_81 ( .A(_55_), .Y(_59__4_) );
BUFX2 BUFX2_82 ( .A(1'b1), .Y(_60__0_) );
BUFX2 BUFX2_83 ( .A(_56_), .Y(_60__4_) );
BUFX2 BUFX2_84 ( .A(1'b0), .Y(w_cout_0_) );
endmodule
