module CSkipA_40bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [39:0] i_add_term1;
input [39:0] i_add_term2;
output [39:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

AND2X2 AND2X2_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_425_) );
OAI21X1 OAI21X1_1 ( .A(_424_), .B(_425_), .C(gnd), .Y(_426_) );
NAND2X1 NAND2X1_1 ( .A(_426_), .B(_430_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_2 ( .A(_427_), .B(_424_), .C(_429_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_1 ( .A(rca_inst_fa3_i_carry), .Y(_434_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_435_) );
NAND2X1 NAND2X1_2 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_436_) );
NAND3X1 NAND3X1_1 ( .A(_434_), .B(_436_), .C(_435_), .Y(_437_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_431_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_432_) );
OAI21X1 OAI21X1_3 ( .A(_431_), .B(_432_), .C(rca_inst_fa3_i_carry), .Y(_433_) );
NAND2X1 NAND2X1_3 ( .A(_433_), .B(_437_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_4 ( .A(_434_), .B(_431_), .C(_436_), .Y(cout0) );
INVX1 INVX1_2 ( .A(rca_inst_fa0_o_carry), .Y(_441_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_442_) );
NAND2X1 NAND2X1_4 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_443_) );
NAND3X1 NAND3X1_2 ( .A(_441_), .B(_443_), .C(_442_), .Y(_444_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_438_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_439_) );
OAI21X1 OAI21X1_5 ( .A(_438_), .B(_439_), .C(rca_inst_fa0_o_carry), .Y(_440_) );
NAND2X1 NAND2X1_5 ( .A(_440_), .B(_444_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_6 ( .A(_441_), .B(_438_), .C(_443_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_3 ( .A(rca_inst_fa_1__o_carry), .Y(_448_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_449_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_450_) );
NAND3X1 NAND3X1_3 ( .A(_448_), .B(_450_), .C(_449_), .Y(_451_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_445_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_446_) );
OAI21X1 OAI21X1_7 ( .A(_445_), .B(_446_), .C(rca_inst_fa_1__o_carry), .Y(_447_) );
NAND2X1 NAND2X1_7 ( .A(_447_), .B(_451_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_8 ( .A(_448_), .B(_445_), .C(_450_), .Y(rca_inst_fa3_i_carry) );
INVX1 INVX1_4 ( .A(i_add_term1[0]), .Y(_452_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[0]), .B(_452_), .Y(_453_) );
INVX1 INVX1_5 ( .A(i_add_term2[0]), .Y(_454_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term1[0]), .B(_454_), .Y(_455_) );
INVX1 INVX1_6 ( .A(i_add_term1[1]), .Y(_456_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[1]), .B(_456_), .Y(_457_) );
INVX1 INVX1_7 ( .A(i_add_term2[1]), .Y(_458_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term1[1]), .B(_458_), .Y(_459_) );
OAI22X1 OAI22X1_1 ( .A(_453_), .B(_455_), .C(_457_), .D(_459_), .Y(_460_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_461_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_462_) );
NOR2X1 NOR2X1_9 ( .A(_461_), .B(_462_), .Y(_463_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_464_) );
NAND2X1 NAND2X1_8 ( .A(_463_), .B(_464_), .Y(_465_) );
NOR2X1 NOR2X1_10 ( .A(_460_), .B(_465_), .Y(skip0_P) );
INVX1 INVX1_8 ( .A(cout0), .Y(_466_) );
NAND2X1 NAND2X1_9 ( .A(gnd), .B(skip0_P), .Y(_467_) );
OAI21X1 OAI21X1_9 ( .A(skip0_P), .B(_466_), .C(_467_), .Y(skip0_cin_next) );
BUFX2 BUFX2_1 ( .A(w_cout_9_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
INVX1 INVX1_9 ( .A(skip0_cin_next), .Y(_31_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_32_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_33_) );
NAND3X1 NAND3X1_4 ( .A(_31_), .B(_33_), .C(_32_), .Y(_34_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_28_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_29_) );
OAI21X1 OAI21X1_10 ( .A(_28_), .B(_29_), .C(skip0_cin_next), .Y(_30_) );
NAND2X1 NAND2X1_11 ( .A(_30_), .B(_34_), .Y(_0__4_) );
OAI21X1 OAI21X1_11 ( .A(_31_), .B(_28_), .C(_33_), .Y(_2__1_) );
INVX1 INVX1_10 ( .A(_2__3_), .Y(_38_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_39_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_40_) );
NAND3X1 NAND3X1_5 ( .A(_38_), .B(_40_), .C(_39_), .Y(_41_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_35_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_36_) );
OAI21X1 OAI21X1_12 ( .A(_35_), .B(_36_), .C(_2__3_), .Y(_37_) );
NAND2X1 NAND2X1_13 ( .A(_37_), .B(_41_), .Y(_0__7_) );
OAI21X1 OAI21X1_13 ( .A(_38_), .B(_35_), .C(_40_), .Y(_1_) );
INVX1 INVX1_11 ( .A(_2__1_), .Y(_45_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_46_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_47_) );
NAND3X1 NAND3X1_6 ( .A(_45_), .B(_47_), .C(_46_), .Y(_48_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_42_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_43_) );
OAI21X1 OAI21X1_14 ( .A(_42_), .B(_43_), .C(_2__1_), .Y(_44_) );
NAND2X1 NAND2X1_15 ( .A(_44_), .B(_48_), .Y(_0__5_) );
OAI21X1 OAI21X1_15 ( .A(_45_), .B(_42_), .C(_47_), .Y(_2__2_) );
INVX1 INVX1_12 ( .A(_2__2_), .Y(_52_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_53_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_54_) );
NAND3X1 NAND3X1_7 ( .A(_52_), .B(_54_), .C(_53_), .Y(_55_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_49_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_50_) );
OAI21X1 OAI21X1_16 ( .A(_49_), .B(_50_), .C(_2__2_), .Y(_51_) );
NAND2X1 NAND2X1_17 ( .A(_51_), .B(_55_), .Y(_0__6_) );
OAI21X1 OAI21X1_17 ( .A(_52_), .B(_49_), .C(_54_), .Y(_2__3_) );
INVX1 INVX1_13 ( .A(i_add_term1[4]), .Y(_56_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[4]), .B(_56_), .Y(_57_) );
INVX1 INVX1_14 ( .A(i_add_term2[4]), .Y(_58_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term1[4]), .B(_58_), .Y(_59_) );
INVX1 INVX1_15 ( .A(i_add_term1[5]), .Y(_60_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[5]), .B(_60_), .Y(_61_) );
INVX1 INVX1_16 ( .A(i_add_term2[5]), .Y(_62_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term1[5]), .B(_62_), .Y(_63_) );
OAI22X1 OAI22X1_2 ( .A(_57_), .B(_59_), .C(_61_), .D(_63_), .Y(_64_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_65_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_66_) );
NOR2X1 NOR2X1_20 ( .A(_65_), .B(_66_), .Y(_67_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_68_) );
NAND2X1 NAND2X1_18 ( .A(_67_), .B(_68_), .Y(_69_) );
NOR2X1 NOR2X1_21 ( .A(_64_), .B(_69_), .Y(_3_) );
INVX1 INVX1_17 ( .A(_1_), .Y(_70_) );
NAND2X1 NAND2X1_19 ( .A(gnd), .B(_3_), .Y(_71_) );
OAI21X1 OAI21X1_18 ( .A(_3_), .B(_70_), .C(_71_), .Y(w_cout_1_) );
INVX1 INVX1_18 ( .A(w_cout_1_), .Y(_75_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_76_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_77_) );
NAND3X1 NAND3X1_8 ( .A(_75_), .B(_77_), .C(_76_), .Y(_78_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_72_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_73_) );
OAI21X1 OAI21X1_19 ( .A(_72_), .B(_73_), .C(w_cout_1_), .Y(_74_) );
NAND2X1 NAND2X1_21 ( .A(_74_), .B(_78_), .Y(_0__8_) );
OAI21X1 OAI21X1_20 ( .A(_75_), .B(_72_), .C(_77_), .Y(_5__1_) );
INVX1 INVX1_19 ( .A(_5__3_), .Y(_82_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_83_) );
NAND2X1 NAND2X1_22 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_84_) );
NAND3X1 NAND3X1_9 ( .A(_82_), .B(_84_), .C(_83_), .Y(_85_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_79_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_80_) );
OAI21X1 OAI21X1_21 ( .A(_79_), .B(_80_), .C(_5__3_), .Y(_81_) );
NAND2X1 NAND2X1_23 ( .A(_81_), .B(_85_), .Y(_0__11_) );
OAI21X1 OAI21X1_22 ( .A(_82_), .B(_79_), .C(_84_), .Y(_4_) );
INVX1 INVX1_20 ( .A(_5__1_), .Y(_89_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_90_) );
NAND2X1 NAND2X1_24 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_91_) );
NAND3X1 NAND3X1_10 ( .A(_89_), .B(_91_), .C(_90_), .Y(_92_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_86_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_87_) );
OAI21X1 OAI21X1_23 ( .A(_86_), .B(_87_), .C(_5__1_), .Y(_88_) );
NAND2X1 NAND2X1_25 ( .A(_88_), .B(_92_), .Y(_0__9_) );
OAI21X1 OAI21X1_24 ( .A(_89_), .B(_86_), .C(_91_), .Y(_5__2_) );
INVX1 INVX1_21 ( .A(_5__2_), .Y(_96_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_97_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_98_) );
NAND3X1 NAND3X1_11 ( .A(_96_), .B(_98_), .C(_97_), .Y(_99_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_93_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_94_) );
OAI21X1 OAI21X1_25 ( .A(_93_), .B(_94_), .C(_5__2_), .Y(_95_) );
NAND2X1 NAND2X1_27 ( .A(_95_), .B(_99_), .Y(_0__10_) );
OAI21X1 OAI21X1_26 ( .A(_96_), .B(_93_), .C(_98_), .Y(_5__3_) );
INVX1 INVX1_22 ( .A(i_add_term1[8]), .Y(_100_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[8]), .B(_100_), .Y(_101_) );
INVX1 INVX1_23 ( .A(i_add_term2[8]), .Y(_102_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term1[8]), .B(_102_), .Y(_103_) );
INVX1 INVX1_24 ( .A(i_add_term1[9]), .Y(_104_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[9]), .B(_104_), .Y(_105_) );
INVX1 INVX1_25 ( .A(i_add_term2[9]), .Y(_106_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term1[9]), .B(_106_), .Y(_107_) );
OAI22X1 OAI22X1_3 ( .A(_101_), .B(_103_), .C(_105_), .D(_107_), .Y(_108_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_109_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_110_) );
NOR2X1 NOR2X1_31 ( .A(_109_), .B(_110_), .Y(_111_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_112_) );
NAND2X1 NAND2X1_28 ( .A(_111_), .B(_112_), .Y(_113_) );
NOR2X1 NOR2X1_32 ( .A(_108_), .B(_113_), .Y(_6_) );
INVX1 INVX1_26 ( .A(_4_), .Y(_114_) );
NAND2X1 NAND2X1_29 ( .A(gnd), .B(_6_), .Y(_115_) );
OAI21X1 OAI21X1_27 ( .A(_6_), .B(_114_), .C(_115_), .Y(w_cout_2_) );
INVX1 INVX1_27 ( .A(w_cout_2_), .Y(_119_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_120_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_121_) );
NAND3X1 NAND3X1_12 ( .A(_119_), .B(_121_), .C(_120_), .Y(_122_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_116_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_117_) );
OAI21X1 OAI21X1_28 ( .A(_116_), .B(_117_), .C(w_cout_2_), .Y(_118_) );
NAND2X1 NAND2X1_31 ( .A(_118_), .B(_122_), .Y(_0__12_) );
OAI21X1 OAI21X1_29 ( .A(_119_), .B(_116_), .C(_121_), .Y(_8__1_) );
INVX1 INVX1_28 ( .A(_8__3_), .Y(_126_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_127_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_128_) );
NAND3X1 NAND3X1_13 ( .A(_126_), .B(_128_), .C(_127_), .Y(_129_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_123_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_124_) );
OAI21X1 OAI21X1_30 ( .A(_123_), .B(_124_), .C(_8__3_), .Y(_125_) );
NAND2X1 NAND2X1_33 ( .A(_125_), .B(_129_), .Y(_0__15_) );
OAI21X1 OAI21X1_31 ( .A(_126_), .B(_123_), .C(_128_), .Y(_7_) );
INVX1 INVX1_29 ( .A(_8__1_), .Y(_133_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_134_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_135_) );
NAND3X1 NAND3X1_14 ( .A(_133_), .B(_135_), .C(_134_), .Y(_136_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_130_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_131_) );
OAI21X1 OAI21X1_32 ( .A(_130_), .B(_131_), .C(_8__1_), .Y(_132_) );
NAND2X1 NAND2X1_35 ( .A(_132_), .B(_136_), .Y(_0__13_) );
OAI21X1 OAI21X1_33 ( .A(_133_), .B(_130_), .C(_135_), .Y(_8__2_) );
INVX1 INVX1_30 ( .A(_8__2_), .Y(_140_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_141_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_142_) );
NAND3X1 NAND3X1_15 ( .A(_140_), .B(_142_), .C(_141_), .Y(_143_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_137_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_138_) );
OAI21X1 OAI21X1_34 ( .A(_137_), .B(_138_), .C(_8__2_), .Y(_139_) );
NAND2X1 NAND2X1_37 ( .A(_139_), .B(_143_), .Y(_0__14_) );
OAI21X1 OAI21X1_35 ( .A(_140_), .B(_137_), .C(_142_), .Y(_8__3_) );
INVX1 INVX1_31 ( .A(i_add_term1[12]), .Y(_144_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[12]), .B(_144_), .Y(_145_) );
INVX1 INVX1_32 ( .A(i_add_term2[12]), .Y(_146_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term1[12]), .B(_146_), .Y(_147_) );
INVX1 INVX1_33 ( .A(i_add_term1[13]), .Y(_148_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[13]), .B(_148_), .Y(_149_) );
INVX1 INVX1_34 ( .A(i_add_term2[13]), .Y(_150_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term1[13]), .B(_150_), .Y(_151_) );
OAI22X1 OAI22X1_4 ( .A(_145_), .B(_147_), .C(_149_), .D(_151_), .Y(_152_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_153_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_154_) );
NOR2X1 NOR2X1_42 ( .A(_153_), .B(_154_), .Y(_155_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_156_) );
NAND2X1 NAND2X1_38 ( .A(_155_), .B(_156_), .Y(_157_) );
NOR2X1 NOR2X1_43 ( .A(_152_), .B(_157_), .Y(_9_) );
INVX1 INVX1_35 ( .A(_7_), .Y(_158_) );
NAND2X1 NAND2X1_39 ( .A(gnd), .B(_9_), .Y(_159_) );
OAI21X1 OAI21X1_36 ( .A(_9_), .B(_158_), .C(_159_), .Y(w_cout_3_) );
INVX1 INVX1_36 ( .A(w_cout_3_), .Y(_163_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_164_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_165_) );
NAND3X1 NAND3X1_16 ( .A(_163_), .B(_165_), .C(_164_), .Y(_166_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_160_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_161_) );
OAI21X1 OAI21X1_37 ( .A(_160_), .B(_161_), .C(w_cout_3_), .Y(_162_) );
NAND2X1 NAND2X1_41 ( .A(_162_), .B(_166_), .Y(_0__16_) );
OAI21X1 OAI21X1_38 ( .A(_163_), .B(_160_), .C(_165_), .Y(_11__1_) );
INVX1 INVX1_37 ( .A(_11__3_), .Y(_170_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_171_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_172_) );
NAND3X1 NAND3X1_17 ( .A(_170_), .B(_172_), .C(_171_), .Y(_173_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_167_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_168_) );
OAI21X1 OAI21X1_39 ( .A(_167_), .B(_168_), .C(_11__3_), .Y(_169_) );
NAND2X1 NAND2X1_43 ( .A(_169_), .B(_173_), .Y(_0__19_) );
OAI21X1 OAI21X1_40 ( .A(_170_), .B(_167_), .C(_172_), .Y(_10_) );
INVX1 INVX1_38 ( .A(_11__1_), .Y(_177_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_178_) );
NAND2X1 NAND2X1_44 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_179_) );
NAND3X1 NAND3X1_18 ( .A(_177_), .B(_179_), .C(_178_), .Y(_180_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_174_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_175_) );
OAI21X1 OAI21X1_41 ( .A(_174_), .B(_175_), .C(_11__1_), .Y(_176_) );
NAND2X1 NAND2X1_45 ( .A(_176_), .B(_180_), .Y(_0__17_) );
OAI21X1 OAI21X1_42 ( .A(_177_), .B(_174_), .C(_179_), .Y(_11__2_) );
INVX1 INVX1_39 ( .A(_11__2_), .Y(_184_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_185_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_186_) );
NAND3X1 NAND3X1_19 ( .A(_184_), .B(_186_), .C(_185_), .Y(_187_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_181_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_182_) );
OAI21X1 OAI21X1_43 ( .A(_181_), .B(_182_), .C(_11__2_), .Y(_183_) );
NAND2X1 NAND2X1_47 ( .A(_183_), .B(_187_), .Y(_0__18_) );
OAI21X1 OAI21X1_44 ( .A(_184_), .B(_181_), .C(_186_), .Y(_11__3_) );
INVX1 INVX1_40 ( .A(i_add_term1[16]), .Y(_188_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[16]), .B(_188_), .Y(_189_) );
INVX1 INVX1_41 ( .A(i_add_term2[16]), .Y(_190_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term1[16]), .B(_190_), .Y(_191_) );
INVX1 INVX1_42 ( .A(i_add_term1[17]), .Y(_192_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[17]), .B(_192_), .Y(_193_) );
INVX1 INVX1_43 ( .A(i_add_term2[17]), .Y(_194_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term1[17]), .B(_194_), .Y(_195_) );
OAI22X1 OAI22X1_5 ( .A(_189_), .B(_191_), .C(_193_), .D(_195_), .Y(_196_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_197_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_198_) );
NOR2X1 NOR2X1_53 ( .A(_197_), .B(_198_), .Y(_199_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_200_) );
NAND2X1 NAND2X1_48 ( .A(_199_), .B(_200_), .Y(_201_) );
NOR2X1 NOR2X1_54 ( .A(_196_), .B(_201_), .Y(_12_) );
INVX1 INVX1_44 ( .A(_10_), .Y(_202_) );
NAND2X1 NAND2X1_49 ( .A(gnd), .B(_12_), .Y(_203_) );
OAI21X1 OAI21X1_45 ( .A(_12_), .B(_202_), .C(_203_), .Y(w_cout_4_) );
INVX1 INVX1_45 ( .A(w_cout_4_), .Y(_207_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_208_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_209_) );
NAND3X1 NAND3X1_20 ( .A(_207_), .B(_209_), .C(_208_), .Y(_210_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_204_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_205_) );
OAI21X1 OAI21X1_46 ( .A(_204_), .B(_205_), .C(w_cout_4_), .Y(_206_) );
NAND2X1 NAND2X1_51 ( .A(_206_), .B(_210_), .Y(_0__20_) );
OAI21X1 OAI21X1_47 ( .A(_207_), .B(_204_), .C(_209_), .Y(_14__1_) );
INVX1 INVX1_46 ( .A(_14__3_), .Y(_214_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_215_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_216_) );
NAND3X1 NAND3X1_21 ( .A(_214_), .B(_216_), .C(_215_), .Y(_217_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_211_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_212_) );
OAI21X1 OAI21X1_48 ( .A(_211_), .B(_212_), .C(_14__3_), .Y(_213_) );
NAND2X1 NAND2X1_53 ( .A(_213_), .B(_217_), .Y(_0__23_) );
OAI21X1 OAI21X1_49 ( .A(_214_), .B(_211_), .C(_216_), .Y(_13_) );
INVX1 INVX1_47 ( .A(_14__1_), .Y(_221_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_222_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_223_) );
NAND3X1 NAND3X1_22 ( .A(_221_), .B(_223_), .C(_222_), .Y(_224_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_218_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_219_) );
OAI21X1 OAI21X1_50 ( .A(_218_), .B(_219_), .C(_14__1_), .Y(_220_) );
NAND2X1 NAND2X1_55 ( .A(_220_), .B(_224_), .Y(_0__21_) );
OAI21X1 OAI21X1_51 ( .A(_221_), .B(_218_), .C(_223_), .Y(_14__2_) );
INVX1 INVX1_48 ( .A(_14__2_), .Y(_228_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_229_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_230_) );
NAND3X1 NAND3X1_23 ( .A(_228_), .B(_230_), .C(_229_), .Y(_231_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_225_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_226_) );
OAI21X1 OAI21X1_52 ( .A(_225_), .B(_226_), .C(_14__2_), .Y(_227_) );
NAND2X1 NAND2X1_57 ( .A(_227_), .B(_231_), .Y(_0__22_) );
OAI21X1 OAI21X1_53 ( .A(_228_), .B(_225_), .C(_230_), .Y(_14__3_) );
INVX1 INVX1_49 ( .A(i_add_term1[20]), .Y(_232_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[20]), .B(_232_), .Y(_233_) );
INVX1 INVX1_50 ( .A(i_add_term2[20]), .Y(_234_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term1[20]), .B(_234_), .Y(_235_) );
INVX1 INVX1_51 ( .A(i_add_term1[21]), .Y(_236_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[21]), .B(_236_), .Y(_237_) );
INVX1 INVX1_52 ( .A(i_add_term2[21]), .Y(_238_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term1[21]), .B(_238_), .Y(_239_) );
OAI22X1 OAI22X1_6 ( .A(_233_), .B(_235_), .C(_237_), .D(_239_), .Y(_240_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_241_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_242_) );
NOR2X1 NOR2X1_64 ( .A(_241_), .B(_242_), .Y(_243_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_244_) );
NAND2X1 NAND2X1_58 ( .A(_243_), .B(_244_), .Y(_245_) );
NOR2X1 NOR2X1_65 ( .A(_240_), .B(_245_), .Y(_15_) );
INVX1 INVX1_53 ( .A(_13_), .Y(_246_) );
NAND2X1 NAND2X1_59 ( .A(gnd), .B(_15_), .Y(_247_) );
OAI21X1 OAI21X1_54 ( .A(_15_), .B(_246_), .C(_247_), .Y(w_cout_5_) );
INVX1 INVX1_54 ( .A(w_cout_5_), .Y(_251_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_252_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_253_) );
NAND3X1 NAND3X1_24 ( .A(_251_), .B(_253_), .C(_252_), .Y(_254_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_248_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_249_) );
OAI21X1 OAI21X1_55 ( .A(_248_), .B(_249_), .C(w_cout_5_), .Y(_250_) );
NAND2X1 NAND2X1_61 ( .A(_250_), .B(_254_), .Y(_0__24_) );
OAI21X1 OAI21X1_56 ( .A(_251_), .B(_248_), .C(_253_), .Y(_17__1_) );
INVX1 INVX1_55 ( .A(_17__3_), .Y(_258_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_259_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_260_) );
NAND3X1 NAND3X1_25 ( .A(_258_), .B(_260_), .C(_259_), .Y(_261_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_255_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_256_) );
OAI21X1 OAI21X1_57 ( .A(_255_), .B(_256_), .C(_17__3_), .Y(_257_) );
NAND2X1 NAND2X1_63 ( .A(_257_), .B(_261_), .Y(_0__27_) );
OAI21X1 OAI21X1_58 ( .A(_258_), .B(_255_), .C(_260_), .Y(_16_) );
INVX1 INVX1_56 ( .A(_17__1_), .Y(_265_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_266_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_267_) );
NAND3X1 NAND3X1_26 ( .A(_265_), .B(_267_), .C(_266_), .Y(_268_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_262_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_263_) );
OAI21X1 OAI21X1_59 ( .A(_262_), .B(_263_), .C(_17__1_), .Y(_264_) );
NAND2X1 NAND2X1_65 ( .A(_264_), .B(_268_), .Y(_0__25_) );
OAI21X1 OAI21X1_60 ( .A(_265_), .B(_262_), .C(_267_), .Y(_17__2_) );
INVX1 INVX1_57 ( .A(_17__2_), .Y(_272_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_273_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_274_) );
NAND3X1 NAND3X1_27 ( .A(_272_), .B(_274_), .C(_273_), .Y(_275_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_269_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_270_) );
OAI21X1 OAI21X1_61 ( .A(_269_), .B(_270_), .C(_17__2_), .Y(_271_) );
NAND2X1 NAND2X1_67 ( .A(_271_), .B(_275_), .Y(_0__26_) );
OAI21X1 OAI21X1_62 ( .A(_272_), .B(_269_), .C(_274_), .Y(_17__3_) );
INVX1 INVX1_58 ( .A(i_add_term1[24]), .Y(_276_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[24]), .B(_276_), .Y(_277_) );
INVX1 INVX1_59 ( .A(i_add_term2[24]), .Y(_278_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term1[24]), .B(_278_), .Y(_279_) );
INVX1 INVX1_60 ( .A(i_add_term1[25]), .Y(_280_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[25]), .B(_280_), .Y(_281_) );
INVX1 INVX1_61 ( .A(i_add_term2[25]), .Y(_282_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term1[25]), .B(_282_), .Y(_283_) );
OAI22X1 OAI22X1_7 ( .A(_277_), .B(_279_), .C(_281_), .D(_283_), .Y(_284_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_285_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_286_) );
NOR2X1 NOR2X1_75 ( .A(_285_), .B(_286_), .Y(_287_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_288_) );
NAND2X1 NAND2X1_68 ( .A(_287_), .B(_288_), .Y(_289_) );
NOR2X1 NOR2X1_76 ( .A(_284_), .B(_289_), .Y(_18_) );
INVX1 INVX1_62 ( .A(_16_), .Y(_290_) );
NAND2X1 NAND2X1_69 ( .A(gnd), .B(_18_), .Y(_291_) );
OAI21X1 OAI21X1_63 ( .A(_18_), .B(_290_), .C(_291_), .Y(w_cout_6_) );
INVX1 INVX1_63 ( .A(w_cout_6_), .Y(_295_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_296_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_297_) );
NAND3X1 NAND3X1_28 ( .A(_295_), .B(_297_), .C(_296_), .Y(_298_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_292_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_293_) );
OAI21X1 OAI21X1_64 ( .A(_292_), .B(_293_), .C(w_cout_6_), .Y(_294_) );
NAND2X1 NAND2X1_71 ( .A(_294_), .B(_298_), .Y(_0__28_) );
OAI21X1 OAI21X1_65 ( .A(_295_), .B(_292_), .C(_297_), .Y(_20__1_) );
INVX1 INVX1_64 ( .A(_20__3_), .Y(_302_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_303_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_304_) );
NAND3X1 NAND3X1_29 ( .A(_302_), .B(_304_), .C(_303_), .Y(_305_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_299_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_300_) );
OAI21X1 OAI21X1_66 ( .A(_299_), .B(_300_), .C(_20__3_), .Y(_301_) );
NAND2X1 NAND2X1_73 ( .A(_301_), .B(_305_), .Y(_0__31_) );
OAI21X1 OAI21X1_67 ( .A(_302_), .B(_299_), .C(_304_), .Y(_19_) );
INVX1 INVX1_65 ( .A(_20__1_), .Y(_309_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_310_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_311_) );
NAND3X1 NAND3X1_30 ( .A(_309_), .B(_311_), .C(_310_), .Y(_312_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_306_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_307_) );
OAI21X1 OAI21X1_68 ( .A(_306_), .B(_307_), .C(_20__1_), .Y(_308_) );
NAND2X1 NAND2X1_75 ( .A(_308_), .B(_312_), .Y(_0__29_) );
OAI21X1 OAI21X1_69 ( .A(_309_), .B(_306_), .C(_311_), .Y(_20__2_) );
INVX1 INVX1_66 ( .A(_20__2_), .Y(_316_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_317_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_318_) );
NAND3X1 NAND3X1_31 ( .A(_316_), .B(_318_), .C(_317_), .Y(_319_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_313_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_314_) );
OAI21X1 OAI21X1_70 ( .A(_313_), .B(_314_), .C(_20__2_), .Y(_315_) );
NAND2X1 NAND2X1_77 ( .A(_315_), .B(_319_), .Y(_0__30_) );
OAI21X1 OAI21X1_71 ( .A(_316_), .B(_313_), .C(_318_), .Y(_20__3_) );
INVX1 INVX1_67 ( .A(i_add_term1[28]), .Y(_320_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[28]), .B(_320_), .Y(_321_) );
INVX1 INVX1_68 ( .A(i_add_term2[28]), .Y(_322_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term1[28]), .B(_322_), .Y(_323_) );
INVX1 INVX1_69 ( .A(i_add_term1[29]), .Y(_324_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[29]), .B(_324_), .Y(_325_) );
INVX1 INVX1_70 ( .A(i_add_term2[29]), .Y(_326_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term1[29]), .B(_326_), .Y(_327_) );
OAI22X1 OAI22X1_8 ( .A(_321_), .B(_323_), .C(_325_), .D(_327_), .Y(_328_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_329_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_330_) );
NOR2X1 NOR2X1_86 ( .A(_329_), .B(_330_), .Y(_331_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_332_) );
NAND2X1 NAND2X1_78 ( .A(_331_), .B(_332_), .Y(_333_) );
NOR2X1 NOR2X1_87 ( .A(_328_), .B(_333_), .Y(_21_) );
INVX1 INVX1_71 ( .A(_19_), .Y(_334_) );
NAND2X1 NAND2X1_79 ( .A(gnd), .B(_21_), .Y(_335_) );
OAI21X1 OAI21X1_72 ( .A(_21_), .B(_334_), .C(_335_), .Y(w_cout_7_) );
INVX1 INVX1_72 ( .A(w_cout_7_), .Y(_339_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_340_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_341_) );
NAND3X1 NAND3X1_32 ( .A(_339_), .B(_341_), .C(_340_), .Y(_342_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_336_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_337_) );
OAI21X1 OAI21X1_73 ( .A(_336_), .B(_337_), .C(w_cout_7_), .Y(_338_) );
NAND2X1 NAND2X1_81 ( .A(_338_), .B(_342_), .Y(_0__32_) );
OAI21X1 OAI21X1_74 ( .A(_339_), .B(_336_), .C(_341_), .Y(_23__1_) );
INVX1 INVX1_73 ( .A(_23__3_), .Y(_346_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_347_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_348_) );
NAND3X1 NAND3X1_33 ( .A(_346_), .B(_348_), .C(_347_), .Y(_349_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_343_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_344_) );
OAI21X1 OAI21X1_75 ( .A(_343_), .B(_344_), .C(_23__3_), .Y(_345_) );
NAND2X1 NAND2X1_83 ( .A(_345_), .B(_349_), .Y(_0__35_) );
OAI21X1 OAI21X1_76 ( .A(_346_), .B(_343_), .C(_348_), .Y(_22_) );
INVX1 INVX1_74 ( .A(_23__1_), .Y(_353_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_354_) );
NAND2X1 NAND2X1_84 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_355_) );
NAND3X1 NAND3X1_34 ( .A(_353_), .B(_355_), .C(_354_), .Y(_356_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_350_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_351_) );
OAI21X1 OAI21X1_77 ( .A(_350_), .B(_351_), .C(_23__1_), .Y(_352_) );
NAND2X1 NAND2X1_85 ( .A(_352_), .B(_356_), .Y(_0__33_) );
OAI21X1 OAI21X1_78 ( .A(_353_), .B(_350_), .C(_355_), .Y(_23__2_) );
INVX1 INVX1_75 ( .A(_23__2_), .Y(_360_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_361_) );
NAND2X1 NAND2X1_86 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_362_) );
NAND3X1 NAND3X1_35 ( .A(_360_), .B(_362_), .C(_361_), .Y(_363_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_357_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_358_) );
OAI21X1 OAI21X1_79 ( .A(_357_), .B(_358_), .C(_23__2_), .Y(_359_) );
NAND2X1 NAND2X1_87 ( .A(_359_), .B(_363_), .Y(_0__34_) );
OAI21X1 OAI21X1_80 ( .A(_360_), .B(_357_), .C(_362_), .Y(_23__3_) );
INVX1 INVX1_76 ( .A(i_add_term1[32]), .Y(_364_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[32]), .B(_364_), .Y(_365_) );
INVX1 INVX1_77 ( .A(i_add_term2[32]), .Y(_366_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term1[32]), .B(_366_), .Y(_367_) );
INVX1 INVX1_78 ( .A(i_add_term1[33]), .Y(_368_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[33]), .B(_368_), .Y(_369_) );
INVX1 INVX1_79 ( .A(i_add_term2[33]), .Y(_370_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term1[33]), .B(_370_), .Y(_371_) );
OAI22X1 OAI22X1_9 ( .A(_365_), .B(_367_), .C(_369_), .D(_371_), .Y(_372_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_373_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_374_) );
NOR2X1 NOR2X1_97 ( .A(_373_), .B(_374_), .Y(_375_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_376_) );
NAND2X1 NAND2X1_88 ( .A(_375_), .B(_376_), .Y(_377_) );
NOR2X1 NOR2X1_98 ( .A(_372_), .B(_377_), .Y(_24_) );
INVX1 INVX1_80 ( .A(_22_), .Y(_378_) );
NAND2X1 NAND2X1_89 ( .A(gnd), .B(_24_), .Y(_379_) );
OAI21X1 OAI21X1_81 ( .A(_24_), .B(_378_), .C(_379_), .Y(w_cout_8_) );
INVX1 INVX1_81 ( .A(w_cout_8_), .Y(_383_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_384_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_385_) );
NAND3X1 NAND3X1_36 ( .A(_383_), .B(_385_), .C(_384_), .Y(_386_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_380_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_381_) );
OAI21X1 OAI21X1_82 ( .A(_380_), .B(_381_), .C(w_cout_8_), .Y(_382_) );
NAND2X1 NAND2X1_91 ( .A(_382_), .B(_386_), .Y(_0__36_) );
OAI21X1 OAI21X1_83 ( .A(_383_), .B(_380_), .C(_385_), .Y(_26__1_) );
INVX1 INVX1_82 ( .A(_26__3_), .Y(_390_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_391_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_392_) );
NAND3X1 NAND3X1_37 ( .A(_390_), .B(_392_), .C(_391_), .Y(_393_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_387_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_388_) );
OAI21X1 OAI21X1_84 ( .A(_387_), .B(_388_), .C(_26__3_), .Y(_389_) );
NAND2X1 NAND2X1_93 ( .A(_389_), .B(_393_), .Y(_0__39_) );
OAI21X1 OAI21X1_85 ( .A(_390_), .B(_387_), .C(_392_), .Y(_25_) );
INVX1 INVX1_83 ( .A(_26__1_), .Y(_397_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_398_) );
NAND2X1 NAND2X1_94 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_399_) );
NAND3X1 NAND3X1_38 ( .A(_397_), .B(_399_), .C(_398_), .Y(_400_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_394_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_395_) );
OAI21X1 OAI21X1_86 ( .A(_394_), .B(_395_), .C(_26__1_), .Y(_396_) );
NAND2X1 NAND2X1_95 ( .A(_396_), .B(_400_), .Y(_0__37_) );
OAI21X1 OAI21X1_87 ( .A(_397_), .B(_394_), .C(_399_), .Y(_26__2_) );
INVX1 INVX1_84 ( .A(_26__2_), .Y(_404_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_405_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_406_) );
NAND3X1 NAND3X1_39 ( .A(_404_), .B(_406_), .C(_405_), .Y(_407_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_401_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_402_) );
OAI21X1 OAI21X1_88 ( .A(_401_), .B(_402_), .C(_26__2_), .Y(_403_) );
NAND2X1 NAND2X1_97 ( .A(_403_), .B(_407_), .Y(_0__38_) );
OAI21X1 OAI21X1_89 ( .A(_404_), .B(_401_), .C(_406_), .Y(_26__3_) );
INVX1 INVX1_85 ( .A(i_add_term1[36]), .Y(_408_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[36]), .B(_408_), .Y(_409_) );
INVX1 INVX1_86 ( .A(i_add_term2[36]), .Y(_410_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term1[36]), .B(_410_), .Y(_411_) );
INVX1 INVX1_87 ( .A(i_add_term1[37]), .Y(_412_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[37]), .B(_412_), .Y(_413_) );
INVX1 INVX1_88 ( .A(i_add_term2[37]), .Y(_414_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term1[37]), .B(_414_), .Y(_415_) );
OAI22X1 OAI22X1_10 ( .A(_409_), .B(_411_), .C(_413_), .D(_415_), .Y(_416_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_417_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_418_) );
NOR2X1 NOR2X1_108 ( .A(_417_), .B(_418_), .Y(_419_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_420_) );
NAND2X1 NAND2X1_98 ( .A(_419_), .B(_420_), .Y(_421_) );
NOR2X1 NOR2X1_109 ( .A(_416_), .B(_421_), .Y(_27_) );
INVX1 INVX1_89 ( .A(_25_), .Y(_422_) );
NAND2X1 NAND2X1_99 ( .A(gnd), .B(_27_), .Y(_423_) );
OAI21X1 OAI21X1_90 ( .A(_27_), .B(_422_), .C(_423_), .Y(w_cout_9_) );
INVX1 INVX1_90 ( .A(gnd), .Y(_427_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_428_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_429_) );
NAND3X1 NAND3X1_40 ( .A(_427_), .B(_429_), .C(_428_), .Y(_430_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_424_) );
BUFX2 BUFX2_42 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_43 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_44 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_45 ( .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_46 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
