module cla_21bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add1[19], i_add1[20], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], i_add2[19], i_add2[20], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add1[19];
input i_add1[20];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
input i_add2[19];
input i_add2[20];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];

NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_74_) );
INVX1 INVX1_1 ( .A(_74_), .Y(w_C_1_) );
NAND2X1 NAND2X1_2 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_75_) );
NAND2X1 NAND2X1_3 ( .A(_74_), .B(_75_), .Y(_76_) );
OAI21X1 OAI21X1_1 ( .A(i_add2[1]), .B(i_add1[1]), .C(_76_), .Y(_77_) );
INVX1 INVX1_2 ( .A(_77_), .Y(w_C_2_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_78_) );
OR2X2 OR2X2_1 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_79_) );
OR2X2 OR2X2_2 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_80_) );
NAND3X1 NAND3X1_1 ( .A(_79_), .B(_80_), .C(_76_), .Y(_81_) );
NAND2X1 NAND2X1_5 ( .A(_78_), .B(_81_), .Y(w_C_3_) );
INVX1 INVX1_3 ( .A(i_add2[3]), .Y(_82_) );
INVX1 INVX1_4 ( .A(i_add1[3]), .Y(_83_) );
NAND2X1 NAND2X1_6 ( .A(_82_), .B(_83_), .Y(_84_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_85_) );
NAND3X1 NAND3X1_2 ( .A(_78_), .B(_85_), .C(_81_), .Y(_86_) );
AND2X2 AND2X2_1 ( .A(_86_), .B(_84_), .Y(w_C_4_) );
NAND2X1 NAND2X1_8 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_87_) );
OR2X2 OR2X2_3 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_88_) );
NAND3X1 NAND3X1_3 ( .A(_84_), .B(_88_), .C(_86_), .Y(_89_) );
NAND2X1 NAND2X1_9 ( .A(_87_), .B(_89_), .Y(w_C_5_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_90_) );
INVX1 INVX1_5 ( .A(_90_), .Y(_91_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_92_) );
NAND3X1 NAND3X1_4 ( .A(_87_), .B(_92_), .C(_89_), .Y(_93_) );
AND2X2 AND2X2_2 ( .A(_93_), .B(_91_), .Y(w_C_6_) );
INVX1 INVX1_6 ( .A(i_add2[6]), .Y(_94_) );
INVX1 INVX1_7 ( .A(i_add1[6]), .Y(_95_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_96_) );
INVX1 INVX1_8 ( .A(_96_), .Y(_97_) );
NAND3X1 NAND3X1_5 ( .A(_91_), .B(_97_), .C(_93_), .Y(_98_) );
OAI21X1 OAI21X1_2 ( .A(_94_), .B(_95_), .C(_98_), .Y(w_C_7_) );
NOR2X1 NOR2X1_3 ( .A(_94_), .B(_95_), .Y(_99_) );
INVX1 INVX1_9 ( .A(_99_), .Y(_100_) );
AND2X2 AND2X2_3 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_101_) );
INVX1 INVX1_10 ( .A(_101_), .Y(_102_) );
NAND3X1 NAND3X1_6 ( .A(_100_), .B(_102_), .C(_98_), .Y(_0_) );
OAI21X1 OAI21X1_3 ( .A(i_add2[7]), .B(i_add1[7]), .C(_0_), .Y(_1_) );
INVX1 INVX1_11 ( .A(_1_), .Y(w_C_8_) );
INVX1 INVX1_12 ( .A(i_add2[8]), .Y(_2_) );
INVX1 INVX1_13 ( .A(i_add1[8]), .Y(_3_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_4_) );
INVX1 INVX1_14 ( .A(_4_), .Y(_5_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_6_) );
INVX1 INVX1_15 ( .A(_6_), .Y(_7_) );
NAND3X1 NAND3X1_7 ( .A(_5_), .B(_7_), .C(_0_), .Y(_8_) );
OAI21X1 OAI21X1_4 ( .A(_2_), .B(_3_), .C(_8_), .Y(w_C_9_) );
NOR2X1 NOR2X1_6 ( .A(_2_), .B(_3_), .Y(_9_) );
INVX1 INVX1_16 ( .A(_9_), .Y(_10_) );
AND2X2 AND2X2_4 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_11_) );
INVX1 INVX1_17 ( .A(_11_), .Y(_12_) );
NAND3X1 NAND3X1_8 ( .A(_10_), .B(_12_), .C(_8_), .Y(_13_) );
OAI21X1 OAI21X1_5 ( .A(i_add2[9]), .B(i_add1[9]), .C(_13_), .Y(_14_) );
INVX1 INVX1_18 ( .A(_14_), .Y(w_C_10_) );
INVX1 INVX1_19 ( .A(i_add2[10]), .Y(_15_) );
INVX1 INVX1_20 ( .A(i_add1[10]), .Y(_16_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_17_) );
INVX1 INVX1_21 ( .A(_17_), .Y(_18_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_19_) );
INVX1 INVX1_22 ( .A(_19_), .Y(_20_) );
NAND3X1 NAND3X1_9 ( .A(_18_), .B(_20_), .C(_13_), .Y(_21_) );
OAI21X1 OAI21X1_6 ( .A(_15_), .B(_16_), .C(_21_), .Y(w_C_11_) );
NOR2X1 NOR2X1_9 ( .A(_15_), .B(_16_), .Y(_22_) );
INVX1 INVX1_23 ( .A(_22_), .Y(_23_) );
AND2X2 AND2X2_5 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_24_) );
INVX1 INVX1_24 ( .A(_24_), .Y(_25_) );
NAND3X1 NAND3X1_10 ( .A(_23_), .B(_25_), .C(_21_), .Y(_26_) );
OAI21X1 OAI21X1_7 ( .A(i_add2[11]), .B(i_add1[11]), .C(_26_), .Y(_27_) );
INVX1 INVX1_25 ( .A(_27_), .Y(w_C_12_) );
INVX1 INVX1_26 ( .A(i_add2[12]), .Y(_28_) );
INVX1 INVX1_27 ( .A(i_add1[12]), .Y(_29_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_30_) );
INVX1 INVX1_28 ( .A(_30_), .Y(_31_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_32_) );
INVX1 INVX1_29 ( .A(_32_), .Y(_33_) );
NAND3X1 NAND3X1_11 ( .A(_31_), .B(_33_), .C(_26_), .Y(_34_) );
OAI21X1 OAI21X1_8 ( .A(_28_), .B(_29_), .C(_34_), .Y(w_C_13_) );
NOR2X1 NOR2X1_12 ( .A(_28_), .B(_29_), .Y(_35_) );
INVX1 INVX1_30 ( .A(_35_), .Y(_36_) );
AND2X2 AND2X2_6 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_37_) );
INVX1 INVX1_31 ( .A(_37_), .Y(_38_) );
NAND3X1 NAND3X1_12 ( .A(_36_), .B(_38_), .C(_34_), .Y(_39_) );
OAI21X1 OAI21X1_9 ( .A(i_add2[13]), .B(i_add1[13]), .C(_39_), .Y(_40_) );
INVX1 INVX1_32 ( .A(_40_), .Y(w_C_14_) );
INVX1 INVX1_33 ( .A(i_add2[14]), .Y(_41_) );
INVX1 INVX1_34 ( .A(i_add1[14]), .Y(_42_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_43_) );
INVX1 INVX1_35 ( .A(_43_), .Y(_44_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_45_) );
INVX1 INVX1_36 ( .A(_45_), .Y(_46_) );
NAND3X1 NAND3X1_13 ( .A(_44_), .B(_46_), .C(_39_), .Y(_47_) );
OAI21X1 OAI21X1_10 ( .A(_41_), .B(_42_), .C(_47_), .Y(w_C_15_) );
NOR2X1 NOR2X1_15 ( .A(_41_), .B(_42_), .Y(_48_) );
INVX1 INVX1_37 ( .A(_48_), .Y(_49_) );
AND2X2 AND2X2_7 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_50_) );
INVX1 INVX1_38 ( .A(_50_), .Y(_51_) );
NAND3X1 NAND3X1_14 ( .A(_49_), .B(_51_), .C(_47_), .Y(_52_) );
OAI21X1 OAI21X1_11 ( .A(i_add2[15]), .B(i_add1[15]), .C(_52_), .Y(_53_) );
INVX1 INVX1_39 ( .A(_53_), .Y(w_C_16_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_54_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_55_) );
OAI21X1 OAI21X1_12 ( .A(_55_), .B(_53_), .C(_54_), .Y(w_C_17_) );
OR2X2 OR2X2_4 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_56_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_57_) );
INVX1 INVX1_40 ( .A(_57_), .Y(_58_) );
INVX1 INVX1_41 ( .A(_55_), .Y(_59_) );
NAND3X1 NAND3X1_15 ( .A(_58_), .B(_59_), .C(_52_), .Y(_60_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_61_) );
NAND3X1 NAND3X1_16 ( .A(_54_), .B(_61_), .C(_60_), .Y(_62_) );
AND2X2 AND2X2_8 ( .A(_62_), .B(_56_), .Y(w_C_18_) );
INVX1 INVX1_42 ( .A(i_add2[18]), .Y(_63_) );
INVX1 INVX1_43 ( .A(i_add1[18]), .Y(_64_) );
NAND2X1 NAND2X1_13 ( .A(_63_), .B(_64_), .Y(_65_) );
NAND3X1 NAND3X1_17 ( .A(_56_), .B(_65_), .C(_62_), .Y(_66_) );
OAI21X1 OAI21X1_13 ( .A(_63_), .B(_64_), .C(_66_), .Y(w_C_19_) );
OR2X2 OR2X2_5 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_67_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_68_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_69_) );
NAND3X1 NAND3X1_18 ( .A(_68_), .B(_69_), .C(_66_), .Y(_70_) );
AND2X2 AND2X2_9 ( .A(_70_), .B(_67_), .Y(w_C_20_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_71_) );
OR2X2 OR2X2_6 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_72_) );
NAND3X1 NAND3X1_19 ( .A(_67_), .B(_72_), .C(_70_), .Y(_73_) );
NAND2X1 NAND2X1_17 ( .A(_71_), .B(_73_), .Y(w_C_21_) );
BUFX2 BUFX2_1 ( .A(_103__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_103__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_103__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_103__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_103__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_103__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_103__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_103__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_103__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_103__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_103__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_103__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_103__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_103__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_103__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_103__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_103__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_103__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_103__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_103__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_103__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(w_C_21_), .Y(o_result[21]) );
INVX1 INVX1_44 ( .A(w_C_4_), .Y(_107_) );
OR2X2 OR2X2_7 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_108_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_109_) );
NAND3X1 NAND3X1_20 ( .A(_107_), .B(_109_), .C(_108_), .Y(_110_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_104_) );
AND2X2 AND2X2_10 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_105_) );
OAI21X1 OAI21X1_14 ( .A(_104_), .B(_105_), .C(w_C_4_), .Y(_106_) );
NAND2X1 NAND2X1_19 ( .A(_106_), .B(_110_), .Y(_103__4_) );
INVX1 INVX1_45 ( .A(w_C_5_), .Y(_114_) );
OR2X2 OR2X2_8 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_115_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_116_) );
NAND3X1 NAND3X1_21 ( .A(_114_), .B(_116_), .C(_115_), .Y(_117_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_111_) );
AND2X2 AND2X2_11 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_112_) );
OAI21X1 OAI21X1_15 ( .A(_111_), .B(_112_), .C(w_C_5_), .Y(_113_) );
NAND2X1 NAND2X1_21 ( .A(_113_), .B(_117_), .Y(_103__5_) );
INVX1 INVX1_46 ( .A(w_C_6_), .Y(_121_) );
OR2X2 OR2X2_9 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_122_) );
NAND2X1 NAND2X1_22 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_123_) );
NAND3X1 NAND3X1_22 ( .A(_121_), .B(_123_), .C(_122_), .Y(_124_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_118_) );
AND2X2 AND2X2_12 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_119_) );
OAI21X1 OAI21X1_16 ( .A(_118_), .B(_119_), .C(w_C_6_), .Y(_120_) );
NAND2X1 NAND2X1_23 ( .A(_120_), .B(_124_), .Y(_103__6_) );
INVX1 INVX1_47 ( .A(w_C_7_), .Y(_128_) );
OR2X2 OR2X2_10 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_129_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_130_) );
NAND3X1 NAND3X1_23 ( .A(_128_), .B(_130_), .C(_129_), .Y(_131_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_125_) );
AND2X2 AND2X2_13 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_126_) );
OAI21X1 OAI21X1_17 ( .A(_125_), .B(_126_), .C(w_C_7_), .Y(_127_) );
NAND2X1 NAND2X1_25 ( .A(_127_), .B(_131_), .Y(_103__7_) );
INVX1 INVX1_48 ( .A(w_C_8_), .Y(_135_) );
OR2X2 OR2X2_11 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_136_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_137_) );
NAND3X1 NAND3X1_24 ( .A(_135_), .B(_137_), .C(_136_), .Y(_138_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_132_) );
AND2X2 AND2X2_14 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_133_) );
OAI21X1 OAI21X1_18 ( .A(_132_), .B(_133_), .C(w_C_8_), .Y(_134_) );
NAND2X1 NAND2X1_27 ( .A(_134_), .B(_138_), .Y(_103__8_) );
INVX1 INVX1_49 ( .A(w_C_9_), .Y(_142_) );
OR2X2 OR2X2_12 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_143_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_144_) );
NAND3X1 NAND3X1_25 ( .A(_142_), .B(_144_), .C(_143_), .Y(_145_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_139_) );
AND2X2 AND2X2_15 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_140_) );
OAI21X1 OAI21X1_19 ( .A(_139_), .B(_140_), .C(w_C_9_), .Y(_141_) );
NAND2X1 NAND2X1_29 ( .A(_141_), .B(_145_), .Y(_103__9_) );
INVX1 INVX1_50 ( .A(w_C_10_), .Y(_149_) );
OR2X2 OR2X2_13 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_150_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_151_) );
NAND3X1 NAND3X1_26 ( .A(_149_), .B(_151_), .C(_150_), .Y(_152_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_146_) );
AND2X2 AND2X2_16 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_147_) );
OAI21X1 OAI21X1_20 ( .A(_146_), .B(_147_), .C(w_C_10_), .Y(_148_) );
NAND2X1 NAND2X1_31 ( .A(_148_), .B(_152_), .Y(_103__10_) );
INVX1 INVX1_51 ( .A(w_C_11_), .Y(_156_) );
OR2X2 OR2X2_14 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_157_) );
NAND2X1 NAND2X1_32 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_158_) );
NAND3X1 NAND3X1_27 ( .A(_156_), .B(_158_), .C(_157_), .Y(_159_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_153_) );
AND2X2 AND2X2_17 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_154_) );
OAI21X1 OAI21X1_21 ( .A(_153_), .B(_154_), .C(w_C_11_), .Y(_155_) );
NAND2X1 NAND2X1_33 ( .A(_155_), .B(_159_), .Y(_103__11_) );
INVX1 INVX1_52 ( .A(w_C_12_), .Y(_163_) );
OR2X2 OR2X2_15 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_164_) );
NAND2X1 NAND2X1_34 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_165_) );
NAND3X1 NAND3X1_28 ( .A(_163_), .B(_165_), .C(_164_), .Y(_166_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_160_) );
AND2X2 AND2X2_18 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_161_) );
OAI21X1 OAI21X1_22 ( .A(_160_), .B(_161_), .C(w_C_12_), .Y(_162_) );
NAND2X1 NAND2X1_35 ( .A(_162_), .B(_166_), .Y(_103__12_) );
INVX1 INVX1_53 ( .A(w_C_13_), .Y(_170_) );
OR2X2 OR2X2_16 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_171_) );
NAND2X1 NAND2X1_36 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_172_) );
NAND3X1 NAND3X1_29 ( .A(_170_), .B(_172_), .C(_171_), .Y(_173_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_167_) );
AND2X2 AND2X2_19 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_168_) );
OAI21X1 OAI21X1_23 ( .A(_167_), .B(_168_), .C(w_C_13_), .Y(_169_) );
NAND2X1 NAND2X1_37 ( .A(_169_), .B(_173_), .Y(_103__13_) );
INVX1 INVX1_54 ( .A(w_C_14_), .Y(_177_) );
OR2X2 OR2X2_17 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_178_) );
NAND2X1 NAND2X1_38 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_179_) );
NAND3X1 NAND3X1_30 ( .A(_177_), .B(_179_), .C(_178_), .Y(_180_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_174_) );
AND2X2 AND2X2_20 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_175_) );
OAI21X1 OAI21X1_24 ( .A(_174_), .B(_175_), .C(w_C_14_), .Y(_176_) );
NAND2X1 NAND2X1_39 ( .A(_176_), .B(_180_), .Y(_103__14_) );
INVX1 INVX1_55 ( .A(w_C_15_), .Y(_184_) );
OR2X2 OR2X2_18 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_185_) );
NAND2X1 NAND2X1_40 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_186_) );
NAND3X1 NAND3X1_31 ( .A(_184_), .B(_186_), .C(_185_), .Y(_187_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_181_) );
AND2X2 AND2X2_21 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_182_) );
OAI21X1 OAI21X1_25 ( .A(_181_), .B(_182_), .C(w_C_15_), .Y(_183_) );
NAND2X1 NAND2X1_41 ( .A(_183_), .B(_187_), .Y(_103__15_) );
INVX1 INVX1_56 ( .A(w_C_16_), .Y(_191_) );
OR2X2 OR2X2_19 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_192_) );
NAND2X1 NAND2X1_42 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_193_) );
NAND3X1 NAND3X1_32 ( .A(_191_), .B(_193_), .C(_192_), .Y(_194_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_188_) );
AND2X2 AND2X2_22 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_189_) );
OAI21X1 OAI21X1_26 ( .A(_188_), .B(_189_), .C(w_C_16_), .Y(_190_) );
NAND2X1 NAND2X1_43 ( .A(_190_), .B(_194_), .Y(_103__16_) );
INVX1 INVX1_57 ( .A(w_C_17_), .Y(_198_) );
OR2X2 OR2X2_20 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_199_) );
NAND2X1 NAND2X1_44 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_200_) );
NAND3X1 NAND3X1_33 ( .A(_198_), .B(_200_), .C(_199_), .Y(_201_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_195_) );
AND2X2 AND2X2_23 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_196_) );
OAI21X1 OAI21X1_27 ( .A(_195_), .B(_196_), .C(w_C_17_), .Y(_197_) );
NAND2X1 NAND2X1_45 ( .A(_197_), .B(_201_), .Y(_103__17_) );
INVX1 INVX1_58 ( .A(w_C_18_), .Y(_205_) );
OR2X2 OR2X2_21 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_206_) );
NAND2X1 NAND2X1_46 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_207_) );
NAND3X1 NAND3X1_34 ( .A(_205_), .B(_207_), .C(_206_), .Y(_208_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_202_) );
AND2X2 AND2X2_24 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_203_) );
OAI21X1 OAI21X1_28 ( .A(_202_), .B(_203_), .C(w_C_18_), .Y(_204_) );
NAND2X1 NAND2X1_47 ( .A(_204_), .B(_208_), .Y(_103__18_) );
INVX1 INVX1_59 ( .A(w_C_19_), .Y(_212_) );
OR2X2 OR2X2_22 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_213_) );
NAND2X1 NAND2X1_48 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_214_) );
NAND3X1 NAND3X1_35 ( .A(_212_), .B(_214_), .C(_213_), .Y(_215_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_209_) );
AND2X2 AND2X2_25 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_210_) );
OAI21X1 OAI21X1_29 ( .A(_209_), .B(_210_), .C(w_C_19_), .Y(_211_) );
NAND2X1 NAND2X1_49 ( .A(_211_), .B(_215_), .Y(_103__19_) );
INVX1 INVX1_60 ( .A(w_C_20_), .Y(_219_) );
OR2X2 OR2X2_23 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_220_) );
NAND2X1 NAND2X1_50 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_221_) );
NAND3X1 NAND3X1_36 ( .A(_219_), .B(_221_), .C(_220_), .Y(_222_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_216_) );
AND2X2 AND2X2_26 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_217_) );
OAI21X1 OAI21X1_30 ( .A(_216_), .B(_217_), .C(w_C_20_), .Y(_218_) );
NAND2X1 NAND2X1_51 ( .A(_218_), .B(_222_), .Y(_103__20_) );
INVX1 INVX1_61 ( .A(1'b0), .Y(_226_) );
OR2X2 OR2X2_24 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_227_) );
NAND2X1 NAND2X1_52 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_228_) );
NAND3X1 NAND3X1_37 ( .A(_226_), .B(_228_), .C(_227_), .Y(_229_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_223_) );
AND2X2 AND2X2_27 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_224_) );
OAI21X1 OAI21X1_31 ( .A(_223_), .B(_224_), .C(1'b0), .Y(_225_) );
NAND2X1 NAND2X1_53 ( .A(_225_), .B(_229_), .Y(_103__0_) );
INVX1 INVX1_62 ( .A(w_C_1_), .Y(_233_) );
OR2X2 OR2X2_25 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_234_) );
NAND2X1 NAND2X1_54 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_235_) );
NAND3X1 NAND3X1_38 ( .A(_233_), .B(_235_), .C(_234_), .Y(_236_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_230_) );
AND2X2 AND2X2_28 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_231_) );
OAI21X1 OAI21X1_32 ( .A(_230_), .B(_231_), .C(w_C_1_), .Y(_232_) );
NAND2X1 NAND2X1_55 ( .A(_232_), .B(_236_), .Y(_103__1_) );
INVX1 INVX1_63 ( .A(w_C_2_), .Y(_240_) );
OR2X2 OR2X2_26 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_241_) );
NAND2X1 NAND2X1_56 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_242_) );
NAND3X1 NAND3X1_39 ( .A(_240_), .B(_242_), .C(_241_), .Y(_243_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_237_) );
AND2X2 AND2X2_29 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_238_) );
OAI21X1 OAI21X1_33 ( .A(_237_), .B(_238_), .C(w_C_2_), .Y(_239_) );
NAND2X1 NAND2X1_57 ( .A(_239_), .B(_243_), .Y(_103__2_) );
INVX1 INVX1_64 ( .A(w_C_3_), .Y(_247_) );
OR2X2 OR2X2_27 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_248_) );
NAND2X1 NAND2X1_58 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_249_) );
NAND3X1 NAND3X1_40 ( .A(_247_), .B(_249_), .C(_248_), .Y(_250_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_244_) );
AND2X2 AND2X2_30 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_245_) );
OAI21X1 OAI21X1_34 ( .A(_244_), .B(_245_), .C(w_C_3_), .Y(_246_) );
NAND2X1 NAND2X1_59 ( .A(_246_), .B(_250_), .Y(_103__3_) );
BUFX2 BUFX2_23 ( .A(w_C_21_), .Y(_103__21_) );
BUFX2 BUFX2_24 ( .A(1'b0), .Y(w_C_0_) );
endmodule
