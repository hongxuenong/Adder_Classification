module cla_44bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [43:0] i_add1;
input [43:0] i_add2;
output [44:0] o_result;

INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(w_C_16_), .Y(_341_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_342_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_343_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_343_), .C(_342_), .Y(_344_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_338_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_339_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_339_), .C(w_C_16_), .Y(_340_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_344_), .Y(_253__16_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(w_C_17_), .Y(_348_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_349_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_350_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_350_), .C(_349_), .Y(_351_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_345_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_346_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_346_), .C(w_C_17_), .Y(_347_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_351_), .Y(_253__17_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(w_C_18_), .Y(_355_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_356_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_357_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_357_), .C(_356_), .Y(_358_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_352_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_353_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_353_), .C(w_C_18_), .Y(_354_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_358_), .Y(_253__18_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(w_C_19_), .Y(_362_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_363_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_364_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_364_), .C(_363_), .Y(_365_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_359_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_360_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_360_), .C(w_C_19_), .Y(_361_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_365_), .Y(_253__19_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(w_C_20_), .Y(_369_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_370_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_371_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_371_), .C(_370_), .Y(_372_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_366_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_367_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_367_), .C(w_C_20_), .Y(_368_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_372_), .Y(_253__20_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(w_C_21_), .Y(_376_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_377_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_378_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_378_), .C(_377_), .Y(_379_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_373_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_374_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_373_), .B(_374_), .C(w_C_21_), .Y(_375_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_379_), .Y(_253__21_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(w_C_22_), .Y(_383_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_384_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_385_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_385_), .C(_384_), .Y(_386_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_380_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_381_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_381_), .C(w_C_22_), .Y(_382_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_382_), .B(_386_), .Y(_253__22_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(w_C_23_), .Y(_390_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_391_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_392_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_392_), .C(_391_), .Y(_393_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_387_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_388_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_388_), .C(w_C_23_), .Y(_389_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_393_), .Y(_253__23_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(w_C_24_), .Y(_397_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_398_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_399_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_399_), .C(_398_), .Y(_400_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_394_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_395_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_395_), .C(w_C_24_), .Y(_396_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_400_), .Y(_253__24_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(w_C_25_), .Y(_404_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_405_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_406_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_406_), .C(_405_), .Y(_407_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_401_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_402_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_402_), .C(w_C_25_), .Y(_403_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_407_), .Y(_253__25_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(w_C_26_), .Y(_411_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_412_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_413_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_413_), .C(_412_), .Y(_414_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_408_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_409_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_409_), .C(w_C_26_), .Y(_410_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(_414_), .Y(_253__26_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(w_C_27_), .Y(_418_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_419_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_420_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_420_), .C(_419_), .Y(_421_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_415_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_416_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_415_), .B(_416_), .C(w_C_27_), .Y(_417_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_421_), .Y(_253__27_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(w_C_28_), .Y(_425_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_426_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_427_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(_427_), .C(_426_), .Y(_428_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_422_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_423_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_422_), .B(_423_), .C(w_C_28_), .Y(_424_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_428_), .Y(_253__28_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(w_C_29_), .Y(_432_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_433_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_434_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_432_), .B(_434_), .C(_433_), .Y(_435_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_429_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_430_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(_430_), .C(w_C_29_), .Y(_431_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_435_), .Y(_253__29_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(w_C_30_), .Y(_439_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_440_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_441_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_441_), .C(_440_), .Y(_442_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_436_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_437_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_437_), .C(w_C_30_), .Y(_438_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_442_), .Y(_253__30_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(w_C_31_), .Y(_446_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_447_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_448_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(_448_), .C(_447_), .Y(_449_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_443_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_444_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_444_), .C(w_C_31_), .Y(_445_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_445_), .B(_449_), .Y(_253__31_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(w_C_32_), .Y(_453_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_454_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_455_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(_455_), .C(_454_), .Y(_456_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_450_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_451_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_451_), .C(w_C_32_), .Y(_452_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_456_), .Y(_253__32_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(w_C_33_), .Y(_460_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_461_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_462_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_462_), .C(_461_), .Y(_463_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_457_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_458_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_458_), .C(w_C_33_), .Y(_459_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_459_), .B(_463_), .Y(_253__33_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(w_C_34_), .Y(_467_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_468_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_469_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_467_), .B(_469_), .C(_468_), .Y(_470_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_464_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_465_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_465_), .C(w_C_34_), .Y(_466_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_466_), .B(_470_), .Y(_253__34_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(w_C_35_), .Y(_474_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_475_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_476_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_474_), .B(_476_), .C(_475_), .Y(_477_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_471_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_472_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_472_), .C(w_C_35_), .Y(_473_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_477_), .Y(_253__35_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(w_C_36_), .Y(_481_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_482_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_483_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_483_), .C(_482_), .Y(_484_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_478_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_479_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_479_), .C(w_C_36_), .Y(_480_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_484_), .Y(_253__36_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(w_C_37_), .Y(_488_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_489_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_490_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_490_), .C(_489_), .Y(_491_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_485_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_486_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_486_), .C(w_C_37_), .Y(_487_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_491_), .Y(_253__37_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(w_C_38_), .Y(_495_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_496_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_497_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_495_), .B(_497_), .C(_496_), .Y(_498_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_492_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_493_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_492_), .B(_493_), .C(w_C_38_), .Y(_494_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_498_), .Y(_253__38_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(w_C_39_), .Y(_502_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_503_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_504_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_502_), .B(_504_), .C(_503_), .Y(_505_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_499_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_500_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_500_), .C(w_C_39_), .Y(_501_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_501_), .B(_505_), .Y(_253__39_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(w_C_40_), .Y(_509_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_510_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_511_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_511_), .C(_510_), .Y(_512_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_506_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_507_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_507_), .C(w_C_40_), .Y(_508_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_512_), .Y(_253__40_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(w_C_41_), .Y(_516_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_517_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_518_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_518_), .C(_517_), .Y(_519_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_513_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_514_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_514_), .C(w_C_41_), .Y(_515_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_519_), .Y(_253__41_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(w_C_42_), .Y(_523_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_524_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_525_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_525_), .C(_524_), .Y(_526_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_520_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_521_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_521_), .C(w_C_42_), .Y(_522_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_522_), .B(_526_), .Y(_253__42_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(w_C_43_), .Y(_530_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_531_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_532_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_532_), .C(_531_), .Y(_533_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_527_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_528_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_528_), .C(w_C_43_), .Y(_529_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_533_), .Y(_253__43_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_537_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_538_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_539_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_539_), .C(_538_), .Y(_540_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_534_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_535_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_535_), .C(gnd), .Y(_536_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_536_), .B(_540_), .Y(_253__0_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_544_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_545_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_546_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_546_), .C(_545_), .Y(_547_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_541_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_542_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_541_), .B(_542_), .C(w_C_1_), .Y(_543_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_547_), .Y(_253__1_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_551_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_552_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_553_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_551_), .B(_553_), .C(_552_), .Y(_554_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_548_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_549_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_549_), .C(w_C_2_), .Y(_550_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_550_), .B(_554_), .Y(_253__2_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_558_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_559_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_560_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_560_), .C(_559_), .Y(_561_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_555_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_556_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_555_), .B(_556_), .C(w_C_3_), .Y(_557_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_557_), .B(_561_), .Y(_253__3_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_2_), .Y(w_C_2_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .Y(_3_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add1[2]), .Y(_4_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_2_), .C(_6_), .Y(_7_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_9_), .C(_7_), .Y(_10_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_8_), .Y(_11_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(w_C_4_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_12_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_11_), .C(_12_), .Y(w_C_5_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_14_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_14_), .Y(_15_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_16_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_12_), .C(_10_), .Y(_17_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_18_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_18_), .Y(_19_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_19_), .C(_17_), .Y(_20_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_15_), .Y(_21_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_21_), .Y(w_C_6_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_23_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_23_), .C(_20_), .Y(_24_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .C(_24_), .Y(_25_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(w_C_7_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .Y(_26_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add1[7]), .Y(_27_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_28_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_28_), .Y(_29_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_30_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_31_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_31_), .C(_24_), .Y(_32_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_27_), .C(_32_), .Y(w_C_8_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_27_), .Y(_33_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_33_), .Y(_34_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_35_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_35_), .Y(_36_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_36_), .C(_32_), .Y(_37_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .C(_37_), .Y(_38_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_38_), .Y(w_C_9_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .Y(_39_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add1[9]), .Y(_40_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_41_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_41_), .Y(_42_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_43_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(_44_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_44_), .C(_37_), .Y(_45_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_40_), .C(_45_), .Y(w_C_10_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_40_), .Y(_46_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_46_), .Y(_47_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_48_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_48_), .Y(_49_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_49_), .C(_45_), .Y(_50_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .C(_50_), .Y(_51_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_51_), .Y(w_C_11_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .Y(_52_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add1[11]), .Y(_53_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_54_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_54_), .Y(_55_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_56_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_56_), .Y(_57_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_57_), .C(_50_), .Y(_58_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_53_), .C(_58_), .Y(w_C_12_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_53_), .Y(_59_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_59_), .Y(_60_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_61_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_61_), .Y(_62_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_62_), .C(_58_), .Y(_63_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .C(_63_), .Y(_64_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_64_), .Y(w_C_13_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .Y(_65_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add1[13]), .Y(_66_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_67_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_67_), .Y(_68_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_69_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(_70_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_70_), .C(_63_), .Y(_71_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_66_), .C(_71_), .Y(w_C_14_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_66_), .Y(_72_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_72_), .Y(_73_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_74_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_74_), .Y(_75_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_75_), .C(_71_), .Y(_76_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .C(_76_), .Y(_77_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_77_), .Y(w_C_15_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .Y(_78_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add1[15]), .Y(_79_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_80_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(_80_), .Y(_81_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_82_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_82_), .Y(_83_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_83_), .C(_76_), .Y(_84_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_79_), .C(_84_), .Y(w_C_16_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_79_), .Y(_85_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_85_), .Y(_86_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_87_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_87_), .Y(_88_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_88_), .C(_84_), .Y(_89_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .C(_89_), .Y(_90_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_90_), .Y(w_C_17_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .Y(_91_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add1[17]), .Y(_92_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_93_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_93_), .Y(_94_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_95_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_95_), .Y(_96_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_96_), .C(_89_), .Y(_97_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_92_), .C(_97_), .Y(w_C_18_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_92_), .Y(_98_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_98_), .Y(_99_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_100_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_100_), .Y(_101_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_101_), .C(_97_), .Y(_102_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .C(_102_), .Y(_103_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(_103_), .Y(w_C_19_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .Y(_104_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add1[19]), .Y(_105_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_106_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(_106_), .Y(_107_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_108_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(_108_), .Y(_109_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_109_), .C(_102_), .Y(_110_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_105_), .C(_110_), .Y(w_C_20_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_105_), .Y(_111_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(_111_), .Y(_112_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_113_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_113_), .Y(_114_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_114_), .C(_110_), .Y(_115_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .C(_115_), .Y(_116_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(_116_), .Y(w_C_21_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .Y(_117_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add1[21]), .Y(_118_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_119_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_119_), .Y(_120_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_121_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_121_), .Y(_122_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_122_), .C(_115_), .Y(_123_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_118_), .C(_123_), .Y(w_C_22_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_118_), .Y(_124_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(_124_), .Y(_125_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_126_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(_126_), .Y(_127_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_127_), .C(_123_), .Y(_128_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .C(_128_), .Y(_129_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(_129_), .Y(w_C_23_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .Y(_130_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add1[23]), .Y(_131_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_132_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(_132_), .Y(_133_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_134_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(_134_), .Y(_135_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_135_), .C(_128_), .Y(_136_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_131_), .C(_136_), .Y(w_C_24_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_131_), .Y(_137_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_137_), .Y(_138_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_139_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(_139_), .Y(_140_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_140_), .C(_136_), .Y(_141_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .C(_141_), .Y(_142_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_142_), .Y(w_C_25_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .Y(_143_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add1[25]), .Y(_144_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_145_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_145_), .Y(_146_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_147_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_147_), .Y(_148_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_148_), .C(_141_), .Y(_149_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_144_), .C(_149_), .Y(w_C_26_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_144_), .Y(_150_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(_150_), .Y(_151_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_152_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_152_), .Y(_153_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_153_), .C(_149_), .Y(_154_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .C(_154_), .Y(_155_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(w_C_27_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .Y(_156_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(i_add1[27]), .Y(_157_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_158_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(_158_), .Y(_159_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_160_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(_160_), .Y(_161_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_159_), .B(_161_), .C(_154_), .Y(_162_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_157_), .C(_162_), .Y(w_C_28_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_157_), .Y(_163_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(_163_), .Y(_164_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_165_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(_165_), .Y(_166_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_166_), .C(_162_), .Y(_167_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .C(_167_), .Y(_168_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(_168_), .Y(w_C_29_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .Y(_169_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(i_add1[29]), .Y(_170_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_171_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(_171_), .Y(_172_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_173_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(_173_), .Y(_174_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_174_), .C(_167_), .Y(_175_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_170_), .C(_175_), .Y(w_C_30_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_170_), .Y(_176_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(_176_), .Y(_177_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_178_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(_178_), .Y(_179_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_179_), .C(_175_), .Y(_180_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .C(_180_), .Y(_181_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(_181_), .Y(w_C_31_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .Y(_182_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(i_add1[31]), .Y(_183_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_184_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(_184_), .Y(_185_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_186_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(_186_), .Y(_187_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_187_), .C(_180_), .Y(_188_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_183_), .C(_188_), .Y(w_C_32_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_183_), .Y(_189_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(_189_), .Y(_190_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_191_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(_191_), .Y(_192_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_192_), .C(_188_), .Y(_193_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .C(_193_), .Y(_194_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(_194_), .Y(w_C_33_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .Y(_195_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(i_add1[33]), .Y(_196_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_197_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(_197_), .Y(_198_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_199_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(_199_), .Y(_200_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_200_), .C(_193_), .Y(_201_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_196_), .C(_201_), .Y(w_C_34_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_202_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(_202_), .Y(_203_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_196_), .Y(_204_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(_204_), .Y(_205_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_206_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_206_), .C(_201_), .Y(_207_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_203_), .Y(w_C_35_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .Y(_208_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(i_add1[35]), .Y(_209_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_209_), .Y(_210_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_210_), .C(_207_), .Y(_211_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_209_), .C(_211_), .Y(w_C_36_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .Y(_212_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(i_add1[36]), .Y(_213_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .C(w_C_36_), .Y(_214_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_213_), .C(_214_), .Y(w_C_37_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .Y(_215_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(i_add1[37]), .Y(_216_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_216_), .Y(_217_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(w_C_37_), .B(_217_), .Y(_218_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .C(_218_), .Y(_219_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(_219_), .Y(w_C_38_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(_217_), .Y(_220_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_213_), .Y(_221_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_222_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_223_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_223_), .C(_211_), .Y(_224_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_216_), .Y(_225_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_225_), .C(_224_), .Y(_226_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_227_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_227_), .C(_226_), .Y(_228_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .C(_228_), .Y(_229_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(_229_), .Y(w_C_39_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .Y(_230_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(i_add1[39]), .Y(_231_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_231_), .C(_229_), .Y(_232_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .C(_232_), .Y(_233_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(_233_), .Y(w_C_40_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_234_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[40]), .B(i_add1[40]), .Y(_235_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_233_), .C(_234_), .Y(w_C_41_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_236_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(_235_), .Y(_237_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_231_), .Y(_238_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(_238_), .Y(_239_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_240_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(_240_), .Y(_241_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_231_), .Y(_242_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_242_), .C(_228_), .Y(_243_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_234_), .C(_243_), .Y(_244_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[41]), .B(i_add1[41]), .Y(_245_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_245_), .C(_244_), .Y(_246_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_246_), .Y(w_C_42_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_247_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[42]), .B(i_add1[42]), .Y(_248_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_248_), .C(_246_), .Y(_249_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_247_), .Y(w_C_43_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_250_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[43]), .B(i_add1[43]), .Y(_251_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_251_), .C(_249_), .Y(_252_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_252_), .Y(w_C_44_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_253__2_), .Y(o_result[2]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_253__3_), .Y(o_result[3]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_253__4_), .Y(o_result[4]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_253__5_), .Y(o_result[5]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_253__6_), .Y(o_result[6]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_253__7_), .Y(o_result[7]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_253__8_), .Y(o_result[8]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_253__9_), .Y(o_result[9]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_253__10_), .Y(o_result[10]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_253__11_), .Y(o_result[11]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_253__12_), .Y(o_result[12]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_253__13_), .Y(o_result[13]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_253__14_), .Y(o_result[14]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_253__15_), .Y(o_result[15]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_253__16_), .Y(o_result[16]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_253__17_), .Y(o_result[17]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_253__18_), .Y(o_result[18]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_253__19_), .Y(o_result[19]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_253__20_), .Y(o_result[20]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_253__21_), .Y(o_result[21]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_253__22_), .Y(o_result[22]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_253__23_), .Y(o_result[23]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_253__24_), .Y(o_result[24]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_253__25_), .Y(o_result[25]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_253__26_), .Y(o_result[26]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_253__27_), .Y(o_result[27]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_253__28_), .Y(o_result[28]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_253__29_), .Y(o_result[29]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_253__30_), .Y(o_result[30]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_253__31_), .Y(o_result[31]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_253__32_), .Y(o_result[32]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_253__33_), .Y(o_result[33]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_253__34_), .Y(o_result[34]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_253__35_), .Y(o_result[35]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_253__36_), .Y(o_result[36]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_253__37_), .Y(o_result[37]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_253__38_), .Y(o_result[38]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_253__39_), .Y(o_result[39]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_253__40_), .Y(o_result[40]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_253__41_), .Y(o_result[41]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_253__42_), .Y(o_result[42]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_253__43_), .Y(o_result[43]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(w_C_44_), .Y(o_result[44]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_253__0_), .Y(o_result[0]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_253__1_), .Y(o_result[1]) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_257_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_258_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_259_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_259_), .C(_258_), .Y(_260_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_254_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_255_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_255_), .C(w_C_4_), .Y(_256_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_260_), .Y(_253__4_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_264_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_265_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_266_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_266_), .C(_265_), .Y(_267_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_261_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_262_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_262_), .C(w_C_5_), .Y(_263_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_267_), .Y(_253__5_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_271_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_272_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_273_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_273_), .C(_272_), .Y(_274_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_268_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_269_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_269_), .C(w_C_6_), .Y(_270_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_274_), .Y(_253__6_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_278_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_279_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_280_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_280_), .C(_279_), .Y(_281_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_275_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_276_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_276_), .C(w_C_7_), .Y(_277_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_281_), .Y(_253__7_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_285_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_286_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_287_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_287_), .C(_286_), .Y(_288_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_282_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_283_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_283_), .C(w_C_8_), .Y(_284_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_288_), .Y(_253__8_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_292_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_293_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_294_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_292_), .B(_294_), .C(_293_), .Y(_295_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_289_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_290_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_290_), .C(w_C_9_), .Y(_291_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_295_), .Y(_253__9_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_299_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_300_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_301_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_301_), .C(_300_), .Y(_302_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_296_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_297_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_297_), .C(w_C_10_), .Y(_298_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_302_), .Y(_253__10_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_306_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_307_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_308_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_308_), .C(_307_), .Y(_309_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_303_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_304_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_304_), .C(w_C_11_), .Y(_305_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_309_), .Y(_253__11_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(w_C_12_), .Y(_313_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_314_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_315_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_315_), .C(_314_), .Y(_316_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_310_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_311_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_311_), .C(w_C_12_), .Y(_312_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_316_), .Y(_253__12_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(w_C_13_), .Y(_320_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_321_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_322_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_322_), .C(_321_), .Y(_323_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_317_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_318_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_318_), .C(w_C_13_), .Y(_319_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_323_), .Y(_253__13_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(w_C_14_), .Y(_327_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_328_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_329_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_329_), .C(_328_), .Y(_330_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_324_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_325_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_325_), .C(w_C_14_), .Y(_326_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_330_), .Y(_253__14_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(_334_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_335_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_336_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_336_), .C(_335_), .Y(_337_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_331_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_332_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_332_), .C(w_C_15_), .Y(_333_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_337_), .Y(_253__15_) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(w_C_44_), .Y(_253__44_) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
