module cla_58bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add1[19], i_add1[20], i_add1[21], i_add1[22], i_add1[23], i_add1[24], i_add1[25], i_add1[26], i_add1[27], i_add1[28], i_add1[29], i_add1[30], i_add1[31], i_add1[32], i_add1[33], i_add1[34], i_add1[35], i_add1[36], i_add1[37], i_add1[38], i_add1[39], i_add1[40], i_add1[41], i_add1[42], i_add1[43], i_add1[44], i_add1[45], i_add1[46], i_add1[47], i_add1[48], i_add1[49], i_add1[50], i_add1[51], i_add1[52], i_add1[53], i_add1[54], i_add1[55], i_add1[56], i_add1[57], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], i_add2[19], i_add2[20], i_add2[21], i_add2[22], i_add2[23], i_add2[24], i_add2[25], i_add2[26], i_add2[27], i_add2[28], i_add2[29], i_add2[30], i_add2[31], i_add2[32], i_add2[33], i_add2[34], i_add2[35], i_add2[36], i_add2[37], i_add2[38], i_add2[39], i_add2[40], i_add2[41], i_add2[42], i_add2[43], i_add2[44], i_add2[45], i_add2[46], i_add2[47], i_add2[48], i_add2[49], i_add2[50], i_add2[51], i_add2[52], i_add2[53], i_add2[54], i_add2[55], i_add2[56], i_add2[57], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21], o_result[22], o_result[23], o_result[24], o_result[25], o_result[26], o_result[27], o_result[28], o_result[29], o_result[30], o_result[31], o_result[32], o_result[33], o_result[34], o_result[35], o_result[36], o_result[37], o_result[38], o_result[39], o_result[40], o_result[41], o_result[42], o_result[43], o_result[44], o_result[45], o_result[46], o_result[47], o_result[48], o_result[49], o_result[50], o_result[51], o_result[52], o_result[53], o_result[54], o_result[55], o_result[56], o_result[57], o_result[58]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add1[19];
input i_add1[20];
input i_add1[21];
input i_add1[22];
input i_add1[23];
input i_add1[24];
input i_add1[25];
input i_add1[26];
input i_add1[27];
input i_add1[28];
input i_add1[29];
input i_add1[30];
input i_add1[31];
input i_add1[32];
input i_add1[33];
input i_add1[34];
input i_add1[35];
input i_add1[36];
input i_add1[37];
input i_add1[38];
input i_add1[39];
input i_add1[40];
input i_add1[41];
input i_add1[42];
input i_add1[43];
input i_add1[44];
input i_add1[45];
input i_add1[46];
input i_add1[47];
input i_add1[48];
input i_add1[49];
input i_add1[50];
input i_add1[51];
input i_add1[52];
input i_add1[53];
input i_add1[54];
input i_add1[55];
input i_add1[56];
input i_add1[57];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
input i_add2[19];
input i_add2[20];
input i_add2[21];
input i_add2[22];
input i_add2[23];
input i_add2[24];
input i_add2[25];
input i_add2[26];
input i_add2[27];
input i_add2[28];
input i_add2[29];
input i_add2[30];
input i_add2[31];
input i_add2[32];
input i_add2[33];
input i_add2[34];
input i_add2[35];
input i_add2[36];
input i_add2[37];
input i_add2[38];
input i_add2[39];
input i_add2[40];
input i_add2[41];
input i_add2[42];
input i_add2[43];
input i_add2[44];
input i_add2[45];
input i_add2[46];
input i_add2[47];
input i_add2[48];
input i_add2[49];
input i_add2[50];
input i_add2[51];
input i_add2[52];
input i_add2[53];
input i_add2[54];
input i_add2[55];
input i_add2[56];
input i_add2[57];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];
output o_result[22];
output o_result[23];
output o_result[24];
output o_result[25];
output o_result[26];
output o_result[27];
output o_result[28];
output o_result[29];
output o_result[30];
output o_result[31];
output o_result[32];
output o_result[33];
output o_result[34];
output o_result[35];
output o_result[36];
output o_result[37];
output o_result[38];
output o_result[39];
output o_result[40];
output o_result[41];
output o_result[42];
output o_result[43];
output o_result[44];
output o_result[45];
output o_result[46];
output o_result[47];
output o_result[48];
output o_result[49];
output o_result[50];
output o_result[51];
output o_result[52];
output o_result[53];
output o_result[54];
output o_result[55];
output o_result[56];
output o_result[57];
output o_result[58];

NAND3X1 NAND3X1_1 ( .A(_299_), .B(_308_), .C(_307_), .Y(_309_) );
OAI21X1 OAI21X1_1 ( .A(_297_), .B(_298_), .C(_309_), .Y(w_C_52_) );
INVX1 INVX1_1 ( .A(i_add2[52]), .Y(_310_) );
INVX1 INVX1_2 ( .A(i_add1[52]), .Y(_311_) );
OAI21X1 OAI21X1_2 ( .A(i_add2[52]), .B(i_add1[52]), .C(w_C_52_), .Y(_312_) );
OAI21X1 OAI21X1_3 ( .A(_310_), .B(_311_), .C(_312_), .Y(w_C_53_) );
NOR2X1 NOR2X1_1 ( .A(_310_), .B(_311_), .Y(_313_) );
INVX1 INVX1_3 ( .A(_313_), .Y(_314_) );
AND2X2 AND2X2_1 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_315_) );
INVX1 INVX1_4 ( .A(_315_), .Y(_316_) );
NAND3X1 NAND3X1_2 ( .A(_314_), .B(_316_), .C(_312_), .Y(_317_) );
OAI21X1 OAI21X1_4 ( .A(i_add2[53]), .B(i_add1[53]), .C(_317_), .Y(_318_) );
INVX1 INVX1_5 ( .A(_318_), .Y(w_C_54_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_319_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_320_) );
OAI21X1 OAI21X1_5 ( .A(_320_), .B(_318_), .C(_319_), .Y(w_C_55_) );
NAND2X1 NAND2X1_2 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_321_) );
INVX1 INVX1_6 ( .A(_320_), .Y(_322_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_323_) );
INVX1 INVX1_7 ( .A(_323_), .Y(_324_) );
NOR2X1 NOR2X1_4 ( .A(_297_), .B(_298_), .Y(_325_) );
INVX1 INVX1_8 ( .A(_325_), .Y(_326_) );
NAND3X1 NAND3X1_3 ( .A(_326_), .B(_314_), .C(_309_), .Y(_327_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_328_) );
INVX1 INVX1_9 ( .A(_328_), .Y(_329_) );
NAND3X1 NAND3X1_4 ( .A(_324_), .B(_329_), .C(_327_), .Y(_330_) );
NAND3X1 NAND3X1_5 ( .A(_316_), .B(_319_), .C(_330_), .Y(_331_) );
OR2X2 OR2X2_1 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_332_) );
NAND3X1 NAND3X1_6 ( .A(_322_), .B(_332_), .C(_331_), .Y(_333_) );
NAND2X1 NAND2X1_3 ( .A(_321_), .B(_333_), .Y(w_C_56_) );
OR2X2 OR2X2_2 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_334_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_335_) );
NAND3X1 NAND3X1_7 ( .A(_321_), .B(_335_), .C(_333_), .Y(_336_) );
AND2X2 AND2X2_2 ( .A(_336_), .B(_334_), .Y(w_C_57_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_337_) );
OR2X2 OR2X2_3 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_338_) );
NAND3X1 NAND3X1_8 ( .A(_334_), .B(_338_), .C(_336_), .Y(_339_) );
NAND2X1 NAND2X1_6 ( .A(_337_), .B(_339_), .Y(w_C_58_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_10 ( .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_7 ( .A(_1_), .B(_2_), .Y(w_C_2_) );
INVX1 INVX1_11 ( .A(i_add2[2]), .Y(_3_) );
INVX1 INVX1_12 ( .A(i_add1[2]), .Y(_4_) );
NAND2X1 NAND2X1_8 ( .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
OAI21X1 OAI21X1_6 ( .A(_1_), .B(_2_), .C(_6_), .Y(_7_) );
AND2X2 AND2X2_3 ( .A(_7_), .B(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
OR2X2 OR2X2_4 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_9 ( .A(_5_), .B(_9_), .C(_7_), .Y(_10_) );
NAND2X1 NAND2X1_11 ( .A(_8_), .B(_10_), .Y(w_C_4_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
INVX1 INVX1_13 ( .A(_11_), .Y(_12_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
NAND3X1 NAND3X1_10 ( .A(_8_), .B(_13_), .C(_10_), .Y(_14_) );
AND2X2 AND2X2_4 ( .A(_14_), .B(_12_), .Y(w_C_5_) );
AND2X2 AND2X2_5 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_15_) );
INVX1 INVX1_14 ( .A(_15_), .Y(_16_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_17_) );
INVX1 INVX1_15 ( .A(_17_), .Y(_18_) );
NAND3X1 NAND3X1_11 ( .A(_12_), .B(_18_), .C(_14_), .Y(_19_) );
AND2X2 AND2X2_6 ( .A(_19_), .B(_16_), .Y(_20_) );
INVX1 INVX1_16 ( .A(_20_), .Y(w_C_6_) );
AND2X2 AND2X2_7 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_21_) );
INVX1 INVX1_17 ( .A(_21_), .Y(_22_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_23_) );
OAI21X1 OAI21X1_7 ( .A(_23_), .B(_20_), .C(_22_), .Y(w_C_7_) );
AND2X2 AND2X2_8 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_24_) );
INVX1 INVX1_18 ( .A(_24_), .Y(_25_) );
INVX1 INVX1_19 ( .A(_23_), .Y(_26_) );
NAND3X1 NAND3X1_12 ( .A(_16_), .B(_22_), .C(_19_), .Y(_27_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_28_) );
INVX1 INVX1_20 ( .A(_28_), .Y(_29_) );
NAND3X1 NAND3X1_13 ( .A(_26_), .B(_29_), .C(_27_), .Y(_30_) );
AND2X2 AND2X2_9 ( .A(_30_), .B(_25_), .Y(_31_) );
INVX1 INVX1_21 ( .A(_31_), .Y(w_C_8_) );
AND2X2 AND2X2_10 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_32_) );
INVX1 INVX1_22 ( .A(_32_), .Y(_33_) );
NAND3X1 NAND3X1_14 ( .A(_25_), .B(_33_), .C(_30_), .Y(_34_) );
OAI21X1 OAI21X1_8 ( .A(i_add2[8]), .B(i_add1[8]), .C(_34_), .Y(_35_) );
INVX1 INVX1_23 ( .A(_35_), .Y(w_C_9_) );
INVX1 INVX1_24 ( .A(i_add2[9]), .Y(_36_) );
INVX1 INVX1_25 ( .A(i_add1[9]), .Y(_37_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_38_) );
INVX1 INVX1_26 ( .A(_38_), .Y(_39_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_40_) );
INVX1 INVX1_27 ( .A(_40_), .Y(_41_) );
NAND3X1 NAND3X1_15 ( .A(_39_), .B(_41_), .C(_34_), .Y(_42_) );
OAI21X1 OAI21X1_9 ( .A(_36_), .B(_37_), .C(_42_), .Y(w_C_10_) );
NOR2X1 NOR2X1_14 ( .A(_36_), .B(_37_), .Y(_43_) );
INVX1 INVX1_28 ( .A(_43_), .Y(_44_) );
AND2X2 AND2X2_11 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_45_) );
INVX1 INVX1_29 ( .A(_45_), .Y(_46_) );
NAND3X1 NAND3X1_16 ( .A(_44_), .B(_46_), .C(_42_), .Y(_47_) );
OAI21X1 OAI21X1_10 ( .A(i_add2[10]), .B(i_add1[10]), .C(_47_), .Y(_48_) );
INVX1 INVX1_30 ( .A(_48_), .Y(w_C_11_) );
INVX1 INVX1_31 ( .A(i_add2[11]), .Y(_49_) );
INVX1 INVX1_32 ( .A(i_add1[11]), .Y(_50_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_51_) );
INVX1 INVX1_33 ( .A(_51_), .Y(_52_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_53_) );
INVX1 INVX1_34 ( .A(_53_), .Y(_54_) );
NAND3X1 NAND3X1_17 ( .A(_52_), .B(_54_), .C(_47_), .Y(_55_) );
OAI21X1 OAI21X1_11 ( .A(_49_), .B(_50_), .C(_55_), .Y(w_C_12_) );
NOR2X1 NOR2X1_17 ( .A(_49_), .B(_50_), .Y(_56_) );
INVX1 INVX1_35 ( .A(_56_), .Y(_57_) );
AND2X2 AND2X2_12 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_58_) );
INVX1 INVX1_36 ( .A(_58_), .Y(_59_) );
NAND3X1 NAND3X1_18 ( .A(_57_), .B(_59_), .C(_55_), .Y(_60_) );
OAI21X1 OAI21X1_12 ( .A(i_add2[12]), .B(i_add1[12]), .C(_60_), .Y(_61_) );
INVX1 INVX1_37 ( .A(_61_), .Y(w_C_13_) );
INVX1 INVX1_38 ( .A(i_add2[13]), .Y(_62_) );
INVX1 INVX1_39 ( .A(i_add1[13]), .Y(_63_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_64_) );
INVX1 INVX1_40 ( .A(_64_), .Y(_65_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_66_) );
INVX1 INVX1_41 ( .A(_66_), .Y(_67_) );
NAND3X1 NAND3X1_19 ( .A(_65_), .B(_67_), .C(_60_), .Y(_68_) );
OAI21X1 OAI21X1_13 ( .A(_62_), .B(_63_), .C(_68_), .Y(w_C_14_) );
NOR2X1 NOR2X1_20 ( .A(_62_), .B(_63_), .Y(_69_) );
INVX1 INVX1_42 ( .A(_69_), .Y(_70_) );
AND2X2 AND2X2_13 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_71_) );
INVX1 INVX1_43 ( .A(_71_), .Y(_72_) );
NAND3X1 NAND3X1_20 ( .A(_70_), .B(_72_), .C(_68_), .Y(_73_) );
OAI21X1 OAI21X1_14 ( .A(i_add2[14]), .B(i_add1[14]), .C(_73_), .Y(_74_) );
INVX1 INVX1_44 ( .A(_74_), .Y(w_C_15_) );
INVX1 INVX1_45 ( .A(i_add2[15]), .Y(_75_) );
INVX1 INVX1_46 ( .A(i_add1[15]), .Y(_76_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_77_) );
INVX1 INVX1_47 ( .A(_77_), .Y(_78_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_79_) );
INVX1 INVX1_48 ( .A(_79_), .Y(_80_) );
NAND3X1 NAND3X1_21 ( .A(_78_), .B(_80_), .C(_73_), .Y(_81_) );
OAI21X1 OAI21X1_15 ( .A(_75_), .B(_76_), .C(_81_), .Y(w_C_16_) );
NOR2X1 NOR2X1_23 ( .A(_75_), .B(_76_), .Y(_82_) );
INVX1 INVX1_49 ( .A(_82_), .Y(_83_) );
AND2X2 AND2X2_14 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_84_) );
INVX1 INVX1_50 ( .A(_84_), .Y(_85_) );
NAND3X1 NAND3X1_22 ( .A(_83_), .B(_85_), .C(_81_), .Y(_86_) );
OAI21X1 OAI21X1_16 ( .A(i_add2[16]), .B(i_add1[16]), .C(_86_), .Y(_87_) );
INVX1 INVX1_51 ( .A(_87_), .Y(w_C_17_) );
INVX1 INVX1_52 ( .A(i_add2[17]), .Y(_88_) );
INVX1 INVX1_53 ( .A(i_add1[17]), .Y(_89_) );
BUFX2 BUFX2_1 ( .A(_340__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_340__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_340__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_340__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_340__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_340__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_340__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_340__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_340__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_340__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_340__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_340__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_340__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_340__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_340__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_340__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_340__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_340__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_340__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_340__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_340__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_340__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_340__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_340__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_340__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_340__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_340__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_340__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_340__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_340__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_340__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_340__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_340__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_340__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_340__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_340__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_340__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(_340__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .A(_340__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .A(_340__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .A(_340__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .A(_340__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .A(_340__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .A(_340__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .A(_340__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .A(_340__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .A(_340__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .A(_340__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .A(_340__48_), .Y(o_result[48]) );
BUFX2 BUFX2_50 ( .A(_340__49_), .Y(o_result[49]) );
BUFX2 BUFX2_51 ( .A(_340__50_), .Y(o_result[50]) );
BUFX2 BUFX2_52 ( .A(_340__51_), .Y(o_result[51]) );
BUFX2 BUFX2_53 ( .A(_340__52_), .Y(o_result[52]) );
BUFX2 BUFX2_54 ( .A(_340__53_), .Y(o_result[53]) );
BUFX2 BUFX2_55 ( .A(_340__54_), .Y(o_result[54]) );
BUFX2 BUFX2_56 ( .A(_340__55_), .Y(o_result[55]) );
BUFX2 BUFX2_57 ( .A(_340__56_), .Y(o_result[56]) );
BUFX2 BUFX2_58 ( .A(_340__57_), .Y(o_result[57]) );
BUFX2 BUFX2_59 ( .A(w_C_58_), .Y(o_result[58]) );
INVX1 INVX1_54 ( .A(w_C_4_), .Y(_344_) );
OR2X2 OR2X2_5 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_345_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_346_) );
NAND3X1 NAND3X1_23 ( .A(_344_), .B(_346_), .C(_345_), .Y(_347_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_341_) );
AND2X2 AND2X2_15 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_342_) );
OAI21X1 OAI21X1_17 ( .A(_341_), .B(_342_), .C(w_C_4_), .Y(_343_) );
NAND2X1 NAND2X1_14 ( .A(_343_), .B(_347_), .Y(_340__4_) );
INVX1 INVX1_55 ( .A(w_C_5_), .Y(_351_) );
OR2X2 OR2X2_6 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_352_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_353_) );
NAND3X1 NAND3X1_24 ( .A(_351_), .B(_353_), .C(_352_), .Y(_354_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_348_) );
AND2X2 AND2X2_16 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_349_) );
OAI21X1 OAI21X1_18 ( .A(_348_), .B(_349_), .C(w_C_5_), .Y(_350_) );
NAND2X1 NAND2X1_16 ( .A(_350_), .B(_354_), .Y(_340__5_) );
INVX1 INVX1_56 ( .A(w_C_6_), .Y(_358_) );
OR2X2 OR2X2_7 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_359_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_360_) );
NAND3X1 NAND3X1_25 ( .A(_358_), .B(_360_), .C(_359_), .Y(_361_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_355_) );
AND2X2 AND2X2_17 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_356_) );
OAI21X1 OAI21X1_19 ( .A(_355_), .B(_356_), .C(w_C_6_), .Y(_357_) );
NAND2X1 NAND2X1_18 ( .A(_357_), .B(_361_), .Y(_340__6_) );
INVX1 INVX1_57 ( .A(w_C_7_), .Y(_365_) );
OR2X2 OR2X2_8 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_366_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_367_) );
NAND3X1 NAND3X1_26 ( .A(_365_), .B(_367_), .C(_366_), .Y(_368_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_362_) );
AND2X2 AND2X2_18 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_363_) );
OAI21X1 OAI21X1_20 ( .A(_362_), .B(_363_), .C(w_C_7_), .Y(_364_) );
NAND2X1 NAND2X1_20 ( .A(_364_), .B(_368_), .Y(_340__7_) );
INVX1 INVX1_58 ( .A(w_C_8_), .Y(_372_) );
OR2X2 OR2X2_9 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_373_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_374_) );
NAND3X1 NAND3X1_27 ( .A(_372_), .B(_374_), .C(_373_), .Y(_375_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_369_) );
AND2X2 AND2X2_19 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_370_) );
OAI21X1 OAI21X1_21 ( .A(_369_), .B(_370_), .C(w_C_8_), .Y(_371_) );
NAND2X1 NAND2X1_22 ( .A(_371_), .B(_375_), .Y(_340__8_) );
INVX1 INVX1_59 ( .A(w_C_9_), .Y(_379_) );
OR2X2 OR2X2_10 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_380_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_381_) );
NAND3X1 NAND3X1_28 ( .A(_379_), .B(_381_), .C(_380_), .Y(_382_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_376_) );
AND2X2 AND2X2_20 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_377_) );
OAI21X1 OAI21X1_22 ( .A(_376_), .B(_377_), .C(w_C_9_), .Y(_378_) );
NAND2X1 NAND2X1_24 ( .A(_378_), .B(_382_), .Y(_340__9_) );
INVX1 INVX1_60 ( .A(w_C_10_), .Y(_386_) );
OR2X2 OR2X2_11 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_387_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_388_) );
NAND3X1 NAND3X1_29 ( .A(_386_), .B(_388_), .C(_387_), .Y(_389_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_383_) );
AND2X2 AND2X2_21 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_384_) );
OAI21X1 OAI21X1_23 ( .A(_383_), .B(_384_), .C(w_C_10_), .Y(_385_) );
NAND2X1 NAND2X1_26 ( .A(_385_), .B(_389_), .Y(_340__10_) );
INVX1 INVX1_61 ( .A(w_C_11_), .Y(_393_) );
OR2X2 OR2X2_12 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_394_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_395_) );
NAND3X1 NAND3X1_30 ( .A(_393_), .B(_395_), .C(_394_), .Y(_396_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_390_) );
AND2X2 AND2X2_22 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_391_) );
OAI21X1 OAI21X1_24 ( .A(_390_), .B(_391_), .C(w_C_11_), .Y(_392_) );
NAND2X1 NAND2X1_28 ( .A(_392_), .B(_396_), .Y(_340__11_) );
INVX1 INVX1_62 ( .A(w_C_12_), .Y(_400_) );
OR2X2 OR2X2_13 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_401_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_402_) );
NAND3X1 NAND3X1_31 ( .A(_400_), .B(_402_), .C(_401_), .Y(_403_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_397_) );
AND2X2 AND2X2_23 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_398_) );
OAI21X1 OAI21X1_25 ( .A(_397_), .B(_398_), .C(w_C_12_), .Y(_399_) );
NAND2X1 NAND2X1_30 ( .A(_399_), .B(_403_), .Y(_340__12_) );
INVX1 INVX1_63 ( .A(w_C_13_), .Y(_407_) );
OR2X2 OR2X2_14 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_408_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_409_) );
NAND3X1 NAND3X1_32 ( .A(_407_), .B(_409_), .C(_408_), .Y(_410_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_404_) );
AND2X2 AND2X2_24 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_405_) );
OAI21X1 OAI21X1_26 ( .A(_404_), .B(_405_), .C(w_C_13_), .Y(_406_) );
NAND2X1 NAND2X1_32 ( .A(_406_), .B(_410_), .Y(_340__13_) );
INVX1 INVX1_64 ( .A(w_C_14_), .Y(_414_) );
OR2X2 OR2X2_15 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_415_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_416_) );
NAND3X1 NAND3X1_33 ( .A(_414_), .B(_416_), .C(_415_), .Y(_417_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_411_) );
AND2X2 AND2X2_25 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_412_) );
OAI21X1 OAI21X1_27 ( .A(_411_), .B(_412_), .C(w_C_14_), .Y(_413_) );
NAND2X1 NAND2X1_34 ( .A(_413_), .B(_417_), .Y(_340__14_) );
INVX1 INVX1_65 ( .A(w_C_15_), .Y(_421_) );
OR2X2 OR2X2_16 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_422_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_423_) );
NAND3X1 NAND3X1_34 ( .A(_421_), .B(_423_), .C(_422_), .Y(_424_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_418_) );
AND2X2 AND2X2_26 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_419_) );
OAI21X1 OAI21X1_28 ( .A(_418_), .B(_419_), .C(w_C_15_), .Y(_420_) );
NAND2X1 NAND2X1_36 ( .A(_420_), .B(_424_), .Y(_340__15_) );
INVX1 INVX1_66 ( .A(w_C_16_), .Y(_428_) );
OR2X2 OR2X2_17 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_429_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_430_) );
NAND3X1 NAND3X1_35 ( .A(_428_), .B(_430_), .C(_429_), .Y(_431_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_425_) );
AND2X2 AND2X2_27 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_426_) );
OAI21X1 OAI21X1_29 ( .A(_425_), .B(_426_), .C(w_C_16_), .Y(_427_) );
NAND2X1 NAND2X1_38 ( .A(_427_), .B(_431_), .Y(_340__16_) );
INVX1 INVX1_67 ( .A(w_C_17_), .Y(_435_) );
OR2X2 OR2X2_18 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_436_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_437_) );
NAND3X1 NAND3X1_36 ( .A(_435_), .B(_437_), .C(_436_), .Y(_438_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_432_) );
AND2X2 AND2X2_28 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_433_) );
OAI21X1 OAI21X1_30 ( .A(_432_), .B(_433_), .C(w_C_17_), .Y(_434_) );
NAND2X1 NAND2X1_40 ( .A(_434_), .B(_438_), .Y(_340__17_) );
INVX1 INVX1_68 ( .A(w_C_18_), .Y(_442_) );
OR2X2 OR2X2_19 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_443_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_444_) );
NAND3X1 NAND3X1_37 ( .A(_442_), .B(_444_), .C(_443_), .Y(_445_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_439_) );
AND2X2 AND2X2_29 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_440_) );
OAI21X1 OAI21X1_31 ( .A(_439_), .B(_440_), .C(w_C_18_), .Y(_441_) );
NAND2X1 NAND2X1_42 ( .A(_441_), .B(_445_), .Y(_340__18_) );
INVX1 INVX1_69 ( .A(w_C_19_), .Y(_449_) );
OR2X2 OR2X2_20 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_450_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_451_) );
NAND3X1 NAND3X1_38 ( .A(_449_), .B(_451_), .C(_450_), .Y(_452_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_446_) );
AND2X2 AND2X2_30 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_447_) );
OAI21X1 OAI21X1_32 ( .A(_446_), .B(_447_), .C(w_C_19_), .Y(_448_) );
NAND2X1 NAND2X1_44 ( .A(_448_), .B(_452_), .Y(_340__19_) );
INVX1 INVX1_70 ( .A(w_C_20_), .Y(_456_) );
OR2X2 OR2X2_21 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_457_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_458_) );
NAND3X1 NAND3X1_39 ( .A(_456_), .B(_458_), .C(_457_), .Y(_459_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_453_) );
AND2X2 AND2X2_31 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_454_) );
OAI21X1 OAI21X1_33 ( .A(_453_), .B(_454_), .C(w_C_20_), .Y(_455_) );
NAND2X1 NAND2X1_46 ( .A(_455_), .B(_459_), .Y(_340__20_) );
INVX1 INVX1_71 ( .A(w_C_21_), .Y(_463_) );
OR2X2 OR2X2_22 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_464_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_465_) );
NAND3X1 NAND3X1_40 ( .A(_463_), .B(_465_), .C(_464_), .Y(_466_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_460_) );
AND2X2 AND2X2_32 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_461_) );
OAI21X1 OAI21X1_34 ( .A(_460_), .B(_461_), .C(w_C_21_), .Y(_462_) );
NAND2X1 NAND2X1_48 ( .A(_462_), .B(_466_), .Y(_340__21_) );
INVX1 INVX1_72 ( .A(w_C_22_), .Y(_470_) );
OR2X2 OR2X2_23 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_471_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_472_) );
NAND3X1 NAND3X1_41 ( .A(_470_), .B(_472_), .C(_471_), .Y(_473_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_467_) );
AND2X2 AND2X2_33 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_468_) );
OAI21X1 OAI21X1_35 ( .A(_467_), .B(_468_), .C(w_C_22_), .Y(_469_) );
NAND2X1 NAND2X1_50 ( .A(_469_), .B(_473_), .Y(_340__22_) );
INVX1 INVX1_73 ( .A(w_C_23_), .Y(_477_) );
OR2X2 OR2X2_24 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_478_) );
NAND2X1 NAND2X1_51 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_479_) );
NAND3X1 NAND3X1_42 ( .A(_477_), .B(_479_), .C(_478_), .Y(_480_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_474_) );
AND2X2 AND2X2_34 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_475_) );
OAI21X1 OAI21X1_36 ( .A(_474_), .B(_475_), .C(w_C_23_), .Y(_476_) );
NAND2X1 NAND2X1_52 ( .A(_476_), .B(_480_), .Y(_340__23_) );
INVX1 INVX1_74 ( .A(w_C_24_), .Y(_484_) );
OR2X2 OR2X2_25 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_485_) );
NAND2X1 NAND2X1_53 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_486_) );
NAND3X1 NAND3X1_43 ( .A(_484_), .B(_486_), .C(_485_), .Y(_487_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_481_) );
AND2X2 AND2X2_35 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_482_) );
OAI21X1 OAI21X1_37 ( .A(_481_), .B(_482_), .C(w_C_24_), .Y(_483_) );
NAND2X1 NAND2X1_54 ( .A(_483_), .B(_487_), .Y(_340__24_) );
INVX1 INVX1_75 ( .A(w_C_25_), .Y(_491_) );
OR2X2 OR2X2_26 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_492_) );
NAND2X1 NAND2X1_55 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_493_) );
NAND3X1 NAND3X1_44 ( .A(_491_), .B(_493_), .C(_492_), .Y(_494_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_488_) );
AND2X2 AND2X2_36 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_489_) );
OAI21X1 OAI21X1_38 ( .A(_488_), .B(_489_), .C(w_C_25_), .Y(_490_) );
NAND2X1 NAND2X1_56 ( .A(_490_), .B(_494_), .Y(_340__25_) );
INVX1 INVX1_76 ( .A(w_C_26_), .Y(_498_) );
OR2X2 OR2X2_27 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_499_) );
NAND2X1 NAND2X1_57 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_500_) );
NAND3X1 NAND3X1_45 ( .A(_498_), .B(_500_), .C(_499_), .Y(_501_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_495_) );
AND2X2 AND2X2_37 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_496_) );
OAI21X1 OAI21X1_39 ( .A(_495_), .B(_496_), .C(w_C_26_), .Y(_497_) );
NAND2X1 NAND2X1_58 ( .A(_497_), .B(_501_), .Y(_340__26_) );
INVX1 INVX1_77 ( .A(w_C_27_), .Y(_505_) );
OR2X2 OR2X2_28 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_506_) );
NAND2X1 NAND2X1_59 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_507_) );
NAND3X1 NAND3X1_46 ( .A(_505_), .B(_507_), .C(_506_), .Y(_508_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_502_) );
AND2X2 AND2X2_38 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_503_) );
OAI21X1 OAI21X1_40 ( .A(_502_), .B(_503_), .C(w_C_27_), .Y(_504_) );
NAND2X1 NAND2X1_60 ( .A(_504_), .B(_508_), .Y(_340__27_) );
INVX1 INVX1_78 ( .A(w_C_28_), .Y(_512_) );
OR2X2 OR2X2_29 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_513_) );
NAND2X1 NAND2X1_61 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_514_) );
NAND3X1 NAND3X1_47 ( .A(_512_), .B(_514_), .C(_513_), .Y(_515_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_509_) );
AND2X2 AND2X2_39 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_510_) );
OAI21X1 OAI21X1_41 ( .A(_509_), .B(_510_), .C(w_C_28_), .Y(_511_) );
NAND2X1 NAND2X1_62 ( .A(_511_), .B(_515_), .Y(_340__28_) );
INVX1 INVX1_79 ( .A(w_C_29_), .Y(_519_) );
OR2X2 OR2X2_30 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_520_) );
NAND2X1 NAND2X1_63 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_521_) );
NAND3X1 NAND3X1_48 ( .A(_519_), .B(_521_), .C(_520_), .Y(_522_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_516_) );
AND2X2 AND2X2_40 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_517_) );
OAI21X1 OAI21X1_42 ( .A(_516_), .B(_517_), .C(w_C_29_), .Y(_518_) );
NAND2X1 NAND2X1_64 ( .A(_518_), .B(_522_), .Y(_340__29_) );
INVX1 INVX1_80 ( .A(w_C_30_), .Y(_526_) );
OR2X2 OR2X2_31 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_527_) );
NAND2X1 NAND2X1_65 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_528_) );
NAND3X1 NAND3X1_49 ( .A(_526_), .B(_528_), .C(_527_), .Y(_529_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_523_) );
AND2X2 AND2X2_41 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_524_) );
OAI21X1 OAI21X1_43 ( .A(_523_), .B(_524_), .C(w_C_30_), .Y(_525_) );
NAND2X1 NAND2X1_66 ( .A(_525_), .B(_529_), .Y(_340__30_) );
INVX1 INVX1_81 ( .A(w_C_31_), .Y(_533_) );
OR2X2 OR2X2_32 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_534_) );
NAND2X1 NAND2X1_67 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_535_) );
NAND3X1 NAND3X1_50 ( .A(_533_), .B(_535_), .C(_534_), .Y(_536_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_530_) );
AND2X2 AND2X2_42 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_531_) );
OAI21X1 OAI21X1_44 ( .A(_530_), .B(_531_), .C(w_C_31_), .Y(_532_) );
NAND2X1 NAND2X1_68 ( .A(_532_), .B(_536_), .Y(_340__31_) );
INVX1 INVX1_82 ( .A(w_C_32_), .Y(_540_) );
OR2X2 OR2X2_33 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_541_) );
NAND2X1 NAND2X1_69 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_542_) );
NAND3X1 NAND3X1_51 ( .A(_540_), .B(_542_), .C(_541_), .Y(_543_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_537_) );
AND2X2 AND2X2_43 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_538_) );
OAI21X1 OAI21X1_45 ( .A(_537_), .B(_538_), .C(w_C_32_), .Y(_539_) );
NAND2X1 NAND2X1_70 ( .A(_539_), .B(_543_), .Y(_340__32_) );
INVX1 INVX1_83 ( .A(w_C_33_), .Y(_547_) );
OR2X2 OR2X2_34 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_548_) );
NAND2X1 NAND2X1_71 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_549_) );
NAND3X1 NAND3X1_52 ( .A(_547_), .B(_549_), .C(_548_), .Y(_550_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_544_) );
AND2X2 AND2X2_44 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_545_) );
OAI21X1 OAI21X1_46 ( .A(_544_), .B(_545_), .C(w_C_33_), .Y(_546_) );
NAND2X1 NAND2X1_72 ( .A(_546_), .B(_550_), .Y(_340__33_) );
INVX1 INVX1_84 ( .A(w_C_34_), .Y(_554_) );
OR2X2 OR2X2_35 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_555_) );
NAND2X1 NAND2X1_73 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_556_) );
NAND3X1 NAND3X1_53 ( .A(_554_), .B(_556_), .C(_555_), .Y(_557_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_551_) );
AND2X2 AND2X2_45 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_552_) );
OAI21X1 OAI21X1_47 ( .A(_551_), .B(_552_), .C(w_C_34_), .Y(_553_) );
NAND2X1 NAND2X1_74 ( .A(_553_), .B(_557_), .Y(_340__34_) );
INVX1 INVX1_85 ( .A(w_C_35_), .Y(_561_) );
OR2X2 OR2X2_36 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_562_) );
NAND2X1 NAND2X1_75 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_563_) );
NAND3X1 NAND3X1_54 ( .A(_561_), .B(_563_), .C(_562_), .Y(_564_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_558_) );
AND2X2 AND2X2_46 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_559_) );
OAI21X1 OAI21X1_48 ( .A(_558_), .B(_559_), .C(w_C_35_), .Y(_560_) );
NAND2X1 NAND2X1_76 ( .A(_560_), .B(_564_), .Y(_340__35_) );
INVX1 INVX1_86 ( .A(w_C_36_), .Y(_568_) );
OR2X2 OR2X2_37 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_569_) );
NAND2X1 NAND2X1_77 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_570_) );
NAND3X1 NAND3X1_55 ( .A(_568_), .B(_570_), .C(_569_), .Y(_571_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_565_) );
AND2X2 AND2X2_47 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_566_) );
OAI21X1 OAI21X1_49 ( .A(_565_), .B(_566_), .C(w_C_36_), .Y(_567_) );
NAND2X1 NAND2X1_78 ( .A(_567_), .B(_571_), .Y(_340__36_) );
INVX1 INVX1_87 ( .A(w_C_37_), .Y(_575_) );
OR2X2 OR2X2_38 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_576_) );
NAND2X1 NAND2X1_79 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_577_) );
NAND3X1 NAND3X1_56 ( .A(_575_), .B(_577_), .C(_576_), .Y(_578_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_572_) );
AND2X2 AND2X2_48 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_573_) );
OAI21X1 OAI21X1_50 ( .A(_572_), .B(_573_), .C(w_C_37_), .Y(_574_) );
NAND2X1 NAND2X1_80 ( .A(_574_), .B(_578_), .Y(_340__37_) );
INVX1 INVX1_88 ( .A(w_C_38_), .Y(_582_) );
OR2X2 OR2X2_39 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_583_) );
NAND2X1 NAND2X1_81 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_584_) );
NAND3X1 NAND3X1_57 ( .A(_582_), .B(_584_), .C(_583_), .Y(_585_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_579_) );
AND2X2 AND2X2_49 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_580_) );
OAI21X1 OAI21X1_51 ( .A(_579_), .B(_580_), .C(w_C_38_), .Y(_581_) );
NAND2X1 NAND2X1_82 ( .A(_581_), .B(_585_), .Y(_340__38_) );
INVX1 INVX1_89 ( .A(w_C_39_), .Y(_589_) );
OR2X2 OR2X2_40 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_590_) );
NAND2X1 NAND2X1_83 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_591_) );
NAND3X1 NAND3X1_58 ( .A(_589_), .B(_591_), .C(_590_), .Y(_592_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_586_) );
AND2X2 AND2X2_50 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_587_) );
OAI21X1 OAI21X1_52 ( .A(_586_), .B(_587_), .C(w_C_39_), .Y(_588_) );
NAND2X1 NAND2X1_84 ( .A(_588_), .B(_592_), .Y(_340__39_) );
INVX1 INVX1_90 ( .A(w_C_40_), .Y(_596_) );
OR2X2 OR2X2_41 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_597_) );
NAND2X1 NAND2X1_85 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_598_) );
NAND3X1 NAND3X1_59 ( .A(_596_), .B(_598_), .C(_597_), .Y(_599_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_593_) );
AND2X2 AND2X2_51 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_594_) );
OAI21X1 OAI21X1_53 ( .A(_593_), .B(_594_), .C(w_C_40_), .Y(_595_) );
NAND2X1 NAND2X1_86 ( .A(_595_), .B(_599_), .Y(_340__40_) );
INVX1 INVX1_91 ( .A(w_C_41_), .Y(_603_) );
OR2X2 OR2X2_42 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_604_) );
NAND2X1 NAND2X1_87 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_605_) );
NAND3X1 NAND3X1_60 ( .A(_603_), .B(_605_), .C(_604_), .Y(_606_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_600_) );
AND2X2 AND2X2_52 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_601_) );
OAI21X1 OAI21X1_54 ( .A(_600_), .B(_601_), .C(w_C_41_), .Y(_602_) );
NAND2X1 NAND2X1_88 ( .A(_602_), .B(_606_), .Y(_340__41_) );
INVX1 INVX1_92 ( .A(w_C_42_), .Y(_610_) );
OR2X2 OR2X2_43 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_611_) );
NAND2X1 NAND2X1_89 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_612_) );
NAND3X1 NAND3X1_61 ( .A(_610_), .B(_612_), .C(_611_), .Y(_613_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_607_) );
AND2X2 AND2X2_53 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_608_) );
OAI21X1 OAI21X1_55 ( .A(_607_), .B(_608_), .C(w_C_42_), .Y(_609_) );
NAND2X1 NAND2X1_90 ( .A(_609_), .B(_613_), .Y(_340__42_) );
INVX1 INVX1_93 ( .A(w_C_43_), .Y(_617_) );
OR2X2 OR2X2_44 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_618_) );
NAND2X1 NAND2X1_91 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_619_) );
NAND3X1 NAND3X1_62 ( .A(_617_), .B(_619_), .C(_618_), .Y(_620_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_614_) );
AND2X2 AND2X2_54 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_615_) );
OAI21X1 OAI21X1_56 ( .A(_614_), .B(_615_), .C(w_C_43_), .Y(_616_) );
NAND2X1 NAND2X1_92 ( .A(_616_), .B(_620_), .Y(_340__43_) );
INVX1 INVX1_94 ( .A(w_C_44_), .Y(_624_) );
OR2X2 OR2X2_45 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_625_) );
NAND2X1 NAND2X1_93 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_626_) );
NAND3X1 NAND3X1_63 ( .A(_624_), .B(_626_), .C(_625_), .Y(_627_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_621_) );
AND2X2 AND2X2_55 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_622_) );
OAI21X1 OAI21X1_57 ( .A(_621_), .B(_622_), .C(w_C_44_), .Y(_623_) );
NAND2X1 NAND2X1_94 ( .A(_623_), .B(_627_), .Y(_340__44_) );
INVX1 INVX1_95 ( .A(w_C_45_), .Y(_631_) );
OR2X2 OR2X2_46 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_632_) );
NAND2X1 NAND2X1_95 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_633_) );
NAND3X1 NAND3X1_64 ( .A(_631_), .B(_633_), .C(_632_), .Y(_634_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_628_) );
AND2X2 AND2X2_56 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_629_) );
OAI21X1 OAI21X1_58 ( .A(_628_), .B(_629_), .C(w_C_45_), .Y(_630_) );
NAND2X1 NAND2X1_96 ( .A(_630_), .B(_634_), .Y(_340__45_) );
INVX1 INVX1_96 ( .A(w_C_46_), .Y(_638_) );
OR2X2 OR2X2_47 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_639_) );
NAND2X1 NAND2X1_97 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_640_) );
NAND3X1 NAND3X1_65 ( .A(_638_), .B(_640_), .C(_639_), .Y(_641_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_635_) );
AND2X2 AND2X2_57 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_636_) );
OAI21X1 OAI21X1_59 ( .A(_635_), .B(_636_), .C(w_C_46_), .Y(_637_) );
NAND2X1 NAND2X1_98 ( .A(_637_), .B(_641_), .Y(_340__46_) );
INVX1 INVX1_97 ( .A(w_C_47_), .Y(_645_) );
OR2X2 OR2X2_48 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_646_) );
NAND2X1 NAND2X1_99 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_647_) );
NAND3X1 NAND3X1_66 ( .A(_645_), .B(_647_), .C(_646_), .Y(_648_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_642_) );
AND2X2 AND2X2_58 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_643_) );
OAI21X1 OAI21X1_60 ( .A(_642_), .B(_643_), .C(w_C_47_), .Y(_644_) );
NAND2X1 NAND2X1_100 ( .A(_644_), .B(_648_), .Y(_340__47_) );
INVX1 INVX1_98 ( .A(w_C_48_), .Y(_652_) );
OR2X2 OR2X2_49 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_653_) );
NAND2X1 NAND2X1_101 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_654_) );
NAND3X1 NAND3X1_67 ( .A(_652_), .B(_654_), .C(_653_), .Y(_655_) );
NOR2X1 NOR2X1_68 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_649_) );
AND2X2 AND2X2_59 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_650_) );
OAI21X1 OAI21X1_61 ( .A(_649_), .B(_650_), .C(w_C_48_), .Y(_651_) );
NAND2X1 NAND2X1_102 ( .A(_651_), .B(_655_), .Y(_340__48_) );
INVX1 INVX1_99 ( .A(w_C_49_), .Y(_659_) );
OR2X2 OR2X2_50 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_660_) );
NAND2X1 NAND2X1_103 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_661_) );
NAND3X1 NAND3X1_68 ( .A(_659_), .B(_661_), .C(_660_), .Y(_662_) );
NOR2X1 NOR2X1_69 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_656_) );
AND2X2 AND2X2_60 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_657_) );
OAI21X1 OAI21X1_62 ( .A(_656_), .B(_657_), .C(w_C_49_), .Y(_658_) );
NAND2X1 NAND2X1_104 ( .A(_658_), .B(_662_), .Y(_340__49_) );
INVX1 INVX1_100 ( .A(w_C_50_), .Y(_666_) );
OR2X2 OR2X2_51 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_667_) );
NAND2X1 NAND2X1_105 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_668_) );
NAND3X1 NAND3X1_69 ( .A(_666_), .B(_668_), .C(_667_), .Y(_669_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_663_) );
AND2X2 AND2X2_61 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_664_) );
OAI21X1 OAI21X1_63 ( .A(_663_), .B(_664_), .C(w_C_50_), .Y(_665_) );
NAND2X1 NAND2X1_106 ( .A(_665_), .B(_669_), .Y(_340__50_) );
INVX1 INVX1_101 ( .A(w_C_51_), .Y(_673_) );
OR2X2 OR2X2_52 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_674_) );
NAND2X1 NAND2X1_107 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_675_) );
NAND3X1 NAND3X1_70 ( .A(_673_), .B(_675_), .C(_674_), .Y(_676_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_670_) );
AND2X2 AND2X2_62 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_671_) );
OAI21X1 OAI21X1_64 ( .A(_670_), .B(_671_), .C(w_C_51_), .Y(_672_) );
NAND2X1 NAND2X1_108 ( .A(_672_), .B(_676_), .Y(_340__51_) );
INVX1 INVX1_102 ( .A(w_C_52_), .Y(_680_) );
OR2X2 OR2X2_53 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_681_) );
NAND2X1 NAND2X1_109 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_682_) );
NAND3X1 NAND3X1_71 ( .A(_680_), .B(_682_), .C(_681_), .Y(_683_) );
NOR2X1 NOR2X1_72 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_677_) );
AND2X2 AND2X2_63 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_678_) );
OAI21X1 OAI21X1_65 ( .A(_677_), .B(_678_), .C(w_C_52_), .Y(_679_) );
NAND2X1 NAND2X1_110 ( .A(_679_), .B(_683_), .Y(_340__52_) );
INVX1 INVX1_103 ( .A(w_C_53_), .Y(_687_) );
OR2X2 OR2X2_54 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_688_) );
NAND2X1 NAND2X1_111 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_689_) );
NAND3X1 NAND3X1_72 ( .A(_687_), .B(_689_), .C(_688_), .Y(_690_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_684_) );
AND2X2 AND2X2_64 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_685_) );
OAI21X1 OAI21X1_66 ( .A(_684_), .B(_685_), .C(w_C_53_), .Y(_686_) );
NAND2X1 NAND2X1_112 ( .A(_686_), .B(_690_), .Y(_340__53_) );
INVX1 INVX1_104 ( .A(w_C_54_), .Y(_694_) );
OR2X2 OR2X2_55 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_695_) );
NAND2X1 NAND2X1_113 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_696_) );
NAND3X1 NAND3X1_73 ( .A(_694_), .B(_696_), .C(_695_), .Y(_697_) );
NOR2X1 NOR2X1_74 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_691_) );
AND2X2 AND2X2_65 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_692_) );
OAI21X1 OAI21X1_67 ( .A(_691_), .B(_692_), .C(w_C_54_), .Y(_693_) );
NAND2X1 NAND2X1_114 ( .A(_693_), .B(_697_), .Y(_340__54_) );
INVX1 INVX1_105 ( .A(w_C_55_), .Y(_701_) );
OR2X2 OR2X2_56 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_702_) );
NAND2X1 NAND2X1_115 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_703_) );
NAND3X1 NAND3X1_74 ( .A(_701_), .B(_703_), .C(_702_), .Y(_704_) );
NOR2X1 NOR2X1_75 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_698_) );
AND2X2 AND2X2_66 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_699_) );
OAI21X1 OAI21X1_68 ( .A(_698_), .B(_699_), .C(w_C_55_), .Y(_700_) );
NAND2X1 NAND2X1_116 ( .A(_700_), .B(_704_), .Y(_340__55_) );
INVX1 INVX1_106 ( .A(w_C_56_), .Y(_708_) );
OR2X2 OR2X2_57 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_709_) );
NAND2X1 NAND2X1_117 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_710_) );
NAND3X1 NAND3X1_75 ( .A(_708_), .B(_710_), .C(_709_), .Y(_711_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_705_) );
AND2X2 AND2X2_67 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_706_) );
OAI21X1 OAI21X1_69 ( .A(_705_), .B(_706_), .C(w_C_56_), .Y(_707_) );
NAND2X1 NAND2X1_118 ( .A(_707_), .B(_711_), .Y(_340__56_) );
INVX1 INVX1_107 ( .A(w_C_57_), .Y(_715_) );
OR2X2 OR2X2_58 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_716_) );
NAND2X1 NAND2X1_119 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_717_) );
NAND3X1 NAND3X1_76 ( .A(_715_), .B(_717_), .C(_716_), .Y(_718_) );
NOR2X1 NOR2X1_77 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_712_) );
AND2X2 AND2X2_68 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_713_) );
OAI21X1 OAI21X1_70 ( .A(_712_), .B(_713_), .C(w_C_57_), .Y(_714_) );
NAND2X1 NAND2X1_120 ( .A(_714_), .B(_718_), .Y(_340__57_) );
INVX1 INVX1_108 ( .A(1'b0), .Y(_722_) );
OR2X2 OR2X2_59 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_723_) );
NAND2X1 NAND2X1_121 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_724_) );
NAND3X1 NAND3X1_77 ( .A(_722_), .B(_724_), .C(_723_), .Y(_725_) );
NOR2X1 NOR2X1_78 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_719_) );
AND2X2 AND2X2_69 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_720_) );
OAI21X1 OAI21X1_71 ( .A(_719_), .B(_720_), .C(1'b0), .Y(_721_) );
NAND2X1 NAND2X1_122 ( .A(_721_), .B(_725_), .Y(_340__0_) );
INVX1 INVX1_109 ( .A(w_C_1_), .Y(_729_) );
OR2X2 OR2X2_60 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_730_) );
NAND2X1 NAND2X1_123 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_731_) );
NAND3X1 NAND3X1_78 ( .A(_729_), .B(_731_), .C(_730_), .Y(_732_) );
NOR2X1 NOR2X1_79 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_726_) );
AND2X2 AND2X2_70 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_727_) );
OAI21X1 OAI21X1_72 ( .A(_726_), .B(_727_), .C(w_C_1_), .Y(_728_) );
NAND2X1 NAND2X1_124 ( .A(_728_), .B(_732_), .Y(_340__1_) );
INVX1 INVX1_110 ( .A(w_C_2_), .Y(_736_) );
OR2X2 OR2X2_61 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_737_) );
NAND2X1 NAND2X1_125 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_738_) );
NAND3X1 NAND3X1_79 ( .A(_736_), .B(_738_), .C(_737_), .Y(_739_) );
NOR2X1 NOR2X1_80 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_733_) );
AND2X2 AND2X2_71 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_734_) );
OAI21X1 OAI21X1_73 ( .A(_733_), .B(_734_), .C(w_C_2_), .Y(_735_) );
NAND2X1 NAND2X1_126 ( .A(_735_), .B(_739_), .Y(_340__2_) );
INVX1 INVX1_111 ( .A(w_C_3_), .Y(_743_) );
OR2X2 OR2X2_62 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_744_) );
NAND2X1 NAND2X1_127 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_745_) );
NAND3X1 NAND3X1_80 ( .A(_743_), .B(_745_), .C(_744_), .Y(_746_) );
NOR2X1 NOR2X1_81 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_740_) );
AND2X2 AND2X2_72 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_741_) );
OAI21X1 OAI21X1_74 ( .A(_740_), .B(_741_), .C(w_C_3_), .Y(_742_) );
NAND2X1 NAND2X1_128 ( .A(_742_), .B(_746_), .Y(_340__3_) );
NOR2X1 NOR2X1_82 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_90_) );
INVX1 INVX1_112 ( .A(_90_), .Y(_91_) );
NOR2X1 NOR2X1_83 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_92_) );
INVX1 INVX1_113 ( .A(_92_), .Y(_93_) );
NAND3X1 NAND3X1_81 ( .A(_91_), .B(_93_), .C(_86_), .Y(_94_) );
OAI21X1 OAI21X1_75 ( .A(_88_), .B(_89_), .C(_94_), .Y(w_C_18_) );
NOR2X1 NOR2X1_84 ( .A(_88_), .B(_89_), .Y(_95_) );
INVX1 INVX1_114 ( .A(_95_), .Y(_96_) );
AND2X2 AND2X2_73 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_97_) );
INVX1 INVX1_115 ( .A(_97_), .Y(_98_) );
NAND3X1 NAND3X1_82 ( .A(_96_), .B(_98_), .C(_94_), .Y(_99_) );
OAI21X1 OAI21X1_76 ( .A(i_add2[18]), .B(i_add1[18]), .C(_99_), .Y(_100_) );
INVX1 INVX1_116 ( .A(_100_), .Y(w_C_19_) );
INVX1 INVX1_117 ( .A(i_add2[19]), .Y(_101_) );
INVX1 INVX1_118 ( .A(i_add1[19]), .Y(_102_) );
NOR2X1 NOR2X1_85 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_103_) );
INVX1 INVX1_119 ( .A(_103_), .Y(_104_) );
NOR2X1 NOR2X1_86 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_105_) );
INVX1 INVX1_120 ( .A(_105_), .Y(_106_) );
NAND3X1 NAND3X1_83 ( .A(_104_), .B(_106_), .C(_99_), .Y(_107_) );
OAI21X1 OAI21X1_77 ( .A(_101_), .B(_102_), .C(_107_), .Y(w_C_20_) );
NOR2X1 NOR2X1_87 ( .A(_101_), .B(_102_), .Y(_108_) );
INVX1 INVX1_121 ( .A(_108_), .Y(_109_) );
AND2X2 AND2X2_74 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_110_) );
INVX1 INVX1_122 ( .A(_110_), .Y(_111_) );
NAND3X1 NAND3X1_84 ( .A(_109_), .B(_111_), .C(_107_), .Y(_112_) );
OAI21X1 OAI21X1_78 ( .A(i_add2[20]), .B(i_add1[20]), .C(_112_), .Y(_113_) );
INVX1 INVX1_123 ( .A(_113_), .Y(w_C_21_) );
INVX1 INVX1_124 ( .A(i_add2[21]), .Y(_114_) );
INVX1 INVX1_125 ( .A(i_add1[21]), .Y(_115_) );
NOR2X1 NOR2X1_88 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_116_) );
INVX1 INVX1_126 ( .A(_116_), .Y(_117_) );
NOR2X1 NOR2X1_89 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_118_) );
INVX1 INVX1_127 ( .A(_118_), .Y(_119_) );
NAND3X1 NAND3X1_85 ( .A(_117_), .B(_119_), .C(_112_), .Y(_120_) );
OAI21X1 OAI21X1_79 ( .A(_114_), .B(_115_), .C(_120_), .Y(w_C_22_) );
NOR2X1 NOR2X1_90 ( .A(_114_), .B(_115_), .Y(_121_) );
INVX1 INVX1_128 ( .A(_121_), .Y(_122_) );
AND2X2 AND2X2_75 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_123_) );
INVX1 INVX1_129 ( .A(_123_), .Y(_124_) );
NAND3X1 NAND3X1_86 ( .A(_122_), .B(_124_), .C(_120_), .Y(_125_) );
OAI21X1 OAI21X1_80 ( .A(i_add2[22]), .B(i_add1[22]), .C(_125_), .Y(_126_) );
INVX1 INVX1_130 ( .A(_126_), .Y(w_C_23_) );
INVX1 INVX1_131 ( .A(i_add2[23]), .Y(_127_) );
INVX1 INVX1_132 ( .A(i_add1[23]), .Y(_128_) );
NOR2X1 NOR2X1_91 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_129_) );
INVX1 INVX1_133 ( .A(_129_), .Y(_130_) );
NOR2X1 NOR2X1_92 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_131_) );
INVX1 INVX1_134 ( .A(_131_), .Y(_132_) );
NAND3X1 NAND3X1_87 ( .A(_130_), .B(_132_), .C(_125_), .Y(_133_) );
OAI21X1 OAI21X1_81 ( .A(_127_), .B(_128_), .C(_133_), .Y(w_C_24_) );
NOR2X1 NOR2X1_93 ( .A(_127_), .B(_128_), .Y(_134_) );
INVX1 INVX1_135 ( .A(_134_), .Y(_135_) );
AND2X2 AND2X2_76 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_136_) );
INVX1 INVX1_136 ( .A(_136_), .Y(_137_) );
NAND3X1 NAND3X1_88 ( .A(_135_), .B(_137_), .C(_133_), .Y(_138_) );
OAI21X1 OAI21X1_82 ( .A(i_add2[24]), .B(i_add1[24]), .C(_138_), .Y(_139_) );
INVX1 INVX1_137 ( .A(_139_), .Y(w_C_25_) );
INVX1 INVX1_138 ( .A(i_add2[25]), .Y(_140_) );
INVX1 INVX1_139 ( .A(i_add1[25]), .Y(_141_) );
NOR2X1 NOR2X1_94 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_142_) );
INVX1 INVX1_140 ( .A(_142_), .Y(_143_) );
NOR2X1 NOR2X1_95 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_144_) );
INVX1 INVX1_141 ( .A(_144_), .Y(_145_) );
NAND3X1 NAND3X1_89 ( .A(_143_), .B(_145_), .C(_138_), .Y(_146_) );
OAI21X1 OAI21X1_83 ( .A(_140_), .B(_141_), .C(_146_), .Y(w_C_26_) );
NOR2X1 NOR2X1_96 ( .A(_140_), .B(_141_), .Y(_147_) );
INVX1 INVX1_142 ( .A(_147_), .Y(_148_) );
AND2X2 AND2X2_77 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_149_) );
INVX1 INVX1_143 ( .A(_149_), .Y(_150_) );
NAND3X1 NAND3X1_90 ( .A(_148_), .B(_150_), .C(_146_), .Y(_151_) );
OAI21X1 OAI21X1_84 ( .A(i_add2[26]), .B(i_add1[26]), .C(_151_), .Y(_152_) );
INVX1 INVX1_144 ( .A(_152_), .Y(w_C_27_) );
INVX1 INVX1_145 ( .A(i_add2[27]), .Y(_153_) );
INVX1 INVX1_146 ( .A(i_add1[27]), .Y(_154_) );
NOR2X1 NOR2X1_97 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_155_) );
INVX1 INVX1_147 ( .A(_155_), .Y(_156_) );
NOR2X1 NOR2X1_98 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_157_) );
INVX1 INVX1_148 ( .A(_157_), .Y(_158_) );
NAND3X1 NAND3X1_91 ( .A(_156_), .B(_158_), .C(_151_), .Y(_159_) );
OAI21X1 OAI21X1_85 ( .A(_153_), .B(_154_), .C(_159_), .Y(w_C_28_) );
NOR2X1 NOR2X1_99 ( .A(_153_), .B(_154_), .Y(_160_) );
INVX1 INVX1_149 ( .A(_160_), .Y(_161_) );
AND2X2 AND2X2_78 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_162_) );
INVX1 INVX1_150 ( .A(_162_), .Y(_163_) );
NAND3X1 NAND3X1_92 ( .A(_161_), .B(_163_), .C(_159_), .Y(_164_) );
OAI21X1 OAI21X1_86 ( .A(i_add2[28]), .B(i_add1[28]), .C(_164_), .Y(_165_) );
INVX1 INVX1_151 ( .A(_165_), .Y(w_C_29_) );
INVX1 INVX1_152 ( .A(i_add2[29]), .Y(_166_) );
INVX1 INVX1_153 ( .A(i_add1[29]), .Y(_167_) );
NOR2X1 NOR2X1_100 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_168_) );
INVX1 INVX1_154 ( .A(_168_), .Y(_169_) );
NOR2X1 NOR2X1_101 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_170_) );
INVX1 INVX1_155 ( .A(_170_), .Y(_171_) );
NAND3X1 NAND3X1_93 ( .A(_169_), .B(_171_), .C(_164_), .Y(_172_) );
OAI21X1 OAI21X1_87 ( .A(_166_), .B(_167_), .C(_172_), .Y(w_C_30_) );
NOR2X1 NOR2X1_102 ( .A(_166_), .B(_167_), .Y(_173_) );
INVX1 INVX1_156 ( .A(_173_), .Y(_174_) );
AND2X2 AND2X2_79 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_175_) );
INVX1 INVX1_157 ( .A(_175_), .Y(_176_) );
NAND3X1 NAND3X1_94 ( .A(_174_), .B(_176_), .C(_172_), .Y(_177_) );
OAI21X1 OAI21X1_88 ( .A(i_add2[30]), .B(i_add1[30]), .C(_177_), .Y(_178_) );
INVX1 INVX1_158 ( .A(_178_), .Y(w_C_31_) );
INVX1 INVX1_159 ( .A(i_add2[31]), .Y(_179_) );
INVX1 INVX1_160 ( .A(i_add1[31]), .Y(_180_) );
NOR2X1 NOR2X1_103 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_181_) );
INVX1 INVX1_161 ( .A(_181_), .Y(_182_) );
NOR2X1 NOR2X1_104 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_183_) );
INVX1 INVX1_162 ( .A(_183_), .Y(_184_) );
NAND3X1 NAND3X1_95 ( .A(_182_), .B(_184_), .C(_177_), .Y(_185_) );
OAI21X1 OAI21X1_89 ( .A(_179_), .B(_180_), .C(_185_), .Y(w_C_32_) );
NOR2X1 NOR2X1_105 ( .A(_179_), .B(_180_), .Y(_186_) );
INVX1 INVX1_163 ( .A(_186_), .Y(_187_) );
AND2X2 AND2X2_80 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_188_) );
INVX1 INVX1_164 ( .A(_188_), .Y(_189_) );
NAND3X1 NAND3X1_96 ( .A(_187_), .B(_189_), .C(_185_), .Y(_190_) );
OAI21X1 OAI21X1_90 ( .A(i_add2[32]), .B(i_add1[32]), .C(_190_), .Y(_191_) );
INVX1 INVX1_165 ( .A(_191_), .Y(w_C_33_) );
INVX1 INVX1_166 ( .A(i_add2[33]), .Y(_192_) );
INVX1 INVX1_167 ( .A(i_add1[33]), .Y(_193_) );
NOR2X1 NOR2X1_106 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_194_) );
INVX1 INVX1_168 ( .A(_194_), .Y(_195_) );
NOR2X1 NOR2X1_107 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_196_) );
INVX1 INVX1_169 ( .A(_196_), .Y(_197_) );
NAND3X1 NAND3X1_97 ( .A(_195_), .B(_197_), .C(_190_), .Y(_198_) );
OAI21X1 OAI21X1_91 ( .A(_192_), .B(_193_), .C(_198_), .Y(w_C_34_) );
NOR2X1 NOR2X1_108 ( .A(_192_), .B(_193_), .Y(_199_) );
INVX1 INVX1_170 ( .A(_199_), .Y(_200_) );
AND2X2 AND2X2_81 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_201_) );
INVX1 INVX1_171 ( .A(_201_), .Y(_202_) );
NAND3X1 NAND3X1_98 ( .A(_200_), .B(_202_), .C(_198_), .Y(_203_) );
OAI21X1 OAI21X1_92 ( .A(i_add2[34]), .B(i_add1[34]), .C(_203_), .Y(_204_) );
INVX1 INVX1_172 ( .A(_204_), .Y(w_C_35_) );
INVX1 INVX1_173 ( .A(i_add2[35]), .Y(_205_) );
INVX1 INVX1_174 ( .A(i_add1[35]), .Y(_206_) );
NOR2X1 NOR2X1_109 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_207_) );
INVX1 INVX1_175 ( .A(_207_), .Y(_208_) );
NOR2X1 NOR2X1_110 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_209_) );
INVX1 INVX1_176 ( .A(_209_), .Y(_210_) );
NAND3X1 NAND3X1_99 ( .A(_208_), .B(_210_), .C(_203_), .Y(_211_) );
OAI21X1 OAI21X1_93 ( .A(_205_), .B(_206_), .C(_211_), .Y(w_C_36_) );
NOR2X1 NOR2X1_111 ( .A(_205_), .B(_206_), .Y(_212_) );
INVX1 INVX1_177 ( .A(_212_), .Y(_213_) );
AND2X2 AND2X2_82 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_214_) );
INVX1 INVX1_178 ( .A(_214_), .Y(_215_) );
NAND3X1 NAND3X1_100 ( .A(_213_), .B(_215_), .C(_211_), .Y(_216_) );
OAI21X1 OAI21X1_94 ( .A(i_add2[36]), .B(i_add1[36]), .C(_216_), .Y(_217_) );
INVX1 INVX1_179 ( .A(_217_), .Y(w_C_37_) );
INVX1 INVX1_180 ( .A(i_add2[37]), .Y(_218_) );
INVX1 INVX1_181 ( .A(i_add1[37]), .Y(_219_) );
NOR2X1 NOR2X1_112 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_220_) );
INVX1 INVX1_182 ( .A(_220_), .Y(_221_) );
NOR2X1 NOR2X1_113 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_222_) );
INVX1 INVX1_183 ( .A(_222_), .Y(_223_) );
NAND3X1 NAND3X1_101 ( .A(_221_), .B(_223_), .C(_216_), .Y(_224_) );
OAI21X1 OAI21X1_95 ( .A(_218_), .B(_219_), .C(_224_), .Y(w_C_38_) );
NOR2X1 NOR2X1_114 ( .A(_218_), .B(_219_), .Y(_225_) );
INVX1 INVX1_184 ( .A(_225_), .Y(_226_) );
AND2X2 AND2X2_83 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_227_) );
INVX1 INVX1_185 ( .A(_227_), .Y(_228_) );
NAND3X1 NAND3X1_102 ( .A(_226_), .B(_228_), .C(_224_), .Y(_229_) );
OAI21X1 OAI21X1_96 ( .A(i_add2[38]), .B(i_add1[38]), .C(_229_), .Y(_230_) );
INVX1 INVX1_186 ( .A(_230_), .Y(w_C_39_) );
INVX1 INVX1_187 ( .A(i_add2[39]), .Y(_231_) );
INVX1 INVX1_188 ( .A(i_add1[39]), .Y(_232_) );
NOR2X1 NOR2X1_115 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_233_) );
INVX1 INVX1_189 ( .A(_233_), .Y(_234_) );
NOR2X1 NOR2X1_116 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_235_) );
INVX1 INVX1_190 ( .A(_235_), .Y(_236_) );
NAND3X1 NAND3X1_103 ( .A(_234_), .B(_236_), .C(_229_), .Y(_237_) );
OAI21X1 OAI21X1_97 ( .A(_231_), .B(_232_), .C(_237_), .Y(w_C_40_) );
NOR2X1 NOR2X1_117 ( .A(_231_), .B(_232_), .Y(_238_) );
INVX1 INVX1_191 ( .A(_238_), .Y(_239_) );
AND2X2 AND2X2_84 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_240_) );
INVX1 INVX1_192 ( .A(_240_), .Y(_241_) );
NAND3X1 NAND3X1_104 ( .A(_239_), .B(_241_), .C(_237_), .Y(_242_) );
OAI21X1 OAI21X1_98 ( .A(i_add2[40]), .B(i_add1[40]), .C(_242_), .Y(_243_) );
INVX1 INVX1_193 ( .A(_243_), .Y(w_C_41_) );
INVX1 INVX1_194 ( .A(i_add2[41]), .Y(_244_) );
INVX1 INVX1_195 ( .A(i_add1[41]), .Y(_245_) );
NOR2X1 NOR2X1_118 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_246_) );
INVX1 INVX1_196 ( .A(_246_), .Y(_247_) );
NOR2X1 NOR2X1_119 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_248_) );
INVX1 INVX1_197 ( .A(_248_), .Y(_249_) );
NAND3X1 NAND3X1_105 ( .A(_247_), .B(_249_), .C(_242_), .Y(_250_) );
OAI21X1 OAI21X1_99 ( .A(_244_), .B(_245_), .C(_250_), .Y(w_C_42_) );
NOR2X1 NOR2X1_120 ( .A(_244_), .B(_245_), .Y(_251_) );
INVX1 INVX1_198 ( .A(_251_), .Y(_252_) );
AND2X2 AND2X2_85 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_253_) );
INVX1 INVX1_199 ( .A(_253_), .Y(_254_) );
NAND3X1 NAND3X1_106 ( .A(_252_), .B(_254_), .C(_250_), .Y(_255_) );
OAI21X1 OAI21X1_100 ( .A(i_add2[42]), .B(i_add1[42]), .C(_255_), .Y(_256_) );
INVX1 INVX1_200 ( .A(_256_), .Y(w_C_43_) );
INVX1 INVX1_201 ( .A(i_add2[43]), .Y(_257_) );
INVX1 INVX1_202 ( .A(i_add1[43]), .Y(_258_) );
NOR2X1 NOR2X1_121 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_259_) );
INVX1 INVX1_203 ( .A(_259_), .Y(_260_) );
NOR2X1 NOR2X1_122 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_261_) );
INVX1 INVX1_204 ( .A(_261_), .Y(_262_) );
NAND3X1 NAND3X1_107 ( .A(_260_), .B(_262_), .C(_255_), .Y(_263_) );
OAI21X1 OAI21X1_101 ( .A(_257_), .B(_258_), .C(_263_), .Y(w_C_44_) );
NOR2X1 NOR2X1_123 ( .A(_257_), .B(_258_), .Y(_264_) );
INVX1 INVX1_205 ( .A(_264_), .Y(_265_) );
AND2X2 AND2X2_86 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_266_) );
INVX1 INVX1_206 ( .A(_266_), .Y(_267_) );
NAND3X1 NAND3X1_108 ( .A(_265_), .B(_267_), .C(_263_), .Y(_268_) );
OAI21X1 OAI21X1_102 ( .A(i_add2[44]), .B(i_add1[44]), .C(_268_), .Y(_269_) );
INVX1 INVX1_207 ( .A(_269_), .Y(w_C_45_) );
INVX1 INVX1_208 ( .A(i_add2[45]), .Y(_270_) );
INVX1 INVX1_209 ( .A(i_add1[45]), .Y(_271_) );
NOR2X1 NOR2X1_124 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_272_) );
INVX1 INVX1_210 ( .A(_272_), .Y(_273_) );
NOR2X1 NOR2X1_125 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_274_) );
INVX1 INVX1_211 ( .A(_274_), .Y(_275_) );
NAND3X1 NAND3X1_109 ( .A(_273_), .B(_275_), .C(_268_), .Y(_276_) );
OAI21X1 OAI21X1_103 ( .A(_270_), .B(_271_), .C(_276_), .Y(w_C_46_) );
NOR2X1 NOR2X1_126 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_277_) );
INVX1 INVX1_212 ( .A(_277_), .Y(_278_) );
NOR2X1 NOR2X1_127 ( .A(_270_), .B(_271_), .Y(_279_) );
INVX1 INVX1_213 ( .A(_279_), .Y(_280_) );
NAND2X1 NAND2X1_129 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_281_) );
NAND3X1 NAND3X1_110 ( .A(_280_), .B(_281_), .C(_276_), .Y(_282_) );
AND2X2 AND2X2_87 ( .A(_282_), .B(_278_), .Y(w_C_47_) );
INVX1 INVX1_214 ( .A(i_add2[47]), .Y(_283_) );
INVX1 INVX1_215 ( .A(i_add1[47]), .Y(_284_) );
NAND2X1 NAND2X1_130 ( .A(_283_), .B(_284_), .Y(_285_) );
NAND3X1 NAND3X1_111 ( .A(_278_), .B(_285_), .C(_282_), .Y(_286_) );
OAI21X1 OAI21X1_104 ( .A(_283_), .B(_284_), .C(_286_), .Y(w_C_48_) );
INVX1 INVX1_216 ( .A(i_add2[48]), .Y(_287_) );
INVX1 INVX1_217 ( .A(i_add1[48]), .Y(_288_) );
OAI21X1 OAI21X1_105 ( .A(i_add2[48]), .B(i_add1[48]), .C(w_C_48_), .Y(_289_) );
OAI21X1 OAI21X1_106 ( .A(_287_), .B(_288_), .C(_289_), .Y(w_C_49_) );
INVX1 INVX1_218 ( .A(i_add2[49]), .Y(_290_) );
INVX1 INVX1_219 ( .A(i_add1[49]), .Y(_291_) );
NOR2X1 NOR2X1_128 ( .A(_290_), .B(_291_), .Y(_292_) );
OR2X2 OR2X2_63 ( .A(w_C_49_), .B(_292_), .Y(_293_) );
OAI21X1 OAI21X1_107 ( .A(i_add2[49]), .B(i_add1[49]), .C(_293_), .Y(_294_) );
INVX1 INVX1_220 ( .A(_294_), .Y(w_C_50_) );
NAND2X1 NAND2X1_131 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_295_) );
NOR2X1 NOR2X1_129 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_296_) );
OAI21X1 OAI21X1_108 ( .A(_296_), .B(_294_), .C(_295_), .Y(w_C_51_) );
INVX1 INVX1_221 ( .A(i_add2[51]), .Y(_297_) );
INVX1 INVX1_222 ( .A(i_add1[51]), .Y(_298_) );
INVX1 INVX1_223 ( .A(_296_), .Y(_299_) );
INVX1 INVX1_224 ( .A(_292_), .Y(_300_) );
NAND2X1 NAND2X1_132 ( .A(_287_), .B(_288_), .Y(_301_) );
NAND2X1 NAND2X1_133 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_302_) );
NAND2X1 NAND2X1_134 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_303_) );
NAND3X1 NAND3X1_112 ( .A(_302_), .B(_303_), .C(_286_), .Y(_304_) );
NAND2X1 NAND2X1_135 ( .A(_290_), .B(_291_), .Y(_305_) );
NAND3X1 NAND3X1_113 ( .A(_301_), .B(_305_), .C(_304_), .Y(_306_) );
NAND3X1 NAND3X1_114 ( .A(_300_), .B(_295_), .C(_306_), .Y(_307_) );
NAND2X1 NAND2X1_136 ( .A(_297_), .B(_298_), .Y(_308_) );
BUFX2 BUFX2_60 ( .A(w_C_58_), .Y(_340__58_) );
BUFX2 BUFX2_61 ( .A(1'b0), .Y(w_C_0_) );
endmodule
