module csa_31bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [30:0] i_add_term1;
input [30:0] i_add_term2;
output [30:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

NOR2X1 NOR2X1_1 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_398_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_399_) );
OAI21X1 OAI21X1_1 ( .A(_398_), .B(_399_), .C(_35__2_), .Y(_400_) );
NAND2X1 NAND2X1_1 ( .A(_400_), .B(_404_), .Y(_33__2_) );
OAI21X1 OAI21X1_2 ( .A(_401_), .B(_398_), .C(_403_), .Y(_35__3_) );
INVX1 INVX1_1 ( .A(vdd), .Y(_408_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_409_) );
NAND2X1 NAND2X1_2 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_410_) );
NAND3X1 NAND3X1_1 ( .A(_408_), .B(_410_), .C(_409_), .Y(_411_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_405_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_406_) );
OAI21X1 OAI21X1_3 ( .A(_405_), .B(_406_), .C(vdd), .Y(_407_) );
NAND2X1 NAND2X1_3 ( .A(_407_), .B(_411_), .Y(_34__0_) );
OAI21X1 OAI21X1_4 ( .A(_408_), .B(_405_), .C(_410_), .Y(_36__1_) );
INVX1 INVX1_2 ( .A(_36__3_), .Y(_415_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_416_) );
NAND2X1 NAND2X1_4 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_417_) );
NAND3X1 NAND3X1_2 ( .A(_415_), .B(_417_), .C(_416_), .Y(_418_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_412_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_413_) );
OAI21X1 OAI21X1_5 ( .A(_412_), .B(_413_), .C(_36__3_), .Y(_414_) );
NAND2X1 NAND2X1_5 ( .A(_414_), .B(_418_), .Y(_34__3_) );
OAI21X1 OAI21X1_6 ( .A(_415_), .B(_412_), .C(_417_), .Y(_32_) );
INVX1 INVX1_3 ( .A(_36__1_), .Y(_422_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_423_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_424_) );
NAND3X1 NAND3X1_3 ( .A(_422_), .B(_424_), .C(_423_), .Y(_425_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_419_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_420_) );
OAI21X1 OAI21X1_7 ( .A(_419_), .B(_420_), .C(_36__1_), .Y(_421_) );
NAND2X1 NAND2X1_7 ( .A(_421_), .B(_425_), .Y(_34__1_) );
OAI21X1 OAI21X1_8 ( .A(_422_), .B(_419_), .C(_424_), .Y(_36__2_) );
INVX1 INVX1_4 ( .A(_36__2_), .Y(_429_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_430_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_431_) );
NAND3X1 NAND3X1_4 ( .A(_429_), .B(_431_), .C(_430_), .Y(_432_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_426_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_427_) );
OAI21X1 OAI21X1_9 ( .A(_426_), .B(_427_), .C(_36__2_), .Y(_428_) );
NAND2X1 NAND2X1_9 ( .A(_428_), .B(_432_), .Y(_34__2_) );
OAI21X1 OAI21X1_10 ( .A(_429_), .B(_426_), .C(_431_), .Y(_36__3_) );
INVX1 INVX1_5 ( .A(csa_inst_cout0_0), .Y(_433_) );
NAND2X1 NAND2X1_10 ( .A(csa_inst_cout0_1), .B(csa_inst_cin), .Y(_434_) );
OAI21X1 OAI21X1_11 ( .A(csa_inst_cin), .B(_433_), .C(_434_), .Y(w_cout_7_) );
INVX1 INVX1_6 ( .A(gnd), .Y(_436_) );
NAND2X1 NAND2X1_11 ( .A(gnd), .B(gnd), .Y(_437_) );
NOR2X1 NOR2X1_6 ( .A(gnd), .B(gnd), .Y(_435_) );
OAI21X1 OAI21X1_12 ( .A(_436_), .B(_435_), .C(_437_), .Y(csa_inst_rca0_0_fa0_o_carry) );
INVX1 INVX1_7 ( .A(csa_inst_rca0_0_fa31_i_carry), .Y(_439_) );
NAND2X1 NAND2X1_12 ( .A(gnd), .B(gnd), .Y(_440_) );
NOR2X1 NOR2X1_7 ( .A(gnd), .B(gnd), .Y(_438_) );
OAI21X1 OAI21X1_13 ( .A(_439_), .B(_438_), .C(_440_), .Y(csa_inst_cout0_0) );
INVX1 INVX1_8 ( .A(csa_inst_rca0_0_fa0_o_carry), .Y(_442_) );
NAND2X1 NAND2X1_13 ( .A(gnd), .B(gnd), .Y(_443_) );
NOR2X1 NOR2X1_8 ( .A(gnd), .B(gnd), .Y(_441_) );
OAI21X1 OAI21X1_14 ( .A(_442_), .B(_441_), .C(_443_), .Y(csa_inst_rca0_0_fa_1__o_carry) );
INVX1 INVX1_9 ( .A(csa_inst_rca0_0_fa_1__o_carry), .Y(_445_) );
NAND2X1 NAND2X1_14 ( .A(gnd), .B(gnd), .Y(_446_) );
NOR2X1 NOR2X1_9 ( .A(gnd), .B(gnd), .Y(_444_) );
OAI21X1 OAI21X1_15 ( .A(_445_), .B(_444_), .C(_446_), .Y(csa_inst_rca0_0_fa31_i_carry) );
INVX1 INVX1_10 ( .A(vdd), .Y(_448_) );
NAND2X1 NAND2X1_15 ( .A(gnd), .B(gnd), .Y(_449_) );
NOR2X1 NOR2X1_10 ( .A(gnd), .B(gnd), .Y(_447_) );
OAI21X1 OAI21X1_16 ( .A(_448_), .B(_447_), .C(_449_), .Y(csa_inst_rca0_1_fa0_o_carry) );
INVX1 INVX1_11 ( .A(csa_inst_rca0_1_fa31_i_carry), .Y(_451_) );
NAND2X1 NAND2X1_16 ( .A(gnd), .B(gnd), .Y(_452_) );
NOR2X1 NOR2X1_11 ( .A(gnd), .B(gnd), .Y(_450_) );
OAI21X1 OAI21X1_17 ( .A(_451_), .B(_450_), .C(_452_), .Y(csa_inst_cout0_1) );
INVX1 INVX1_12 ( .A(csa_inst_rca0_1_fa0_o_carry), .Y(_454_) );
NAND2X1 NAND2X1_17 ( .A(gnd), .B(gnd), .Y(_455_) );
NOR2X1 NOR2X1_12 ( .A(gnd), .B(gnd), .Y(_453_) );
OAI21X1 OAI21X1_18 ( .A(_454_), .B(_453_), .C(_455_), .Y(csa_inst_rca0_1_fa_1__o_carry) );
INVX1 INVX1_13 ( .A(csa_inst_rca0_1_fa_1__o_carry), .Y(_457_) );
NAND2X1 NAND2X1_18 ( .A(gnd), .B(gnd), .Y(_458_) );
NOR2X1 NOR2X1_13 ( .A(gnd), .B(gnd), .Y(_456_) );
OAI21X1 OAI21X1_19 ( .A(_457_), .B(_456_), .C(_458_), .Y(csa_inst_rca0_1_fa31_i_carry) );
INVX1 INVX1_14 ( .A(gnd), .Y(_462_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_463_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_464_) );
NAND3X1 NAND3X1_5 ( .A(_462_), .B(_464_), .C(_463_), .Y(_465_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_459_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_460_) );
OAI21X1 OAI21X1_20 ( .A(_459_), .B(_460_), .C(gnd), .Y(_461_) );
NAND2X1 NAND2X1_20 ( .A(_461_), .B(_465_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_21 ( .A(_462_), .B(_459_), .C(_464_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_15 ( .A(rca_inst_fa31_i_carry), .Y(_469_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_470_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_471_) );
NAND3X1 NAND3X1_6 ( .A(_469_), .B(_471_), .C(_470_), .Y(_472_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_466_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_467_) );
OAI21X1 OAI21X1_22 ( .A(_466_), .B(_467_), .C(rca_inst_fa31_i_carry), .Y(_468_) );
NAND2X1 NAND2X1_22 ( .A(_468_), .B(_472_), .Y(rca_inst_fa31_o_sum) );
OAI21X1 OAI21X1_23 ( .A(_469_), .B(_466_), .C(_471_), .Y(rca_inst_cout) );
INVX1 INVX1_16 ( .A(rca_inst_fa0_o_carry), .Y(_476_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_477_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_478_) );
NAND3X1 NAND3X1_7 ( .A(_476_), .B(_478_), .C(_477_), .Y(_479_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_473_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_474_) );
OAI21X1 OAI21X1_24 ( .A(_473_), .B(_474_), .C(rca_inst_fa0_o_carry), .Y(_475_) );
NAND2X1 NAND2X1_24 ( .A(_475_), .B(_479_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_25 ( .A(_476_), .B(_473_), .C(_478_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_17 ( .A(rca_inst_fa_1__o_carry), .Y(_483_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_484_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_485_) );
NAND3X1 NAND3X1_8 ( .A(_483_), .B(_485_), .C(_484_), .Y(_486_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_480_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_481_) );
OAI21X1 OAI21X1_26 ( .A(_480_), .B(_481_), .C(rca_inst_fa_1__o_carry), .Y(_482_) );
NAND2X1 NAND2X1_26 ( .A(_482_), .B(_486_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_27 ( .A(_483_), .B(_480_), .C(_485_), .Y(rca_inst_fa31_i_carry) );
BUFX2 BUFX2_1 ( .A(w_cout_7_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa31_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(gnd), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(gnd), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(gnd), .Y(sum[30]) );
INVX1 INVX1_18 ( .A(_1_), .Y(_37_) );
NAND2X1 NAND2X1_27 ( .A(_2_), .B(rca_inst_cout), .Y(_38_) );
OAI21X1 OAI21X1_28 ( .A(rca_inst_cout), .B(_37_), .C(_38_), .Y(w_cout_1_) );
INVX1 INVX1_19 ( .A(_3__0_), .Y(_39_) );
NAND2X1 NAND2X1_28 ( .A(_4__0_), .B(rca_inst_cout), .Y(_40_) );
OAI21X1 OAI21X1_29 ( .A(rca_inst_cout), .B(_39_), .C(_40_), .Y(_0__4_) );
INVX1 INVX1_20 ( .A(_3__1_), .Y(_41_) );
NAND2X1 NAND2X1_29 ( .A(rca_inst_cout), .B(_4__1_), .Y(_42_) );
OAI21X1 OAI21X1_30 ( .A(rca_inst_cout), .B(_41_), .C(_42_), .Y(_0__5_) );
INVX1 INVX1_21 ( .A(_3__2_), .Y(_43_) );
NAND2X1 NAND2X1_30 ( .A(rca_inst_cout), .B(_4__2_), .Y(_44_) );
OAI21X1 OAI21X1_31 ( .A(rca_inst_cout), .B(_43_), .C(_44_), .Y(_0__6_) );
INVX1 INVX1_22 ( .A(_3__3_), .Y(_45_) );
NAND2X1 NAND2X1_31 ( .A(rca_inst_cout), .B(_4__3_), .Y(_46_) );
OAI21X1 OAI21X1_32 ( .A(rca_inst_cout), .B(_45_), .C(_46_), .Y(_0__7_) );
INVX1 INVX1_23 ( .A(gnd), .Y(_50_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_51_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_52_) );
NAND3X1 NAND3X1_9 ( .A(_50_), .B(_52_), .C(_51_), .Y(_53_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_47_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_48_) );
OAI21X1 OAI21X1_33 ( .A(_47_), .B(_48_), .C(gnd), .Y(_49_) );
NAND2X1 NAND2X1_33 ( .A(_49_), .B(_53_), .Y(_3__0_) );
OAI21X1 OAI21X1_34 ( .A(_50_), .B(_47_), .C(_52_), .Y(_5__1_) );
INVX1 INVX1_24 ( .A(_5__3_), .Y(_57_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_58_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_59_) );
NAND3X1 NAND3X1_10 ( .A(_57_), .B(_59_), .C(_58_), .Y(_60_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_54_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_55_) );
OAI21X1 OAI21X1_35 ( .A(_54_), .B(_55_), .C(_5__3_), .Y(_56_) );
NAND2X1 NAND2X1_35 ( .A(_56_), .B(_60_), .Y(_3__3_) );
OAI21X1 OAI21X1_36 ( .A(_57_), .B(_54_), .C(_59_), .Y(_1_) );
INVX1 INVX1_25 ( .A(_5__1_), .Y(_64_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_65_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_66_) );
NAND3X1 NAND3X1_11 ( .A(_64_), .B(_66_), .C(_65_), .Y(_67_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_61_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_62_) );
OAI21X1 OAI21X1_37 ( .A(_61_), .B(_62_), .C(_5__1_), .Y(_63_) );
NAND2X1 NAND2X1_37 ( .A(_63_), .B(_67_), .Y(_3__1_) );
OAI21X1 OAI21X1_38 ( .A(_64_), .B(_61_), .C(_66_), .Y(_5__2_) );
INVX1 INVX1_26 ( .A(_5__2_), .Y(_71_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_72_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_73_) );
NAND3X1 NAND3X1_12 ( .A(_71_), .B(_73_), .C(_72_), .Y(_74_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_68_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_69_) );
OAI21X1 OAI21X1_39 ( .A(_68_), .B(_69_), .C(_5__2_), .Y(_70_) );
NAND2X1 NAND2X1_39 ( .A(_70_), .B(_74_), .Y(_3__2_) );
OAI21X1 OAI21X1_40 ( .A(_71_), .B(_68_), .C(_73_), .Y(_5__3_) );
INVX1 INVX1_27 ( .A(vdd), .Y(_78_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_79_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_80_) );
NAND3X1 NAND3X1_13 ( .A(_78_), .B(_80_), .C(_79_), .Y(_81_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_75_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_76_) );
OAI21X1 OAI21X1_41 ( .A(_75_), .B(_76_), .C(vdd), .Y(_77_) );
NAND2X1 NAND2X1_41 ( .A(_77_), .B(_81_), .Y(_4__0_) );
OAI21X1 OAI21X1_42 ( .A(_78_), .B(_75_), .C(_80_), .Y(_6__1_) );
INVX1 INVX1_28 ( .A(_6__3_), .Y(_85_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_86_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_87_) );
NAND3X1 NAND3X1_14 ( .A(_85_), .B(_87_), .C(_86_), .Y(_88_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_82_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_83_) );
OAI21X1 OAI21X1_43 ( .A(_82_), .B(_83_), .C(_6__3_), .Y(_84_) );
NAND2X1 NAND2X1_43 ( .A(_84_), .B(_88_), .Y(_4__3_) );
OAI21X1 OAI21X1_44 ( .A(_85_), .B(_82_), .C(_87_), .Y(_2_) );
INVX1 INVX1_29 ( .A(_6__1_), .Y(_92_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_93_) );
NAND2X1 NAND2X1_44 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_94_) );
NAND3X1 NAND3X1_15 ( .A(_92_), .B(_94_), .C(_93_), .Y(_95_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_89_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_90_) );
OAI21X1 OAI21X1_45 ( .A(_89_), .B(_90_), .C(_6__1_), .Y(_91_) );
NAND2X1 NAND2X1_45 ( .A(_91_), .B(_95_), .Y(_4__1_) );
OAI21X1 OAI21X1_46 ( .A(_92_), .B(_89_), .C(_94_), .Y(_6__2_) );
INVX1 INVX1_30 ( .A(_6__2_), .Y(_99_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_100_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_101_) );
NAND3X1 NAND3X1_16 ( .A(_99_), .B(_101_), .C(_100_), .Y(_102_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_96_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_97_) );
OAI21X1 OAI21X1_47 ( .A(_96_), .B(_97_), .C(_6__2_), .Y(_98_) );
NAND2X1 NAND2X1_47 ( .A(_98_), .B(_102_), .Y(_4__2_) );
OAI21X1 OAI21X1_48 ( .A(_99_), .B(_96_), .C(_101_), .Y(_6__3_) );
INVX1 INVX1_31 ( .A(_7_), .Y(_103_) );
NAND2X1 NAND2X1_48 ( .A(_8_), .B(w_cout_1_), .Y(_104_) );
OAI21X1 OAI21X1_49 ( .A(w_cout_1_), .B(_103_), .C(_104_), .Y(w_cout_2_) );
INVX1 INVX1_32 ( .A(_9__0_), .Y(_105_) );
NAND2X1 NAND2X1_49 ( .A(_10__0_), .B(w_cout_1_), .Y(_106_) );
OAI21X1 OAI21X1_50 ( .A(w_cout_1_), .B(_105_), .C(_106_), .Y(_0__8_) );
INVX1 INVX1_33 ( .A(_9__1_), .Y(_107_) );
NAND2X1 NAND2X1_50 ( .A(w_cout_1_), .B(_10__1_), .Y(_108_) );
OAI21X1 OAI21X1_51 ( .A(w_cout_1_), .B(_107_), .C(_108_), .Y(_0__9_) );
INVX1 INVX1_34 ( .A(_9__2_), .Y(_109_) );
NAND2X1 NAND2X1_51 ( .A(w_cout_1_), .B(_10__2_), .Y(_110_) );
OAI21X1 OAI21X1_52 ( .A(w_cout_1_), .B(_109_), .C(_110_), .Y(_0__10_) );
INVX1 INVX1_35 ( .A(_9__3_), .Y(_111_) );
NAND2X1 NAND2X1_52 ( .A(w_cout_1_), .B(_10__3_), .Y(_112_) );
OAI21X1 OAI21X1_53 ( .A(w_cout_1_), .B(_111_), .C(_112_), .Y(_0__11_) );
INVX1 INVX1_36 ( .A(gnd), .Y(_116_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_117_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_118_) );
NAND3X1 NAND3X1_17 ( .A(_116_), .B(_118_), .C(_117_), .Y(_119_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_113_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_114_) );
OAI21X1 OAI21X1_54 ( .A(_113_), .B(_114_), .C(gnd), .Y(_115_) );
NAND2X1 NAND2X1_54 ( .A(_115_), .B(_119_), .Y(_9__0_) );
OAI21X1 OAI21X1_55 ( .A(_116_), .B(_113_), .C(_118_), .Y(_11__1_) );
INVX1 INVX1_37 ( .A(_11__3_), .Y(_123_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_124_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_125_) );
NAND3X1 NAND3X1_18 ( .A(_123_), .B(_125_), .C(_124_), .Y(_126_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_120_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_121_) );
OAI21X1 OAI21X1_56 ( .A(_120_), .B(_121_), .C(_11__3_), .Y(_122_) );
NAND2X1 NAND2X1_56 ( .A(_122_), .B(_126_), .Y(_9__3_) );
OAI21X1 OAI21X1_57 ( .A(_123_), .B(_120_), .C(_125_), .Y(_7_) );
INVX1 INVX1_38 ( .A(_11__1_), .Y(_130_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_131_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_132_) );
NAND3X1 NAND3X1_19 ( .A(_130_), .B(_132_), .C(_131_), .Y(_133_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_127_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_128_) );
OAI21X1 OAI21X1_58 ( .A(_127_), .B(_128_), .C(_11__1_), .Y(_129_) );
NAND2X1 NAND2X1_58 ( .A(_129_), .B(_133_), .Y(_9__1_) );
OAI21X1 OAI21X1_59 ( .A(_130_), .B(_127_), .C(_132_), .Y(_11__2_) );
INVX1 INVX1_39 ( .A(_11__2_), .Y(_137_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_138_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_139_) );
NAND3X1 NAND3X1_20 ( .A(_137_), .B(_139_), .C(_138_), .Y(_140_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_134_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_135_) );
OAI21X1 OAI21X1_60 ( .A(_134_), .B(_135_), .C(_11__2_), .Y(_136_) );
NAND2X1 NAND2X1_60 ( .A(_136_), .B(_140_), .Y(_9__2_) );
OAI21X1 OAI21X1_61 ( .A(_137_), .B(_134_), .C(_139_), .Y(_11__3_) );
INVX1 INVX1_40 ( .A(vdd), .Y(_144_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_145_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_146_) );
NAND3X1 NAND3X1_21 ( .A(_144_), .B(_146_), .C(_145_), .Y(_147_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_141_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_142_) );
OAI21X1 OAI21X1_62 ( .A(_141_), .B(_142_), .C(vdd), .Y(_143_) );
NAND2X1 NAND2X1_62 ( .A(_143_), .B(_147_), .Y(_10__0_) );
OAI21X1 OAI21X1_63 ( .A(_144_), .B(_141_), .C(_146_), .Y(_12__1_) );
INVX1 INVX1_41 ( .A(_12__3_), .Y(_151_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_152_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_153_) );
NAND3X1 NAND3X1_22 ( .A(_151_), .B(_153_), .C(_152_), .Y(_154_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_148_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_149_) );
OAI21X1 OAI21X1_64 ( .A(_148_), .B(_149_), .C(_12__3_), .Y(_150_) );
NAND2X1 NAND2X1_64 ( .A(_150_), .B(_154_), .Y(_10__3_) );
OAI21X1 OAI21X1_65 ( .A(_151_), .B(_148_), .C(_153_), .Y(_8_) );
INVX1 INVX1_42 ( .A(_12__1_), .Y(_158_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_159_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_160_) );
NAND3X1 NAND3X1_23 ( .A(_158_), .B(_160_), .C(_159_), .Y(_161_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_155_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_156_) );
OAI21X1 OAI21X1_66 ( .A(_155_), .B(_156_), .C(_12__1_), .Y(_157_) );
NAND2X1 NAND2X1_66 ( .A(_157_), .B(_161_), .Y(_10__1_) );
OAI21X1 OAI21X1_67 ( .A(_158_), .B(_155_), .C(_160_), .Y(_12__2_) );
INVX1 INVX1_43 ( .A(_12__2_), .Y(_165_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_166_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_167_) );
NAND3X1 NAND3X1_24 ( .A(_165_), .B(_167_), .C(_166_), .Y(_168_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_162_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_163_) );
OAI21X1 OAI21X1_68 ( .A(_162_), .B(_163_), .C(_12__2_), .Y(_164_) );
NAND2X1 NAND2X1_68 ( .A(_164_), .B(_168_), .Y(_10__2_) );
OAI21X1 OAI21X1_69 ( .A(_165_), .B(_162_), .C(_167_), .Y(_12__3_) );
INVX1 INVX1_44 ( .A(_13_), .Y(_169_) );
NAND2X1 NAND2X1_69 ( .A(_14_), .B(w_cout_2_), .Y(_170_) );
OAI21X1 OAI21X1_70 ( .A(w_cout_2_), .B(_169_), .C(_170_), .Y(w_cout_3_) );
INVX1 INVX1_45 ( .A(_15__0_), .Y(_171_) );
NAND2X1 NAND2X1_70 ( .A(_16__0_), .B(w_cout_2_), .Y(_172_) );
OAI21X1 OAI21X1_71 ( .A(w_cout_2_), .B(_171_), .C(_172_), .Y(_0__12_) );
INVX1 INVX1_46 ( .A(_15__1_), .Y(_173_) );
NAND2X1 NAND2X1_71 ( .A(w_cout_2_), .B(_16__1_), .Y(_174_) );
OAI21X1 OAI21X1_72 ( .A(w_cout_2_), .B(_173_), .C(_174_), .Y(_0__13_) );
INVX1 INVX1_47 ( .A(_15__2_), .Y(_175_) );
NAND2X1 NAND2X1_72 ( .A(w_cout_2_), .B(_16__2_), .Y(_176_) );
OAI21X1 OAI21X1_73 ( .A(w_cout_2_), .B(_175_), .C(_176_), .Y(_0__14_) );
INVX1 INVX1_48 ( .A(_15__3_), .Y(_177_) );
NAND2X1 NAND2X1_73 ( .A(w_cout_2_), .B(_16__3_), .Y(_178_) );
OAI21X1 OAI21X1_74 ( .A(w_cout_2_), .B(_177_), .C(_178_), .Y(_0__15_) );
INVX1 INVX1_49 ( .A(gnd), .Y(_182_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_183_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_184_) );
NAND3X1 NAND3X1_25 ( .A(_182_), .B(_184_), .C(_183_), .Y(_185_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_179_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_180_) );
OAI21X1 OAI21X1_75 ( .A(_179_), .B(_180_), .C(gnd), .Y(_181_) );
NAND2X1 NAND2X1_75 ( .A(_181_), .B(_185_), .Y(_15__0_) );
OAI21X1 OAI21X1_76 ( .A(_182_), .B(_179_), .C(_184_), .Y(_17__1_) );
INVX1 INVX1_50 ( .A(_17__3_), .Y(_189_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_190_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_191_) );
NAND3X1 NAND3X1_26 ( .A(_189_), .B(_191_), .C(_190_), .Y(_192_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_186_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_187_) );
OAI21X1 OAI21X1_77 ( .A(_186_), .B(_187_), .C(_17__3_), .Y(_188_) );
NAND2X1 NAND2X1_77 ( .A(_188_), .B(_192_), .Y(_15__3_) );
OAI21X1 OAI21X1_78 ( .A(_189_), .B(_186_), .C(_191_), .Y(_13_) );
INVX1 INVX1_51 ( .A(_17__1_), .Y(_196_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_197_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_198_) );
NAND3X1 NAND3X1_27 ( .A(_196_), .B(_198_), .C(_197_), .Y(_199_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_193_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_194_) );
OAI21X1 OAI21X1_79 ( .A(_193_), .B(_194_), .C(_17__1_), .Y(_195_) );
NAND2X1 NAND2X1_79 ( .A(_195_), .B(_199_), .Y(_15__1_) );
OAI21X1 OAI21X1_80 ( .A(_196_), .B(_193_), .C(_198_), .Y(_17__2_) );
INVX1 INVX1_52 ( .A(_17__2_), .Y(_203_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_204_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_205_) );
NAND3X1 NAND3X1_28 ( .A(_203_), .B(_205_), .C(_204_), .Y(_206_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_200_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_201_) );
OAI21X1 OAI21X1_81 ( .A(_200_), .B(_201_), .C(_17__2_), .Y(_202_) );
NAND2X1 NAND2X1_81 ( .A(_202_), .B(_206_), .Y(_15__2_) );
OAI21X1 OAI21X1_82 ( .A(_203_), .B(_200_), .C(_205_), .Y(_17__3_) );
INVX1 INVX1_53 ( .A(vdd), .Y(_210_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_211_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_212_) );
NAND3X1 NAND3X1_29 ( .A(_210_), .B(_212_), .C(_211_), .Y(_213_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_207_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_208_) );
OAI21X1 OAI21X1_83 ( .A(_207_), .B(_208_), .C(vdd), .Y(_209_) );
NAND2X1 NAND2X1_83 ( .A(_209_), .B(_213_), .Y(_16__0_) );
OAI21X1 OAI21X1_84 ( .A(_210_), .B(_207_), .C(_212_), .Y(_18__1_) );
INVX1 INVX1_54 ( .A(_18__3_), .Y(_217_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_218_) );
NAND2X1 NAND2X1_84 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_219_) );
NAND3X1 NAND3X1_30 ( .A(_217_), .B(_219_), .C(_218_), .Y(_220_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_214_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_215_) );
OAI21X1 OAI21X1_85 ( .A(_214_), .B(_215_), .C(_18__3_), .Y(_216_) );
NAND2X1 NAND2X1_85 ( .A(_216_), .B(_220_), .Y(_16__3_) );
OAI21X1 OAI21X1_86 ( .A(_217_), .B(_214_), .C(_219_), .Y(_14_) );
INVX1 INVX1_55 ( .A(_18__1_), .Y(_224_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_225_) );
NAND2X1 NAND2X1_86 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_226_) );
NAND3X1 NAND3X1_31 ( .A(_224_), .B(_226_), .C(_225_), .Y(_227_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_221_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_222_) );
OAI21X1 OAI21X1_87 ( .A(_221_), .B(_222_), .C(_18__1_), .Y(_223_) );
NAND2X1 NAND2X1_87 ( .A(_223_), .B(_227_), .Y(_16__1_) );
OAI21X1 OAI21X1_88 ( .A(_224_), .B(_221_), .C(_226_), .Y(_18__2_) );
INVX1 INVX1_56 ( .A(_18__2_), .Y(_231_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_232_) );
NAND2X1 NAND2X1_88 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_233_) );
NAND3X1 NAND3X1_32 ( .A(_231_), .B(_233_), .C(_232_), .Y(_234_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_228_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_229_) );
OAI21X1 OAI21X1_89 ( .A(_228_), .B(_229_), .C(_18__2_), .Y(_230_) );
NAND2X1 NAND2X1_89 ( .A(_230_), .B(_234_), .Y(_16__2_) );
OAI21X1 OAI21X1_90 ( .A(_231_), .B(_228_), .C(_233_), .Y(_18__3_) );
INVX1 INVX1_57 ( .A(_19_), .Y(_235_) );
NAND2X1 NAND2X1_90 ( .A(_20_), .B(w_cout_3_), .Y(_236_) );
OAI21X1 OAI21X1_91 ( .A(w_cout_3_), .B(_235_), .C(_236_), .Y(w_cout_4_) );
INVX1 INVX1_58 ( .A(_21__0_), .Y(_237_) );
NAND2X1 NAND2X1_91 ( .A(_22__0_), .B(w_cout_3_), .Y(_238_) );
OAI21X1 OAI21X1_92 ( .A(w_cout_3_), .B(_237_), .C(_238_), .Y(_0__16_) );
INVX1 INVX1_59 ( .A(_21__1_), .Y(_239_) );
NAND2X1 NAND2X1_92 ( .A(w_cout_3_), .B(_22__1_), .Y(_240_) );
OAI21X1 OAI21X1_93 ( .A(w_cout_3_), .B(_239_), .C(_240_), .Y(_0__17_) );
INVX1 INVX1_60 ( .A(_21__2_), .Y(_241_) );
NAND2X1 NAND2X1_93 ( .A(w_cout_3_), .B(_22__2_), .Y(_242_) );
OAI21X1 OAI21X1_94 ( .A(w_cout_3_), .B(_241_), .C(_242_), .Y(_0__18_) );
INVX1 INVX1_61 ( .A(_21__3_), .Y(_243_) );
NAND2X1 NAND2X1_94 ( .A(w_cout_3_), .B(_22__3_), .Y(_244_) );
OAI21X1 OAI21X1_95 ( .A(w_cout_3_), .B(_243_), .C(_244_), .Y(_0__19_) );
INVX1 INVX1_62 ( .A(gnd), .Y(_248_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_249_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_250_) );
NAND3X1 NAND3X1_33 ( .A(_248_), .B(_250_), .C(_249_), .Y(_251_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_245_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_246_) );
OAI21X1 OAI21X1_96 ( .A(_245_), .B(_246_), .C(gnd), .Y(_247_) );
NAND2X1 NAND2X1_96 ( .A(_247_), .B(_251_), .Y(_21__0_) );
OAI21X1 OAI21X1_97 ( .A(_248_), .B(_245_), .C(_250_), .Y(_23__1_) );
INVX1 INVX1_63 ( .A(_23__3_), .Y(_255_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_256_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_257_) );
NAND3X1 NAND3X1_34 ( .A(_255_), .B(_257_), .C(_256_), .Y(_258_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_252_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_253_) );
OAI21X1 OAI21X1_98 ( .A(_252_), .B(_253_), .C(_23__3_), .Y(_254_) );
NAND2X1 NAND2X1_98 ( .A(_254_), .B(_258_), .Y(_21__3_) );
OAI21X1 OAI21X1_99 ( .A(_255_), .B(_252_), .C(_257_), .Y(_19_) );
INVX1 INVX1_64 ( .A(_23__1_), .Y(_262_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_263_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_264_) );
NAND3X1 NAND3X1_35 ( .A(_262_), .B(_264_), .C(_263_), .Y(_265_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_259_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_260_) );
OAI21X1 OAI21X1_100 ( .A(_259_), .B(_260_), .C(_23__1_), .Y(_261_) );
NAND2X1 NAND2X1_100 ( .A(_261_), .B(_265_), .Y(_21__1_) );
OAI21X1 OAI21X1_101 ( .A(_262_), .B(_259_), .C(_264_), .Y(_23__2_) );
INVX1 INVX1_65 ( .A(_23__2_), .Y(_269_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_270_) );
NAND2X1 NAND2X1_101 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_271_) );
NAND3X1 NAND3X1_36 ( .A(_269_), .B(_271_), .C(_270_), .Y(_272_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_266_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_267_) );
OAI21X1 OAI21X1_102 ( .A(_266_), .B(_267_), .C(_23__2_), .Y(_268_) );
NAND2X1 NAND2X1_102 ( .A(_268_), .B(_272_), .Y(_21__2_) );
OAI21X1 OAI21X1_103 ( .A(_269_), .B(_266_), .C(_271_), .Y(_23__3_) );
INVX1 INVX1_66 ( .A(vdd), .Y(_276_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_277_) );
NAND2X1 NAND2X1_103 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_278_) );
NAND3X1 NAND3X1_37 ( .A(_276_), .B(_278_), .C(_277_), .Y(_279_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_273_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_274_) );
OAI21X1 OAI21X1_104 ( .A(_273_), .B(_274_), .C(vdd), .Y(_275_) );
NAND2X1 NAND2X1_104 ( .A(_275_), .B(_279_), .Y(_22__0_) );
OAI21X1 OAI21X1_105 ( .A(_276_), .B(_273_), .C(_278_), .Y(_24__1_) );
INVX1 INVX1_67 ( .A(_24__3_), .Y(_283_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_284_) );
NAND2X1 NAND2X1_105 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_285_) );
NAND3X1 NAND3X1_38 ( .A(_283_), .B(_285_), .C(_284_), .Y(_286_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_280_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_281_) );
OAI21X1 OAI21X1_106 ( .A(_280_), .B(_281_), .C(_24__3_), .Y(_282_) );
NAND2X1 NAND2X1_106 ( .A(_282_), .B(_286_), .Y(_22__3_) );
OAI21X1 OAI21X1_107 ( .A(_283_), .B(_280_), .C(_285_), .Y(_20_) );
INVX1 INVX1_68 ( .A(_24__1_), .Y(_290_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_291_) );
NAND2X1 NAND2X1_107 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_292_) );
NAND3X1 NAND3X1_39 ( .A(_290_), .B(_292_), .C(_291_), .Y(_293_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_287_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_288_) );
OAI21X1 OAI21X1_108 ( .A(_287_), .B(_288_), .C(_24__1_), .Y(_289_) );
NAND2X1 NAND2X1_108 ( .A(_289_), .B(_293_), .Y(_22__1_) );
OAI21X1 OAI21X1_109 ( .A(_290_), .B(_287_), .C(_292_), .Y(_24__2_) );
INVX1 INVX1_69 ( .A(_24__2_), .Y(_297_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_298_) );
NAND2X1 NAND2X1_109 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_299_) );
NAND3X1 NAND3X1_40 ( .A(_297_), .B(_299_), .C(_298_), .Y(_300_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_294_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_295_) );
OAI21X1 OAI21X1_110 ( .A(_294_), .B(_295_), .C(_24__2_), .Y(_296_) );
NAND2X1 NAND2X1_110 ( .A(_296_), .B(_300_), .Y(_22__2_) );
OAI21X1 OAI21X1_111 ( .A(_297_), .B(_294_), .C(_299_), .Y(_24__3_) );
INVX1 INVX1_70 ( .A(_25_), .Y(_301_) );
NAND2X1 NAND2X1_111 ( .A(_26_), .B(w_cout_4_), .Y(_302_) );
OAI21X1 OAI21X1_112 ( .A(w_cout_4_), .B(_301_), .C(_302_), .Y(w_cout_5_) );
INVX1 INVX1_71 ( .A(_27__0_), .Y(_303_) );
NAND2X1 NAND2X1_112 ( .A(_28__0_), .B(w_cout_4_), .Y(_304_) );
OAI21X1 OAI21X1_113 ( .A(w_cout_4_), .B(_303_), .C(_304_), .Y(_0__20_) );
INVX1 INVX1_72 ( .A(_27__1_), .Y(_305_) );
NAND2X1 NAND2X1_113 ( .A(w_cout_4_), .B(_28__1_), .Y(_306_) );
OAI21X1 OAI21X1_114 ( .A(w_cout_4_), .B(_305_), .C(_306_), .Y(_0__21_) );
INVX1 INVX1_73 ( .A(_27__2_), .Y(_307_) );
NAND2X1 NAND2X1_114 ( .A(w_cout_4_), .B(_28__2_), .Y(_308_) );
OAI21X1 OAI21X1_115 ( .A(w_cout_4_), .B(_307_), .C(_308_), .Y(_0__22_) );
INVX1 INVX1_74 ( .A(_27__3_), .Y(_309_) );
NAND2X1 NAND2X1_115 ( .A(w_cout_4_), .B(_28__3_), .Y(_310_) );
OAI21X1 OAI21X1_116 ( .A(w_cout_4_), .B(_309_), .C(_310_), .Y(_0__23_) );
INVX1 INVX1_75 ( .A(gnd), .Y(_314_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_315_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_316_) );
NAND3X1 NAND3X1_41 ( .A(_314_), .B(_316_), .C(_315_), .Y(_317_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_311_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_312_) );
OAI21X1 OAI21X1_117 ( .A(_311_), .B(_312_), .C(gnd), .Y(_313_) );
NAND2X1 NAND2X1_117 ( .A(_313_), .B(_317_), .Y(_27__0_) );
OAI21X1 OAI21X1_118 ( .A(_314_), .B(_311_), .C(_316_), .Y(_29__1_) );
INVX1 INVX1_76 ( .A(_29__3_), .Y(_321_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_322_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_323_) );
NAND3X1 NAND3X1_42 ( .A(_321_), .B(_323_), .C(_322_), .Y(_324_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_318_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_319_) );
OAI21X1 OAI21X1_119 ( .A(_318_), .B(_319_), .C(_29__3_), .Y(_320_) );
NAND2X1 NAND2X1_119 ( .A(_320_), .B(_324_), .Y(_27__3_) );
OAI21X1 OAI21X1_120 ( .A(_321_), .B(_318_), .C(_323_), .Y(_25_) );
INVX1 INVX1_77 ( .A(_29__1_), .Y(_328_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_329_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_330_) );
NAND3X1 NAND3X1_43 ( .A(_328_), .B(_330_), .C(_329_), .Y(_331_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_325_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_326_) );
OAI21X1 OAI21X1_121 ( .A(_325_), .B(_326_), .C(_29__1_), .Y(_327_) );
NAND2X1 NAND2X1_121 ( .A(_327_), .B(_331_), .Y(_27__1_) );
OAI21X1 OAI21X1_122 ( .A(_328_), .B(_325_), .C(_330_), .Y(_29__2_) );
INVX1 INVX1_78 ( .A(_29__2_), .Y(_335_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_336_) );
NAND2X1 NAND2X1_122 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_337_) );
NAND3X1 NAND3X1_44 ( .A(_335_), .B(_337_), .C(_336_), .Y(_338_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_332_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_333_) );
OAI21X1 OAI21X1_123 ( .A(_332_), .B(_333_), .C(_29__2_), .Y(_334_) );
NAND2X1 NAND2X1_123 ( .A(_334_), .B(_338_), .Y(_27__2_) );
OAI21X1 OAI21X1_124 ( .A(_335_), .B(_332_), .C(_337_), .Y(_29__3_) );
INVX1 INVX1_79 ( .A(vdd), .Y(_342_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_343_) );
NAND2X1 NAND2X1_124 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_344_) );
NAND3X1 NAND3X1_45 ( .A(_342_), .B(_344_), .C(_343_), .Y(_345_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_339_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_340_) );
OAI21X1 OAI21X1_125 ( .A(_339_), .B(_340_), .C(vdd), .Y(_341_) );
NAND2X1 NAND2X1_125 ( .A(_341_), .B(_345_), .Y(_28__0_) );
OAI21X1 OAI21X1_126 ( .A(_342_), .B(_339_), .C(_344_), .Y(_30__1_) );
INVX1 INVX1_80 ( .A(_30__3_), .Y(_349_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_350_) );
NAND2X1 NAND2X1_126 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_351_) );
NAND3X1 NAND3X1_46 ( .A(_349_), .B(_351_), .C(_350_), .Y(_352_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_346_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_347_) );
OAI21X1 OAI21X1_127 ( .A(_346_), .B(_347_), .C(_30__3_), .Y(_348_) );
NAND2X1 NAND2X1_127 ( .A(_348_), .B(_352_), .Y(_28__3_) );
OAI21X1 OAI21X1_128 ( .A(_349_), .B(_346_), .C(_351_), .Y(_26_) );
INVX1 INVX1_81 ( .A(_30__1_), .Y(_356_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_357_) );
NAND2X1 NAND2X1_128 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_358_) );
NAND3X1 NAND3X1_47 ( .A(_356_), .B(_358_), .C(_357_), .Y(_359_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_353_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_354_) );
OAI21X1 OAI21X1_129 ( .A(_353_), .B(_354_), .C(_30__1_), .Y(_355_) );
NAND2X1 NAND2X1_129 ( .A(_355_), .B(_359_), .Y(_28__1_) );
OAI21X1 OAI21X1_130 ( .A(_356_), .B(_353_), .C(_358_), .Y(_30__2_) );
INVX1 INVX1_82 ( .A(_30__2_), .Y(_363_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_364_) );
NAND2X1 NAND2X1_130 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_365_) );
NAND3X1 NAND3X1_48 ( .A(_363_), .B(_365_), .C(_364_), .Y(_366_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_360_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_361_) );
OAI21X1 OAI21X1_131 ( .A(_360_), .B(_361_), .C(_30__2_), .Y(_362_) );
NAND2X1 NAND2X1_131 ( .A(_362_), .B(_366_), .Y(_28__2_) );
OAI21X1 OAI21X1_132 ( .A(_363_), .B(_360_), .C(_365_), .Y(_30__3_) );
INVX1 INVX1_83 ( .A(_31_), .Y(_367_) );
NAND2X1 NAND2X1_132 ( .A(_32_), .B(w_cout_5_), .Y(_368_) );
OAI21X1 OAI21X1_133 ( .A(w_cout_5_), .B(_367_), .C(_368_), .Y(csa_inst_cin) );
INVX1 INVX1_84 ( .A(_33__0_), .Y(_369_) );
NAND2X1 NAND2X1_133 ( .A(_34__0_), .B(w_cout_5_), .Y(_370_) );
OAI21X1 OAI21X1_134 ( .A(w_cout_5_), .B(_369_), .C(_370_), .Y(_0__24_) );
INVX1 INVX1_85 ( .A(_33__1_), .Y(_371_) );
NAND2X1 NAND2X1_134 ( .A(w_cout_5_), .B(_34__1_), .Y(_372_) );
OAI21X1 OAI21X1_135 ( .A(w_cout_5_), .B(_371_), .C(_372_), .Y(_0__25_) );
INVX1 INVX1_86 ( .A(_33__2_), .Y(_373_) );
NAND2X1 NAND2X1_135 ( .A(w_cout_5_), .B(_34__2_), .Y(_374_) );
OAI21X1 OAI21X1_136 ( .A(w_cout_5_), .B(_373_), .C(_374_), .Y(_0__26_) );
INVX1 INVX1_87 ( .A(_33__3_), .Y(_375_) );
NAND2X1 NAND2X1_136 ( .A(w_cout_5_), .B(_34__3_), .Y(_376_) );
OAI21X1 OAI21X1_137 ( .A(w_cout_5_), .B(_375_), .C(_376_), .Y(_0__27_) );
INVX1 INVX1_88 ( .A(gnd), .Y(_380_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_381_) );
NAND2X1 NAND2X1_137 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_382_) );
NAND3X1 NAND3X1_49 ( .A(_380_), .B(_382_), .C(_381_), .Y(_383_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_377_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_378_) );
OAI21X1 OAI21X1_138 ( .A(_377_), .B(_378_), .C(gnd), .Y(_379_) );
NAND2X1 NAND2X1_138 ( .A(_379_), .B(_383_), .Y(_33__0_) );
OAI21X1 OAI21X1_139 ( .A(_380_), .B(_377_), .C(_382_), .Y(_35__1_) );
INVX1 INVX1_89 ( .A(_35__3_), .Y(_387_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_388_) );
NAND2X1 NAND2X1_139 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_389_) );
NAND3X1 NAND3X1_50 ( .A(_387_), .B(_389_), .C(_388_), .Y(_390_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_384_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_385_) );
OAI21X1 OAI21X1_140 ( .A(_384_), .B(_385_), .C(_35__3_), .Y(_386_) );
NAND2X1 NAND2X1_140 ( .A(_386_), .B(_390_), .Y(_33__3_) );
OAI21X1 OAI21X1_141 ( .A(_387_), .B(_384_), .C(_389_), .Y(_31_) );
INVX1 INVX1_90 ( .A(_35__1_), .Y(_394_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_395_) );
NAND2X1 NAND2X1_141 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_396_) );
NAND3X1 NAND3X1_51 ( .A(_394_), .B(_396_), .C(_395_), .Y(_397_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_391_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_392_) );
OAI21X1 OAI21X1_142 ( .A(_391_), .B(_392_), .C(_35__1_), .Y(_393_) );
NAND2X1 NAND2X1_142 ( .A(_393_), .B(_397_), .Y(_33__1_) );
OAI21X1 OAI21X1_143 ( .A(_394_), .B(_391_), .C(_396_), .Y(_35__2_) );
INVX1 INVX1_91 ( .A(_35__2_), .Y(_401_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_402_) );
NAND2X1 NAND2X1_143 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_403_) );
NAND3X1 NAND3X1_52 ( .A(_401_), .B(_403_), .C(_402_), .Y(_404_) );
BUFX2 BUFX2_33 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_34 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_35 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_36 ( .A(rca_inst_fa31_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_37 ( .A(gnd), .Y(_0__28_) );
BUFX2 BUFX2_38 ( .A(gnd), .Y(_0__29_) );
BUFX2 BUFX2_39 ( .A(gnd), .Y(_0__30_) );
BUFX2 BUFX2_40 ( .A(rca_inst_cout), .Y(w_cout_0_) );
BUFX2 BUFX2_41 ( .A(csa_inst_cin), .Y(w_cout_6_) );
endmodule
