module csa_22bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_5_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_31_) );
NAND2X1 NAND2X1_1 ( .A(_2_), .B(1'b0), .Y(_32_) );
OAI21X1 OAI21X1_1 ( .A(1'b0), .B(_31_), .C(_32_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3__2_), .Y(_33_) );
NAND2X1 NAND2X1_2 ( .A(_4__2_), .B(1'b0), .Y(_34_) );
OAI21X1 OAI21X1_2 ( .A(1'b0), .B(_33_), .C(_34_), .Y(_0__4_) );
INVX1 INVX1_3 ( .A(_3__3_), .Y(_35_) );
NAND2X1 NAND2X1_3 ( .A(1'b0), .B(_4__3_), .Y(_36_) );
OAI21X1 OAI21X1_3 ( .A(1'b0), .B(_35_), .C(_36_), .Y(_0__5_) );
INVX1 INVX1_4 ( .A(_3__0_), .Y(_37_) );
NAND2X1 NAND2X1_4 ( .A(1'b0), .B(_4__0_), .Y(_38_) );
OAI21X1 OAI21X1_4 ( .A(1'b0), .B(_37_), .C(_38_), .Y(_0__2_) );
INVX1 INVX1_5 ( .A(_3__1_), .Y(_39_) );
NAND2X1 NAND2X1_5 ( .A(1'b0), .B(_4__1_), .Y(_40_) );
OAI21X1 OAI21X1_5 ( .A(1'b0), .B(_39_), .C(_40_), .Y(_0__3_) );
INVX1 INVX1_6 ( .A(_7_), .Y(_41_) );
NAND2X1 NAND2X1_6 ( .A(_8_), .B(w_cout_1_), .Y(_42_) );
OAI21X1 OAI21X1_6 ( .A(w_cout_1_), .B(_41_), .C(_42_), .Y(w_cout_2_) );
INVX1 INVX1_7 ( .A(_9__2_), .Y(_43_) );
NAND2X1 NAND2X1_7 ( .A(_10__2_), .B(w_cout_1_), .Y(_44_) );
OAI21X1 OAI21X1_7 ( .A(w_cout_1_), .B(_43_), .C(_44_), .Y(_0__8_) );
INVX1 INVX1_8 ( .A(_9__3_), .Y(_45_) );
NAND2X1 NAND2X1_8 ( .A(w_cout_1_), .B(_10__3_), .Y(_46_) );
OAI21X1 OAI21X1_8 ( .A(w_cout_1_), .B(_45_), .C(_46_), .Y(_0__9_) );
INVX1 INVX1_9 ( .A(_9__0_), .Y(_47_) );
NAND2X1 NAND2X1_9 ( .A(w_cout_1_), .B(_10__0_), .Y(_48_) );
OAI21X1 OAI21X1_9 ( .A(w_cout_1_), .B(_47_), .C(_48_), .Y(_0__6_) );
INVX1 INVX1_10 ( .A(_9__1_), .Y(_49_) );
NAND2X1 NAND2X1_10 ( .A(w_cout_1_), .B(_10__1_), .Y(_50_) );
OAI21X1 OAI21X1_10 ( .A(w_cout_1_), .B(_49_), .C(_50_), .Y(_0__7_) );
INVX1 INVX1_11 ( .A(_13_), .Y(_51_) );
NAND2X1 NAND2X1_11 ( .A(_14_), .B(w_cout_2_), .Y(_52_) );
OAI21X1 OAI21X1_11 ( .A(w_cout_2_), .B(_51_), .C(_52_), .Y(w_cout_3_) );
INVX1 INVX1_12 ( .A(_15__2_), .Y(_53_) );
NAND2X1 NAND2X1_12 ( .A(_16__2_), .B(w_cout_2_), .Y(_54_) );
OAI21X1 OAI21X1_12 ( .A(w_cout_2_), .B(_53_), .C(_54_), .Y(_0__12_) );
INVX1 INVX1_13 ( .A(_15__3_), .Y(_55_) );
NAND2X1 NAND2X1_13 ( .A(w_cout_2_), .B(_16__3_), .Y(_56_) );
OAI21X1 OAI21X1_13 ( .A(w_cout_2_), .B(_55_), .C(_56_), .Y(_0__13_) );
INVX1 INVX1_14 ( .A(_15__0_), .Y(_57_) );
NAND2X1 NAND2X1_14 ( .A(w_cout_2_), .B(_16__0_), .Y(_58_) );
OAI21X1 OAI21X1_14 ( .A(w_cout_2_), .B(_57_), .C(_58_), .Y(_0__10_) );
INVX1 INVX1_15 ( .A(_15__1_), .Y(_59_) );
NAND2X1 NAND2X1_15 ( .A(w_cout_2_), .B(_16__1_), .Y(_60_) );
OAI21X1 OAI21X1_15 ( .A(w_cout_2_), .B(_59_), .C(_60_), .Y(_0__11_) );
INVX1 INVX1_16 ( .A(_19_), .Y(_61_) );
NAND2X1 NAND2X1_16 ( .A(_20_), .B(w_cout_3_), .Y(_62_) );
OAI21X1 OAI21X1_16 ( .A(w_cout_3_), .B(_61_), .C(_62_), .Y(w_cout_4_) );
INVX1 INVX1_17 ( .A(_21__2_), .Y(_63_) );
NAND2X1 NAND2X1_17 ( .A(_22__2_), .B(w_cout_3_), .Y(_64_) );
OAI21X1 OAI21X1_17 ( .A(w_cout_3_), .B(_63_), .C(_64_), .Y(_0__16_) );
INVX1 INVX1_18 ( .A(_21__3_), .Y(_65_) );
NAND2X1 NAND2X1_18 ( .A(w_cout_3_), .B(_22__3_), .Y(_66_) );
OAI21X1 OAI21X1_18 ( .A(w_cout_3_), .B(_65_), .C(_66_), .Y(_0__17_) );
INVX1 INVX1_19 ( .A(_21__0_), .Y(_67_) );
NAND2X1 NAND2X1_19 ( .A(w_cout_3_), .B(_22__0_), .Y(_68_) );
OAI21X1 OAI21X1_19 ( .A(w_cout_3_), .B(_67_), .C(_68_), .Y(_0__14_) );
INVX1 INVX1_20 ( .A(_21__1_), .Y(_69_) );
NAND2X1 NAND2X1_20 ( .A(w_cout_3_), .B(_22__1_), .Y(_70_) );
OAI21X1 OAI21X1_20 ( .A(w_cout_3_), .B(_69_), .C(_70_), .Y(_0__15_) );
INVX1 INVX1_21 ( .A(_25_), .Y(_71_) );
NAND2X1 NAND2X1_21 ( .A(_26_), .B(w_cout_4_), .Y(_72_) );
OAI21X1 OAI21X1_21 ( .A(w_cout_4_), .B(_71_), .C(_72_), .Y(w_cout_5_) );
INVX1 INVX1_22 ( .A(_27__2_), .Y(_73_) );
NAND2X1 NAND2X1_22 ( .A(_28__2_), .B(w_cout_4_), .Y(_74_) );
OAI21X1 OAI21X1_22 ( .A(w_cout_4_), .B(_73_), .C(_74_), .Y(_0__20_) );
INVX1 INVX1_23 ( .A(_27__3_), .Y(_75_) );
NAND2X1 NAND2X1_23 ( .A(w_cout_4_), .B(_28__3_), .Y(_76_) );
OAI21X1 OAI21X1_23 ( .A(w_cout_4_), .B(_75_), .C(_76_), .Y(_0__21_) );
INVX1 INVX1_24 ( .A(_27__0_), .Y(_77_) );
NAND2X1 NAND2X1_24 ( .A(w_cout_4_), .B(_28__0_), .Y(_78_) );
OAI21X1 OAI21X1_24 ( .A(w_cout_4_), .B(_77_), .C(_78_), .Y(_0__18_) );
INVX1 INVX1_25 ( .A(_27__1_), .Y(_79_) );
NAND2X1 NAND2X1_25 ( .A(w_cout_4_), .B(_28__1_), .Y(_80_) );
OAI21X1 OAI21X1_25 ( .A(w_cout_4_), .B(_79_), .C(_80_), .Y(_0__19_) );
INVX1 INVX1_26 ( .A(1'b0), .Y(_84_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_85_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_86_) );
NAND3X1 NAND3X1_1 ( .A(_84_), .B(_86_), .C(_85_), .Y(_87_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_81_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_82_) );
OAI21X1 OAI21X1_26 ( .A(_81_), .B(_82_), .C(1'b0), .Y(_83_) );
NAND2X1 NAND2X1_27 ( .A(_83_), .B(_87_), .Y(_3__0_) );
OAI21X1 OAI21X1_27 ( .A(_84_), .B(_81_), .C(_86_), .Y(_5__1_) );
INVX1 INVX1_27 ( .A(_5__1_), .Y(_91_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_92_) );
NAND2X1 NAND2X1_28 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_93_) );
NAND3X1 NAND3X1_2 ( .A(_91_), .B(_93_), .C(_92_), .Y(_94_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_88_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_89_) );
OAI21X1 OAI21X1_28 ( .A(_88_), .B(_89_), .C(_5__1_), .Y(_90_) );
NAND2X1 NAND2X1_29 ( .A(_90_), .B(_94_), .Y(_3__1_) );
OAI21X1 OAI21X1_29 ( .A(_91_), .B(_88_), .C(_93_), .Y(_5__2_) );
INVX1 INVX1_28 ( .A(_5__2_), .Y(_98_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_99_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_100_) );
NAND3X1 NAND3X1_3 ( .A(_98_), .B(_100_), .C(_99_), .Y(_101_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_95_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_96_) );
OAI21X1 OAI21X1_30 ( .A(_95_), .B(_96_), .C(_5__2_), .Y(_97_) );
NAND2X1 NAND2X1_31 ( .A(_97_), .B(_101_), .Y(_3__2_) );
OAI21X1 OAI21X1_31 ( .A(_98_), .B(_95_), .C(_100_), .Y(_5__3_) );
INVX1 INVX1_29 ( .A(_5__3_), .Y(_105_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_106_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_107_) );
NAND3X1 NAND3X1_4 ( .A(_105_), .B(_107_), .C(_106_), .Y(_108_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_102_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_103_) );
OAI21X1 OAI21X1_32 ( .A(_102_), .B(_103_), .C(_5__3_), .Y(_104_) );
NAND2X1 NAND2X1_33 ( .A(_104_), .B(_108_), .Y(_3__3_) );
OAI21X1 OAI21X1_33 ( .A(_105_), .B(_102_), .C(_107_), .Y(_1_) );
INVX1 INVX1_30 ( .A(1'b1), .Y(_112_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_113_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_114_) );
NAND3X1 NAND3X1_5 ( .A(_112_), .B(_114_), .C(_113_), .Y(_115_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_109_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_110_) );
OAI21X1 OAI21X1_34 ( .A(_109_), .B(_110_), .C(1'b1), .Y(_111_) );
NAND2X1 NAND2X1_35 ( .A(_111_), .B(_115_), .Y(_4__0_) );
OAI21X1 OAI21X1_35 ( .A(_112_), .B(_109_), .C(_114_), .Y(_6__1_) );
INVX1 INVX1_31 ( .A(_6__1_), .Y(_119_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_120_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_121_) );
NAND3X1 NAND3X1_6 ( .A(_119_), .B(_121_), .C(_120_), .Y(_122_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_116_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_117_) );
OAI21X1 OAI21X1_36 ( .A(_116_), .B(_117_), .C(_6__1_), .Y(_118_) );
NAND2X1 NAND2X1_37 ( .A(_118_), .B(_122_), .Y(_4__1_) );
OAI21X1 OAI21X1_37 ( .A(_119_), .B(_116_), .C(_121_), .Y(_6__2_) );
INVX1 INVX1_32 ( .A(_6__2_), .Y(_126_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_127_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_128_) );
NAND3X1 NAND3X1_7 ( .A(_126_), .B(_128_), .C(_127_), .Y(_129_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_123_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_124_) );
OAI21X1 OAI21X1_38 ( .A(_123_), .B(_124_), .C(_6__2_), .Y(_125_) );
NAND2X1 NAND2X1_39 ( .A(_125_), .B(_129_), .Y(_4__2_) );
OAI21X1 OAI21X1_39 ( .A(_126_), .B(_123_), .C(_128_), .Y(_6__3_) );
INVX1 INVX1_33 ( .A(_6__3_), .Y(_133_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_134_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_135_) );
NAND3X1 NAND3X1_8 ( .A(_133_), .B(_135_), .C(_134_), .Y(_136_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_130_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_131_) );
OAI21X1 OAI21X1_40 ( .A(_130_), .B(_131_), .C(_6__3_), .Y(_132_) );
NAND2X1 NAND2X1_41 ( .A(_132_), .B(_136_), .Y(_4__3_) );
OAI21X1 OAI21X1_41 ( .A(_133_), .B(_130_), .C(_135_), .Y(_2_) );
INVX1 INVX1_34 ( .A(1'b0), .Y(_140_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_141_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_142_) );
NAND3X1 NAND3X1_9 ( .A(_140_), .B(_142_), .C(_141_), .Y(_143_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_137_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_138_) );
OAI21X1 OAI21X1_42 ( .A(_137_), .B(_138_), .C(1'b0), .Y(_139_) );
NAND2X1 NAND2X1_43 ( .A(_139_), .B(_143_), .Y(_9__0_) );
OAI21X1 OAI21X1_43 ( .A(_140_), .B(_137_), .C(_142_), .Y(_11__1_) );
INVX1 INVX1_35 ( .A(_11__1_), .Y(_147_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_148_) );
NAND2X1 NAND2X1_44 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_149_) );
NAND3X1 NAND3X1_10 ( .A(_147_), .B(_149_), .C(_148_), .Y(_150_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_144_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_145_) );
OAI21X1 OAI21X1_44 ( .A(_144_), .B(_145_), .C(_11__1_), .Y(_146_) );
NAND2X1 NAND2X1_45 ( .A(_146_), .B(_150_), .Y(_9__1_) );
OAI21X1 OAI21X1_45 ( .A(_147_), .B(_144_), .C(_149_), .Y(_11__2_) );
INVX1 INVX1_36 ( .A(_11__2_), .Y(_154_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_155_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_156_) );
NAND3X1 NAND3X1_11 ( .A(_154_), .B(_156_), .C(_155_), .Y(_157_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_151_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_152_) );
OAI21X1 OAI21X1_46 ( .A(_151_), .B(_152_), .C(_11__2_), .Y(_153_) );
NAND2X1 NAND2X1_47 ( .A(_153_), .B(_157_), .Y(_9__2_) );
OAI21X1 OAI21X1_47 ( .A(_154_), .B(_151_), .C(_156_), .Y(_11__3_) );
INVX1 INVX1_37 ( .A(_11__3_), .Y(_161_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_162_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_163_) );
NAND3X1 NAND3X1_12 ( .A(_161_), .B(_163_), .C(_162_), .Y(_164_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_158_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_159_) );
OAI21X1 OAI21X1_48 ( .A(_158_), .B(_159_), .C(_11__3_), .Y(_160_) );
NAND2X1 NAND2X1_49 ( .A(_160_), .B(_164_), .Y(_9__3_) );
OAI21X1 OAI21X1_49 ( .A(_161_), .B(_158_), .C(_163_), .Y(_7_) );
INVX1 INVX1_38 ( .A(1'b1), .Y(_168_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_169_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_170_) );
NAND3X1 NAND3X1_13 ( .A(_168_), .B(_170_), .C(_169_), .Y(_171_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_165_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_166_) );
OAI21X1 OAI21X1_50 ( .A(_165_), .B(_166_), .C(1'b1), .Y(_167_) );
NAND2X1 NAND2X1_51 ( .A(_167_), .B(_171_), .Y(_10__0_) );
OAI21X1 OAI21X1_51 ( .A(_168_), .B(_165_), .C(_170_), .Y(_12__1_) );
INVX1 INVX1_39 ( .A(_12__1_), .Y(_175_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_176_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_177_) );
NAND3X1 NAND3X1_14 ( .A(_175_), .B(_177_), .C(_176_), .Y(_178_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_172_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_173_) );
OAI21X1 OAI21X1_52 ( .A(_172_), .B(_173_), .C(_12__1_), .Y(_174_) );
NAND2X1 NAND2X1_53 ( .A(_174_), .B(_178_), .Y(_10__1_) );
OAI21X1 OAI21X1_53 ( .A(_175_), .B(_172_), .C(_177_), .Y(_12__2_) );
INVX1 INVX1_40 ( .A(_12__2_), .Y(_182_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_183_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_184_) );
NAND3X1 NAND3X1_15 ( .A(_182_), .B(_184_), .C(_183_), .Y(_185_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_179_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_180_) );
OAI21X1 OAI21X1_54 ( .A(_179_), .B(_180_), .C(_12__2_), .Y(_181_) );
NAND2X1 NAND2X1_55 ( .A(_181_), .B(_185_), .Y(_10__2_) );
OAI21X1 OAI21X1_55 ( .A(_182_), .B(_179_), .C(_184_), .Y(_12__3_) );
INVX1 INVX1_41 ( .A(_12__3_), .Y(_189_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_190_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_191_) );
NAND3X1 NAND3X1_16 ( .A(_189_), .B(_191_), .C(_190_), .Y(_192_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_186_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_187_) );
OAI21X1 OAI21X1_56 ( .A(_186_), .B(_187_), .C(_12__3_), .Y(_188_) );
NAND2X1 NAND2X1_57 ( .A(_188_), .B(_192_), .Y(_10__3_) );
OAI21X1 OAI21X1_57 ( .A(_189_), .B(_186_), .C(_191_), .Y(_8_) );
INVX1 INVX1_42 ( .A(1'b0), .Y(_196_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_197_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_198_) );
NAND3X1 NAND3X1_17 ( .A(_196_), .B(_198_), .C(_197_), .Y(_199_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_193_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_194_) );
OAI21X1 OAI21X1_58 ( .A(_193_), .B(_194_), .C(1'b0), .Y(_195_) );
NAND2X1 NAND2X1_59 ( .A(_195_), .B(_199_), .Y(_15__0_) );
OAI21X1 OAI21X1_59 ( .A(_196_), .B(_193_), .C(_198_), .Y(_17__1_) );
INVX1 INVX1_43 ( .A(_17__1_), .Y(_203_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_204_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_205_) );
NAND3X1 NAND3X1_18 ( .A(_203_), .B(_205_), .C(_204_), .Y(_206_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_200_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_201_) );
OAI21X1 OAI21X1_60 ( .A(_200_), .B(_201_), .C(_17__1_), .Y(_202_) );
NAND2X1 NAND2X1_61 ( .A(_202_), .B(_206_), .Y(_15__1_) );
OAI21X1 OAI21X1_61 ( .A(_203_), .B(_200_), .C(_205_), .Y(_17__2_) );
INVX1 INVX1_44 ( .A(_17__2_), .Y(_210_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_211_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_212_) );
NAND3X1 NAND3X1_19 ( .A(_210_), .B(_212_), .C(_211_), .Y(_213_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_207_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_208_) );
OAI21X1 OAI21X1_62 ( .A(_207_), .B(_208_), .C(_17__2_), .Y(_209_) );
NAND2X1 NAND2X1_63 ( .A(_209_), .B(_213_), .Y(_15__2_) );
OAI21X1 OAI21X1_63 ( .A(_210_), .B(_207_), .C(_212_), .Y(_17__3_) );
INVX1 INVX1_45 ( .A(_17__3_), .Y(_217_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_218_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_219_) );
NAND3X1 NAND3X1_20 ( .A(_217_), .B(_219_), .C(_218_), .Y(_220_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_214_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_215_) );
OAI21X1 OAI21X1_64 ( .A(_214_), .B(_215_), .C(_17__3_), .Y(_216_) );
NAND2X1 NAND2X1_65 ( .A(_216_), .B(_220_), .Y(_15__3_) );
OAI21X1 OAI21X1_65 ( .A(_217_), .B(_214_), .C(_219_), .Y(_13_) );
INVX1 INVX1_46 ( .A(1'b1), .Y(_224_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_225_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_226_) );
NAND3X1 NAND3X1_21 ( .A(_224_), .B(_226_), .C(_225_), .Y(_227_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_221_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_222_) );
OAI21X1 OAI21X1_66 ( .A(_221_), .B(_222_), .C(1'b1), .Y(_223_) );
NAND2X1 NAND2X1_67 ( .A(_223_), .B(_227_), .Y(_16__0_) );
OAI21X1 OAI21X1_67 ( .A(_224_), .B(_221_), .C(_226_), .Y(_18__1_) );
INVX1 INVX1_47 ( .A(_18__1_), .Y(_231_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_232_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_233_) );
NAND3X1 NAND3X1_22 ( .A(_231_), .B(_233_), .C(_232_), .Y(_234_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_228_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_229_) );
OAI21X1 OAI21X1_68 ( .A(_228_), .B(_229_), .C(_18__1_), .Y(_230_) );
NAND2X1 NAND2X1_69 ( .A(_230_), .B(_234_), .Y(_16__1_) );
OAI21X1 OAI21X1_69 ( .A(_231_), .B(_228_), .C(_233_), .Y(_18__2_) );
INVX1 INVX1_48 ( .A(_18__2_), .Y(_238_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_239_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_240_) );
NAND3X1 NAND3X1_23 ( .A(_238_), .B(_240_), .C(_239_), .Y(_241_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_235_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_236_) );
OAI21X1 OAI21X1_70 ( .A(_235_), .B(_236_), .C(_18__2_), .Y(_237_) );
NAND2X1 NAND2X1_71 ( .A(_237_), .B(_241_), .Y(_16__2_) );
OAI21X1 OAI21X1_71 ( .A(_238_), .B(_235_), .C(_240_), .Y(_18__3_) );
INVX1 INVX1_49 ( .A(_18__3_), .Y(_245_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_246_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_247_) );
NAND3X1 NAND3X1_24 ( .A(_245_), .B(_247_), .C(_246_), .Y(_248_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_242_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_243_) );
OAI21X1 OAI21X1_72 ( .A(_242_), .B(_243_), .C(_18__3_), .Y(_244_) );
NAND2X1 NAND2X1_73 ( .A(_244_), .B(_248_), .Y(_16__3_) );
OAI21X1 OAI21X1_73 ( .A(_245_), .B(_242_), .C(_247_), .Y(_14_) );
INVX1 INVX1_50 ( .A(1'b0), .Y(_252_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_253_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_254_) );
NAND3X1 NAND3X1_25 ( .A(_252_), .B(_254_), .C(_253_), .Y(_255_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_249_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_250_) );
OAI21X1 OAI21X1_74 ( .A(_249_), .B(_250_), .C(1'b0), .Y(_251_) );
NAND2X1 NAND2X1_75 ( .A(_251_), .B(_255_), .Y(_21__0_) );
OAI21X1 OAI21X1_75 ( .A(_252_), .B(_249_), .C(_254_), .Y(_23__1_) );
INVX1 INVX1_51 ( .A(_23__1_), .Y(_259_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_260_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_261_) );
NAND3X1 NAND3X1_26 ( .A(_259_), .B(_261_), .C(_260_), .Y(_262_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_256_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_257_) );
OAI21X1 OAI21X1_76 ( .A(_256_), .B(_257_), .C(_23__1_), .Y(_258_) );
NAND2X1 NAND2X1_77 ( .A(_258_), .B(_262_), .Y(_21__1_) );
OAI21X1 OAI21X1_77 ( .A(_259_), .B(_256_), .C(_261_), .Y(_23__2_) );
INVX1 INVX1_52 ( .A(_23__2_), .Y(_266_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_267_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_268_) );
NAND3X1 NAND3X1_27 ( .A(_266_), .B(_268_), .C(_267_), .Y(_269_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_263_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_264_) );
OAI21X1 OAI21X1_78 ( .A(_263_), .B(_264_), .C(_23__2_), .Y(_265_) );
NAND2X1 NAND2X1_79 ( .A(_265_), .B(_269_), .Y(_21__2_) );
OAI21X1 OAI21X1_79 ( .A(_266_), .B(_263_), .C(_268_), .Y(_23__3_) );
INVX1 INVX1_53 ( .A(_23__3_), .Y(_273_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_274_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_275_) );
NAND3X1 NAND3X1_28 ( .A(_273_), .B(_275_), .C(_274_), .Y(_276_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_270_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_271_) );
OAI21X1 OAI21X1_80 ( .A(_270_), .B(_271_), .C(_23__3_), .Y(_272_) );
NAND2X1 NAND2X1_81 ( .A(_272_), .B(_276_), .Y(_21__3_) );
OAI21X1 OAI21X1_81 ( .A(_273_), .B(_270_), .C(_275_), .Y(_19_) );
INVX1 INVX1_54 ( .A(1'b1), .Y(_280_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_281_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_282_) );
NAND3X1 NAND3X1_29 ( .A(_280_), .B(_282_), .C(_281_), .Y(_283_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_277_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_278_) );
OAI21X1 OAI21X1_82 ( .A(_277_), .B(_278_), .C(1'b1), .Y(_279_) );
NAND2X1 NAND2X1_83 ( .A(_279_), .B(_283_), .Y(_22__0_) );
OAI21X1 OAI21X1_83 ( .A(_280_), .B(_277_), .C(_282_), .Y(_24__1_) );
INVX1 INVX1_55 ( .A(_24__1_), .Y(_287_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_288_) );
NAND2X1 NAND2X1_84 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_289_) );
NAND3X1 NAND3X1_30 ( .A(_287_), .B(_289_), .C(_288_), .Y(_290_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_284_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_285_) );
OAI21X1 OAI21X1_84 ( .A(_284_), .B(_285_), .C(_24__1_), .Y(_286_) );
NAND2X1 NAND2X1_85 ( .A(_286_), .B(_290_), .Y(_22__1_) );
OAI21X1 OAI21X1_85 ( .A(_287_), .B(_284_), .C(_289_), .Y(_24__2_) );
INVX1 INVX1_56 ( .A(_24__2_), .Y(_294_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_295_) );
NAND2X1 NAND2X1_86 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_296_) );
NAND3X1 NAND3X1_31 ( .A(_294_), .B(_296_), .C(_295_), .Y(_297_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_291_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_292_) );
OAI21X1 OAI21X1_86 ( .A(_291_), .B(_292_), .C(_24__2_), .Y(_293_) );
NAND2X1 NAND2X1_87 ( .A(_293_), .B(_297_), .Y(_22__2_) );
OAI21X1 OAI21X1_87 ( .A(_294_), .B(_291_), .C(_296_), .Y(_24__3_) );
INVX1 INVX1_57 ( .A(_24__3_), .Y(_301_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_302_) );
NAND2X1 NAND2X1_88 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_303_) );
NAND3X1 NAND3X1_32 ( .A(_301_), .B(_303_), .C(_302_), .Y(_304_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_298_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_299_) );
OAI21X1 OAI21X1_88 ( .A(_298_), .B(_299_), .C(_24__3_), .Y(_300_) );
NAND2X1 NAND2X1_89 ( .A(_300_), .B(_304_), .Y(_22__3_) );
OAI21X1 OAI21X1_89 ( .A(_301_), .B(_298_), .C(_303_), .Y(_20_) );
INVX1 INVX1_58 ( .A(1'b0), .Y(_308_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_309_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_310_) );
NAND3X1 NAND3X1_33 ( .A(_308_), .B(_310_), .C(_309_), .Y(_311_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_305_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_306_) );
OAI21X1 OAI21X1_90 ( .A(_305_), .B(_306_), .C(1'b0), .Y(_307_) );
NAND2X1 NAND2X1_91 ( .A(_307_), .B(_311_), .Y(_27__0_) );
OAI21X1 OAI21X1_91 ( .A(_308_), .B(_305_), .C(_310_), .Y(_29__1_) );
INVX1 INVX1_59 ( .A(_29__1_), .Y(_315_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_316_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_317_) );
NAND3X1 NAND3X1_34 ( .A(_315_), .B(_317_), .C(_316_), .Y(_318_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_312_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_313_) );
OAI21X1 OAI21X1_92 ( .A(_312_), .B(_313_), .C(_29__1_), .Y(_314_) );
NAND2X1 NAND2X1_93 ( .A(_314_), .B(_318_), .Y(_27__1_) );
OAI21X1 OAI21X1_93 ( .A(_315_), .B(_312_), .C(_317_), .Y(_29__2_) );
INVX1 INVX1_60 ( .A(_29__2_), .Y(_322_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_323_) );
NAND2X1 NAND2X1_94 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_324_) );
NAND3X1 NAND3X1_35 ( .A(_322_), .B(_324_), .C(_323_), .Y(_325_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_319_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_320_) );
OAI21X1 OAI21X1_94 ( .A(_319_), .B(_320_), .C(_29__2_), .Y(_321_) );
NAND2X1 NAND2X1_95 ( .A(_321_), .B(_325_), .Y(_27__2_) );
OAI21X1 OAI21X1_95 ( .A(_322_), .B(_319_), .C(_324_), .Y(_29__3_) );
INVX1 INVX1_61 ( .A(_29__3_), .Y(_329_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_330_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_331_) );
NAND3X1 NAND3X1_36 ( .A(_329_), .B(_331_), .C(_330_), .Y(_332_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_326_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_327_) );
OAI21X1 OAI21X1_96 ( .A(_326_), .B(_327_), .C(_29__3_), .Y(_328_) );
NAND2X1 NAND2X1_97 ( .A(_328_), .B(_332_), .Y(_27__3_) );
OAI21X1 OAI21X1_97 ( .A(_329_), .B(_326_), .C(_331_), .Y(_25_) );
INVX1 INVX1_62 ( .A(1'b1), .Y(_336_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_337_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_338_) );
NAND3X1 NAND3X1_37 ( .A(_336_), .B(_338_), .C(_337_), .Y(_339_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_333_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_334_) );
OAI21X1 OAI21X1_98 ( .A(_333_), .B(_334_), .C(1'b1), .Y(_335_) );
NAND2X1 NAND2X1_99 ( .A(_335_), .B(_339_), .Y(_28__0_) );
OAI21X1 OAI21X1_99 ( .A(_336_), .B(_333_), .C(_338_), .Y(_30__1_) );
INVX1 INVX1_63 ( .A(_30__1_), .Y(_343_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_344_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_345_) );
NAND3X1 NAND3X1_38 ( .A(_343_), .B(_345_), .C(_344_), .Y(_346_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_340_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_341_) );
OAI21X1 OAI21X1_100 ( .A(_340_), .B(_341_), .C(_30__1_), .Y(_342_) );
NAND2X1 NAND2X1_101 ( .A(_342_), .B(_346_), .Y(_28__1_) );
OAI21X1 OAI21X1_101 ( .A(_343_), .B(_340_), .C(_345_), .Y(_30__2_) );
INVX1 INVX1_64 ( .A(_30__2_), .Y(_350_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_351_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_352_) );
NAND3X1 NAND3X1_39 ( .A(_350_), .B(_352_), .C(_351_), .Y(_353_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_347_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_348_) );
OAI21X1 OAI21X1_102 ( .A(_347_), .B(_348_), .C(_30__2_), .Y(_349_) );
NAND2X1 NAND2X1_103 ( .A(_349_), .B(_353_), .Y(_28__2_) );
OAI21X1 OAI21X1_103 ( .A(_350_), .B(_347_), .C(_352_), .Y(_30__3_) );
INVX1 INVX1_65 ( .A(_30__3_), .Y(_357_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_358_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_359_) );
NAND3X1 NAND3X1_40 ( .A(_357_), .B(_359_), .C(_358_), .Y(_360_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_354_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_355_) );
OAI21X1 OAI21X1_104 ( .A(_354_), .B(_355_), .C(_30__3_), .Y(_356_) );
NAND2X1 NAND2X1_105 ( .A(_356_), .B(_360_), .Y(_28__3_) );
OAI21X1 OAI21X1_105 ( .A(_357_), .B(_354_), .C(_359_), .Y(_26_) );
INVX1 INVX1_66 ( .A(1'b0), .Y(_364_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_365_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_366_) );
NAND3X1 NAND3X1_41 ( .A(_364_), .B(_366_), .C(_365_), .Y(_367_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_361_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_362_) );
OAI21X1 OAI21X1_106 ( .A(_361_), .B(_362_), .C(1'b0), .Y(_363_) );
NAND2X1 NAND2X1_107 ( .A(_363_), .B(_367_), .Y(_0__0_) );
OAI21X1 OAI21X1_107 ( .A(_364_), .B(_361_), .C(_366_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_67 ( .A(rca_inst_w_CARRY_1_), .Y(_371_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_372_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_373_) );
NAND3X1 NAND3X1_42 ( .A(_371_), .B(_373_), .C(_372_), .Y(_374_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_368_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_369_) );
OAI21X1 OAI21X1_108 ( .A(_368_), .B(_369_), .C(rca_inst_w_CARRY_1_), .Y(_370_) );
NAND2X1 NAND2X1_109 ( .A(_370_), .B(_374_), .Y(_0__1_) );
BUFX2 BUFX2_24 ( .A(1'b0), .Y(_5__0_) );
BUFX2 BUFX2_25 ( .A(_1_), .Y(_5__4_) );
BUFX2 BUFX2_26 ( .A(1'b1), .Y(_6__0_) );
BUFX2 BUFX2_27 ( .A(_2_), .Y(_6__4_) );
BUFX2 BUFX2_28 ( .A(1'b0), .Y(_11__0_) );
BUFX2 BUFX2_29 ( .A(_7_), .Y(_11__4_) );
BUFX2 BUFX2_30 ( .A(1'b1), .Y(_12__0_) );
BUFX2 BUFX2_31 ( .A(_8_), .Y(_12__4_) );
BUFX2 BUFX2_32 ( .A(1'b0), .Y(_17__0_) );
BUFX2 BUFX2_33 ( .A(_13_), .Y(_17__4_) );
BUFX2 BUFX2_34 ( .A(1'b1), .Y(_18__0_) );
BUFX2 BUFX2_35 ( .A(_14_), .Y(_18__4_) );
BUFX2 BUFX2_36 ( .A(1'b0), .Y(_23__0_) );
BUFX2 BUFX2_37 ( .A(_19_), .Y(_23__4_) );
BUFX2 BUFX2_38 ( .A(1'b1), .Y(_24__0_) );
BUFX2 BUFX2_39 ( .A(_20_), .Y(_24__4_) );
BUFX2 BUFX2_40 ( .A(1'b0), .Y(_29__0_) );
BUFX2 BUFX2_41 ( .A(_25_), .Y(_29__4_) );
BUFX2 BUFX2_42 ( .A(1'b1), .Y(_30__0_) );
BUFX2 BUFX2_43 ( .A(_26_), .Y(_30__4_) );
BUFX2 BUFX2_44 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_45 ( .A(1'b0), .Y(w_cout_0_) );
endmodule
