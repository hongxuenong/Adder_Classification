module cla_17bit (i_add1, i_add2, o_result);

input [16:0] i_add1;
input [16:0] i_add2;
output [17:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_38_) );
INVX1 INVX1_1 ( .A(_38_), .Y(w_C_1_) );
NAND2X1 NAND2X1_2 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_39_) );
NAND2X1 NAND2X1_3 ( .A(_38_), .B(_39_), .Y(_40_) );
OAI21X1 OAI21X1_1 ( .A(i_add2[1]), .B(i_add1[1]), .C(_40_), .Y(_41_) );
INVX1 INVX1_2 ( .A(_41_), .Y(w_C_2_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_42_) );
OR2X2 OR2X2_1 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_43_) );
OR2X2 OR2X2_2 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_44_) );
NAND3X1 NAND3X1_1 ( .A(_43_), .B(_44_), .C(_40_), .Y(_45_) );
NAND2X1 NAND2X1_5 ( .A(_42_), .B(_45_), .Y(w_C_3_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_46_) );
NAND3X1 NAND3X1_2 ( .A(_42_), .B(_46_), .C(_45_), .Y(_47_) );
OAI21X1 OAI21X1_2 ( .A(i_add2[3]), .B(i_add1[3]), .C(_47_), .Y(_48_) );
INVX1 INVX1_3 ( .A(_48_), .Y(w_C_4_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_49_) );
OR2X2 OR2X2_3 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_50_) );
OR2X2 OR2X2_4 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_51_) );
NAND3X1 NAND3X1_3 ( .A(_50_), .B(_51_), .C(_47_), .Y(_52_) );
NAND2X1 NAND2X1_8 ( .A(_49_), .B(_52_), .Y(w_C_5_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_53_) );
NAND3X1 NAND3X1_4 ( .A(_49_), .B(_53_), .C(_52_), .Y(_54_) );
OAI21X1 OAI21X1_3 ( .A(i_add2[5]), .B(i_add1[5]), .C(_54_), .Y(_55_) );
INVX1 INVX1_4 ( .A(_55_), .Y(w_C_6_) );
INVX1 INVX1_5 ( .A(i_add2[6]), .Y(_56_) );
INVX1 INVX1_6 ( .A(i_add1[6]), .Y(_57_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_58_) );
INVX1 INVX1_7 ( .A(_58_), .Y(_59_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_60_) );
INVX1 INVX1_8 ( .A(_60_), .Y(_61_) );
NAND3X1 NAND3X1_5 ( .A(_59_), .B(_61_), .C(_54_), .Y(_62_) );
OAI21X1 OAI21X1_4 ( .A(_56_), .B(_57_), .C(_62_), .Y(w_C_7_) );
NOR2X1 NOR2X1_3 ( .A(_56_), .B(_57_), .Y(_63_) );
INVX1 INVX1_9 ( .A(_63_), .Y(_64_) );
AND2X2 AND2X2_1 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_65_) );
INVX1 INVX1_10 ( .A(_65_), .Y(_66_) );
NAND3X1 NAND3X1_6 ( .A(_64_), .B(_66_), .C(_62_), .Y(_67_) );
OAI21X1 OAI21X1_5 ( .A(i_add2[7]), .B(i_add1[7]), .C(_67_), .Y(_68_) );
INVX1 INVX1_11 ( .A(_68_), .Y(w_C_8_) );
INVX1 INVX1_12 ( .A(i_add2[8]), .Y(_69_) );
INVX1 INVX1_13 ( .A(i_add1[8]), .Y(_70_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_71_) );
INVX1 INVX1_14 ( .A(_71_), .Y(_72_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_73_) );
INVX1 INVX1_15 ( .A(_73_), .Y(_74_) );
NAND3X1 NAND3X1_7 ( .A(_72_), .B(_74_), .C(_67_), .Y(_75_) );
OAI21X1 OAI21X1_6 ( .A(_69_), .B(_70_), .C(_75_), .Y(w_C_9_) );
NOR2X1 NOR2X1_6 ( .A(_69_), .B(_70_), .Y(_76_) );
INVX1 INVX1_16 ( .A(_76_), .Y(_0_) );
AND2X2 AND2X2_2 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_1_) );
INVX1 INVX1_17 ( .A(_1_), .Y(_2_) );
NAND3X1 NAND3X1_8 ( .A(_0_), .B(_2_), .C(_75_), .Y(_3_) );
OAI21X1 OAI21X1_7 ( .A(i_add2[9]), .B(i_add1[9]), .C(_3_), .Y(_4_) );
INVX1 INVX1_18 ( .A(_4_), .Y(w_C_10_) );
INVX1 INVX1_19 ( .A(i_add2[10]), .Y(_5_) );
INVX1 INVX1_20 ( .A(i_add1[10]), .Y(_6_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_7_) );
INVX1 INVX1_21 ( .A(_7_), .Y(_8_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_9_) );
INVX1 INVX1_22 ( .A(_9_), .Y(_10_) );
NAND3X1 NAND3X1_9 ( .A(_8_), .B(_10_), .C(_3_), .Y(_11_) );
OAI21X1 OAI21X1_8 ( .A(_5_), .B(_6_), .C(_11_), .Y(w_C_11_) );
NOR2X1 NOR2X1_9 ( .A(_5_), .B(_6_), .Y(_12_) );
INVX1 INVX1_23 ( .A(_12_), .Y(_13_) );
AND2X2 AND2X2_3 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_14_) );
INVX1 INVX1_24 ( .A(_14_), .Y(_15_) );
NAND3X1 NAND3X1_10 ( .A(_13_), .B(_15_), .C(_11_), .Y(_16_) );
OAI21X1 OAI21X1_9 ( .A(i_add2[11]), .B(i_add1[11]), .C(_16_), .Y(_17_) );
INVX1 INVX1_25 ( .A(_17_), .Y(w_C_12_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_18_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_19_) );
OAI21X1 OAI21X1_10 ( .A(_19_), .B(_17_), .C(_18_), .Y(w_C_13_) );
OR2X2 OR2X2_5 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_20_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_21_) );
INVX1 INVX1_26 ( .A(_21_), .Y(_22_) );
INVX1 INVX1_27 ( .A(_19_), .Y(_23_) );
NAND3X1 NAND3X1_11 ( .A(_22_), .B(_23_), .C(_16_), .Y(_24_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_25_) );
NAND3X1 NAND3X1_12 ( .A(_18_), .B(_25_), .C(_24_), .Y(_26_) );
AND2X2 AND2X2_4 ( .A(_26_), .B(_20_), .Y(w_C_14_) );
INVX1 INVX1_28 ( .A(i_add2[14]), .Y(_27_) );
INVX1 INVX1_29 ( .A(i_add1[14]), .Y(_28_) );
NAND2X1 NAND2X1_12 ( .A(_27_), .B(_28_), .Y(_29_) );
NAND3X1 NAND3X1_13 ( .A(_20_), .B(_29_), .C(_26_), .Y(_30_) );
OAI21X1 OAI21X1_11 ( .A(_27_), .B(_28_), .C(_30_), .Y(w_C_15_) );
OR2X2 OR2X2_6 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_31_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_32_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_33_) );
NAND3X1 NAND3X1_14 ( .A(_32_), .B(_33_), .C(_30_), .Y(_34_) );
AND2X2 AND2X2_5 ( .A(_34_), .B(_31_), .Y(w_C_16_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_35_) );
OR2X2 OR2X2_7 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_36_) );
NAND3X1 NAND3X1_15 ( .A(_31_), .B(_36_), .C(_34_), .Y(_37_) );
NAND2X1 NAND2X1_16 ( .A(_35_), .B(_37_), .Y(w_C_17_) );
BUFX2 BUFX2_1 ( .A(_77__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_77__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_77__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_77__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_77__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_77__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_77__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_77__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_77__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_77__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_77__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_77__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_77__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_77__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_77__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_77__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_77__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(w_C_17_), .Y(o_result[17]) );
INVX1 INVX1_30 ( .A(w_C_4_), .Y(_81_) );
OR2X2 OR2X2_8 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_82_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_83_) );
NAND3X1 NAND3X1_16 ( .A(_81_), .B(_83_), .C(_82_), .Y(_84_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_78_) );
AND2X2 AND2X2_6 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_79_) );
OAI21X1 OAI21X1_12 ( .A(_78_), .B(_79_), .C(w_C_4_), .Y(_80_) );
NAND2X1 NAND2X1_18 ( .A(_80_), .B(_84_), .Y(_77__4_) );
INVX1 INVX1_31 ( .A(w_C_5_), .Y(_88_) );
OR2X2 OR2X2_9 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_89_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_90_) );
NAND3X1 NAND3X1_17 ( .A(_88_), .B(_90_), .C(_89_), .Y(_91_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_85_) );
AND2X2 AND2X2_7 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_86_) );
OAI21X1 OAI21X1_13 ( .A(_85_), .B(_86_), .C(w_C_5_), .Y(_87_) );
NAND2X1 NAND2X1_20 ( .A(_87_), .B(_91_), .Y(_77__5_) );
INVX1 INVX1_32 ( .A(w_C_6_), .Y(_95_) );
OR2X2 OR2X2_10 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_96_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_97_) );
NAND3X1 NAND3X1_18 ( .A(_95_), .B(_97_), .C(_96_), .Y(_98_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_92_) );
AND2X2 AND2X2_8 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_93_) );
OAI21X1 OAI21X1_14 ( .A(_92_), .B(_93_), .C(w_C_6_), .Y(_94_) );
NAND2X1 NAND2X1_22 ( .A(_94_), .B(_98_), .Y(_77__6_) );
INVX1 INVX1_33 ( .A(w_C_7_), .Y(_102_) );
OR2X2 OR2X2_11 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_103_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_104_) );
NAND3X1 NAND3X1_19 ( .A(_102_), .B(_104_), .C(_103_), .Y(_105_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_99_) );
AND2X2 AND2X2_9 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_100_) );
OAI21X1 OAI21X1_15 ( .A(_99_), .B(_100_), .C(w_C_7_), .Y(_101_) );
NAND2X1 NAND2X1_24 ( .A(_101_), .B(_105_), .Y(_77__7_) );
INVX1 INVX1_34 ( .A(w_C_8_), .Y(_109_) );
OR2X2 OR2X2_12 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_110_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_111_) );
NAND3X1 NAND3X1_20 ( .A(_109_), .B(_111_), .C(_110_), .Y(_112_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_106_) );
AND2X2 AND2X2_10 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_107_) );
OAI21X1 OAI21X1_16 ( .A(_106_), .B(_107_), .C(w_C_8_), .Y(_108_) );
NAND2X1 NAND2X1_26 ( .A(_108_), .B(_112_), .Y(_77__8_) );
INVX1 INVX1_35 ( .A(w_C_9_), .Y(_116_) );
OR2X2 OR2X2_13 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_117_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_118_) );
NAND3X1 NAND3X1_21 ( .A(_116_), .B(_118_), .C(_117_), .Y(_119_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_113_) );
AND2X2 AND2X2_11 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_114_) );
OAI21X1 OAI21X1_17 ( .A(_113_), .B(_114_), .C(w_C_9_), .Y(_115_) );
NAND2X1 NAND2X1_28 ( .A(_115_), .B(_119_), .Y(_77__9_) );
INVX1 INVX1_36 ( .A(w_C_10_), .Y(_123_) );
OR2X2 OR2X2_14 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_124_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_125_) );
NAND3X1 NAND3X1_22 ( .A(_123_), .B(_125_), .C(_124_), .Y(_126_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_120_) );
AND2X2 AND2X2_12 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_121_) );
OAI21X1 OAI21X1_18 ( .A(_120_), .B(_121_), .C(w_C_10_), .Y(_122_) );
NAND2X1 NAND2X1_30 ( .A(_122_), .B(_126_), .Y(_77__10_) );
INVX1 INVX1_37 ( .A(w_C_11_), .Y(_130_) );
OR2X2 OR2X2_15 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_131_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_132_) );
NAND3X1 NAND3X1_23 ( .A(_130_), .B(_132_), .C(_131_), .Y(_133_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_127_) );
AND2X2 AND2X2_13 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_128_) );
OAI21X1 OAI21X1_19 ( .A(_127_), .B(_128_), .C(w_C_11_), .Y(_129_) );
NAND2X1 NAND2X1_32 ( .A(_129_), .B(_133_), .Y(_77__11_) );
INVX1 INVX1_38 ( .A(w_C_12_), .Y(_137_) );
OR2X2 OR2X2_16 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_138_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_139_) );
NAND3X1 NAND3X1_24 ( .A(_137_), .B(_139_), .C(_138_), .Y(_140_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_134_) );
AND2X2 AND2X2_14 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_135_) );
OAI21X1 OAI21X1_20 ( .A(_134_), .B(_135_), .C(w_C_12_), .Y(_136_) );
NAND2X1 NAND2X1_34 ( .A(_136_), .B(_140_), .Y(_77__12_) );
INVX1 INVX1_39 ( .A(w_C_13_), .Y(_144_) );
OR2X2 OR2X2_17 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_145_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_146_) );
NAND3X1 NAND3X1_25 ( .A(_144_), .B(_146_), .C(_145_), .Y(_147_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_141_) );
AND2X2 AND2X2_15 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_142_) );
OAI21X1 OAI21X1_21 ( .A(_141_), .B(_142_), .C(w_C_13_), .Y(_143_) );
NAND2X1 NAND2X1_36 ( .A(_143_), .B(_147_), .Y(_77__13_) );
INVX1 INVX1_40 ( .A(w_C_14_), .Y(_151_) );
OR2X2 OR2X2_18 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_152_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_153_) );
NAND3X1 NAND3X1_26 ( .A(_151_), .B(_153_), .C(_152_), .Y(_154_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_148_) );
AND2X2 AND2X2_16 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_149_) );
OAI21X1 OAI21X1_22 ( .A(_148_), .B(_149_), .C(w_C_14_), .Y(_150_) );
NAND2X1 NAND2X1_38 ( .A(_150_), .B(_154_), .Y(_77__14_) );
INVX1 INVX1_41 ( .A(w_C_15_), .Y(_158_) );
OR2X2 OR2X2_19 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_159_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_160_) );
NAND3X1 NAND3X1_27 ( .A(_158_), .B(_160_), .C(_159_), .Y(_161_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_155_) );
AND2X2 AND2X2_17 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_156_) );
OAI21X1 OAI21X1_23 ( .A(_155_), .B(_156_), .C(w_C_15_), .Y(_157_) );
NAND2X1 NAND2X1_40 ( .A(_157_), .B(_161_), .Y(_77__15_) );
INVX1 INVX1_42 ( .A(w_C_16_), .Y(_165_) );
OR2X2 OR2X2_20 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_166_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_167_) );
NAND3X1 NAND3X1_28 ( .A(_165_), .B(_167_), .C(_166_), .Y(_168_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_162_) );
AND2X2 AND2X2_18 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_163_) );
OAI21X1 OAI21X1_24 ( .A(_162_), .B(_163_), .C(w_C_16_), .Y(_164_) );
NAND2X1 NAND2X1_42 ( .A(_164_), .B(_168_), .Y(_77__16_) );
INVX1 INVX1_43 ( .A(gnd), .Y(_172_) );
OR2X2 OR2X2_21 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_173_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_174_) );
NAND3X1 NAND3X1_29 ( .A(_172_), .B(_174_), .C(_173_), .Y(_175_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_169_) );
AND2X2 AND2X2_19 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_170_) );
OAI21X1 OAI21X1_25 ( .A(_169_), .B(_170_), .C(gnd), .Y(_171_) );
NAND2X1 NAND2X1_44 ( .A(_171_), .B(_175_), .Y(_77__0_) );
INVX1 INVX1_44 ( .A(w_C_1_), .Y(_179_) );
OR2X2 OR2X2_22 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_180_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_181_) );
NAND3X1 NAND3X1_30 ( .A(_179_), .B(_181_), .C(_180_), .Y(_182_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_176_) );
AND2X2 AND2X2_20 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_177_) );
OAI21X1 OAI21X1_26 ( .A(_176_), .B(_177_), .C(w_C_1_), .Y(_178_) );
NAND2X1 NAND2X1_46 ( .A(_178_), .B(_182_), .Y(_77__1_) );
INVX1 INVX1_45 ( .A(w_C_2_), .Y(_186_) );
OR2X2 OR2X2_23 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_187_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_188_) );
NAND3X1 NAND3X1_31 ( .A(_186_), .B(_188_), .C(_187_), .Y(_189_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_183_) );
AND2X2 AND2X2_21 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_184_) );
OAI21X1 OAI21X1_27 ( .A(_183_), .B(_184_), .C(w_C_2_), .Y(_185_) );
NAND2X1 NAND2X1_48 ( .A(_185_), .B(_189_), .Y(_77__2_) );
INVX1 INVX1_46 ( .A(w_C_3_), .Y(_193_) );
OR2X2 OR2X2_24 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_194_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_195_) );
NAND3X1 NAND3X1_32 ( .A(_193_), .B(_195_), .C(_194_), .Y(_196_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_190_) );
AND2X2 AND2X2_22 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_191_) );
OAI21X1 OAI21X1_28 ( .A(_190_), .B(_191_), .C(w_C_3_), .Y(_192_) );
NAND2X1 NAND2X1_50 ( .A(_192_), .B(_196_), .Y(_77__3_) );
BUFX2 BUFX2_19 ( .A(w_C_17_), .Y(_77__17_) );
BUFX2 BUFX2_20 ( .A(gnd), .Y(w_C_0_) );
endmodule
