module CSkipA_16bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_3_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
INVX1 INVX1_1 ( .A(skip0_cin_next), .Y(_13_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_14_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_15_) );
NAND3X1 NAND3X1_1 ( .A(_13_), .B(_15_), .C(_14_), .Y(_16_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_10_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_11_) );
OAI21X1 OAI21X1_1 ( .A(_10_), .B(_11_), .C(skip0_cin_next), .Y(_12_) );
NAND2X1 NAND2X1_2 ( .A(_12_), .B(_16_), .Y(_0__4_) );
OAI21X1 OAI21X1_2 ( .A(_13_), .B(_10_), .C(_15_), .Y(_2__1_) );
INVX1 INVX1_2 ( .A(_2__3_), .Y(_20_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_21_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_22_) );
NAND3X1 NAND3X1_2 ( .A(_20_), .B(_22_), .C(_21_), .Y(_23_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_17_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_18_) );
OAI21X1 OAI21X1_3 ( .A(_17_), .B(_18_), .C(_2__3_), .Y(_19_) );
NAND2X1 NAND2X1_4 ( .A(_19_), .B(_23_), .Y(_0__7_) );
OAI21X1 OAI21X1_4 ( .A(_20_), .B(_17_), .C(_22_), .Y(_1_) );
INVX1 INVX1_3 ( .A(_2__1_), .Y(_27_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_28_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_29_) );
NAND3X1 NAND3X1_3 ( .A(_27_), .B(_29_), .C(_28_), .Y(_30_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_24_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_25_) );
OAI21X1 OAI21X1_5 ( .A(_24_), .B(_25_), .C(_2__1_), .Y(_26_) );
NAND2X1 NAND2X1_6 ( .A(_26_), .B(_30_), .Y(_0__5_) );
OAI21X1 OAI21X1_6 ( .A(_27_), .B(_24_), .C(_29_), .Y(_2__2_) );
INVX1 INVX1_4 ( .A(_2__2_), .Y(_34_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_35_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_36_) );
NAND3X1 NAND3X1_4 ( .A(_34_), .B(_36_), .C(_35_), .Y(_37_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_31_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_32_) );
OAI21X1 OAI21X1_7 ( .A(_31_), .B(_32_), .C(_2__2_), .Y(_33_) );
NAND2X1 NAND2X1_8 ( .A(_33_), .B(_37_), .Y(_0__6_) );
OAI21X1 OAI21X1_8 ( .A(_34_), .B(_31_), .C(_36_), .Y(_2__3_) );
INVX1 INVX1_5 ( .A(i_add_term2[4]), .Y(_38_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term1[4]), .B(_38_), .Y(_39_) );
INVX1 INVX1_6 ( .A(i_add_term1[4]), .Y(_40_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[4]), .B(_40_), .Y(_41_) );
INVX1 INVX1_7 ( .A(i_add_term1[5]), .Y(_42_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[5]), .B(_42_), .Y(_43_) );
INVX1 INVX1_8 ( .A(i_add_term2[5]), .Y(_44_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term1[5]), .B(_44_), .Y(_45_) );
OAI22X1 OAI22X1_1 ( .A(_39_), .B(_41_), .C(_43_), .D(_45_), .Y(_46_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_47_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_48_) );
NOR2X1 NOR2X1_10 ( .A(_47_), .B(_48_), .Y(_49_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_50_) );
NAND2X1 NAND2X1_9 ( .A(_49_), .B(_50_), .Y(_51_) );
NOR2X1 NOR2X1_11 ( .A(_46_), .B(_51_), .Y(_3_) );
INVX1 INVX1_9 ( .A(_1_), .Y(_52_) );
NAND2X1 NAND2X1_10 ( .A(1'b0), .B(_3_), .Y(_53_) );
OAI21X1 OAI21X1_9 ( .A(_3_), .B(_52_), .C(_53_), .Y(w_cout_1_) );
INVX1 INVX1_10 ( .A(w_cout_1_), .Y(_57_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_58_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_59_) );
NAND3X1 NAND3X1_5 ( .A(_57_), .B(_59_), .C(_58_), .Y(_60_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_54_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_55_) );
OAI21X1 OAI21X1_10 ( .A(_54_), .B(_55_), .C(w_cout_1_), .Y(_56_) );
NAND2X1 NAND2X1_12 ( .A(_56_), .B(_60_), .Y(_0__8_) );
OAI21X1 OAI21X1_11 ( .A(_57_), .B(_54_), .C(_59_), .Y(_5__1_) );
INVX1 INVX1_11 ( .A(_5__3_), .Y(_64_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_65_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_66_) );
NAND3X1 NAND3X1_6 ( .A(_64_), .B(_66_), .C(_65_), .Y(_67_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_61_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_62_) );
OAI21X1 OAI21X1_12 ( .A(_61_), .B(_62_), .C(_5__3_), .Y(_63_) );
NAND2X1 NAND2X1_14 ( .A(_63_), .B(_67_), .Y(_0__11_) );
OAI21X1 OAI21X1_13 ( .A(_64_), .B(_61_), .C(_66_), .Y(_4_) );
INVX1 INVX1_12 ( .A(_5__1_), .Y(_71_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_72_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_73_) );
NAND3X1 NAND3X1_7 ( .A(_71_), .B(_73_), .C(_72_), .Y(_74_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_68_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_69_) );
OAI21X1 OAI21X1_14 ( .A(_68_), .B(_69_), .C(_5__1_), .Y(_70_) );
NAND2X1 NAND2X1_16 ( .A(_70_), .B(_74_), .Y(_0__9_) );
OAI21X1 OAI21X1_15 ( .A(_71_), .B(_68_), .C(_73_), .Y(_5__2_) );
INVX1 INVX1_13 ( .A(_5__2_), .Y(_78_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_79_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_80_) );
NAND3X1 NAND3X1_8 ( .A(_78_), .B(_80_), .C(_79_), .Y(_81_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_75_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_76_) );
OAI21X1 OAI21X1_16 ( .A(_75_), .B(_76_), .C(_5__2_), .Y(_77_) );
NAND2X1 NAND2X1_18 ( .A(_77_), .B(_81_), .Y(_0__10_) );
OAI21X1 OAI21X1_17 ( .A(_78_), .B(_75_), .C(_80_), .Y(_5__3_) );
INVX1 INVX1_14 ( .A(i_add_term2[8]), .Y(_82_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term1[8]), .B(_82_), .Y(_83_) );
INVX1 INVX1_15 ( .A(i_add_term1[8]), .Y(_84_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[8]), .B(_84_), .Y(_85_) );
INVX1 INVX1_16 ( .A(i_add_term1[9]), .Y(_86_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[9]), .B(_86_), .Y(_87_) );
INVX1 INVX1_17 ( .A(i_add_term2[9]), .Y(_88_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term1[9]), .B(_88_), .Y(_89_) );
OAI22X1 OAI22X1_2 ( .A(_83_), .B(_85_), .C(_87_), .D(_89_), .Y(_90_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_91_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_92_) );
NOR2X1 NOR2X1_21 ( .A(_91_), .B(_92_), .Y(_93_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_94_) );
NAND2X1 NAND2X1_19 ( .A(_93_), .B(_94_), .Y(_95_) );
NOR2X1 NOR2X1_22 ( .A(_90_), .B(_95_), .Y(_6_) );
INVX1 INVX1_18 ( .A(_4_), .Y(_96_) );
NAND2X1 NAND2X1_20 ( .A(1'b0), .B(_6_), .Y(_97_) );
OAI21X1 OAI21X1_18 ( .A(_6_), .B(_96_), .C(_97_), .Y(w_cout_2_) );
INVX1 INVX1_19 ( .A(w_cout_2_), .Y(_101_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_102_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_103_) );
NAND3X1 NAND3X1_9 ( .A(_101_), .B(_103_), .C(_102_), .Y(_104_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_98_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_99_) );
OAI21X1 OAI21X1_19 ( .A(_98_), .B(_99_), .C(w_cout_2_), .Y(_100_) );
NAND2X1 NAND2X1_22 ( .A(_100_), .B(_104_), .Y(_0__12_) );
OAI21X1 OAI21X1_20 ( .A(_101_), .B(_98_), .C(_103_), .Y(_8__1_) );
INVX1 INVX1_20 ( .A(_8__3_), .Y(_108_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_109_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_110_) );
NAND3X1 NAND3X1_10 ( .A(_108_), .B(_110_), .C(_109_), .Y(_111_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_105_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_106_) );
OAI21X1 OAI21X1_21 ( .A(_105_), .B(_106_), .C(_8__3_), .Y(_107_) );
NAND2X1 NAND2X1_24 ( .A(_107_), .B(_111_), .Y(_0__15_) );
OAI21X1 OAI21X1_22 ( .A(_108_), .B(_105_), .C(_110_), .Y(_7_) );
INVX1 INVX1_21 ( .A(_8__1_), .Y(_115_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_116_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_117_) );
NAND3X1 NAND3X1_11 ( .A(_115_), .B(_117_), .C(_116_), .Y(_118_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_112_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_113_) );
OAI21X1 OAI21X1_23 ( .A(_112_), .B(_113_), .C(_8__1_), .Y(_114_) );
NAND2X1 NAND2X1_26 ( .A(_114_), .B(_118_), .Y(_0__13_) );
OAI21X1 OAI21X1_24 ( .A(_115_), .B(_112_), .C(_117_), .Y(_8__2_) );
INVX1 INVX1_22 ( .A(_8__2_), .Y(_122_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_123_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_124_) );
NAND3X1 NAND3X1_12 ( .A(_122_), .B(_124_), .C(_123_), .Y(_125_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_119_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_120_) );
OAI21X1 OAI21X1_25 ( .A(_119_), .B(_120_), .C(_8__2_), .Y(_121_) );
NAND2X1 NAND2X1_28 ( .A(_121_), .B(_125_), .Y(_0__14_) );
OAI21X1 OAI21X1_26 ( .A(_122_), .B(_119_), .C(_124_), .Y(_8__3_) );
INVX1 INVX1_23 ( .A(i_add_term2[12]), .Y(_126_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term1[12]), .B(_126_), .Y(_127_) );
INVX1 INVX1_24 ( .A(i_add_term1[12]), .Y(_128_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[12]), .B(_128_), .Y(_129_) );
INVX1 INVX1_25 ( .A(i_add_term1[13]), .Y(_130_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[13]), .B(_130_), .Y(_131_) );
INVX1 INVX1_26 ( .A(i_add_term2[13]), .Y(_132_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term1[13]), .B(_132_), .Y(_133_) );
OAI22X1 OAI22X1_3 ( .A(_127_), .B(_129_), .C(_131_), .D(_133_), .Y(_134_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_135_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_136_) );
NOR2X1 NOR2X1_32 ( .A(_135_), .B(_136_), .Y(_137_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_138_) );
NAND2X1 NAND2X1_29 ( .A(_137_), .B(_138_), .Y(_139_) );
NOR2X1 NOR2X1_33 ( .A(_134_), .B(_139_), .Y(_9_) );
INVX1 INVX1_27 ( .A(_7_), .Y(_140_) );
NAND2X1 NAND2X1_30 ( .A(1'b0), .B(_9_), .Y(_141_) );
OAI21X1 OAI21X1_27 ( .A(_9_), .B(_140_), .C(_141_), .Y(w_cout_3_) );
INVX1 INVX1_28 ( .A(1'b0), .Y(_145_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_146_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_147_) );
NAND3X1 NAND3X1_13 ( .A(_145_), .B(_147_), .C(_146_), .Y(_148_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_142_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_143_) );
OAI21X1 OAI21X1_28 ( .A(_142_), .B(_143_), .C(1'b0), .Y(_144_) );
NAND2X1 NAND2X1_32 ( .A(_144_), .B(_148_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_29 ( .A(_145_), .B(_142_), .C(_147_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_29 ( .A(rca_inst_fa3_i_carry), .Y(_152_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_153_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_154_) );
NAND3X1 NAND3X1_14 ( .A(_152_), .B(_154_), .C(_153_), .Y(_155_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_149_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_150_) );
OAI21X1 OAI21X1_30 ( .A(_149_), .B(_150_), .C(rca_inst_fa3_i_carry), .Y(_151_) );
NAND2X1 NAND2X1_34 ( .A(_151_), .B(_155_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_31 ( .A(_152_), .B(_149_), .C(_154_), .Y(cout0) );
INVX1 INVX1_30 ( .A(rca_inst_fa0_o_carry), .Y(_159_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_160_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_161_) );
NAND3X1 NAND3X1_15 ( .A(_159_), .B(_161_), .C(_160_), .Y(_162_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_156_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_157_) );
OAI21X1 OAI21X1_32 ( .A(_156_), .B(_157_), .C(rca_inst_fa0_o_carry), .Y(_158_) );
NAND2X1 NAND2X1_36 ( .A(_158_), .B(_162_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_33 ( .A(_159_), .B(_156_), .C(_161_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_31 ( .A(rca_inst_fa_1__o_carry), .Y(_166_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_167_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_168_) );
NAND3X1 NAND3X1_16 ( .A(_166_), .B(_168_), .C(_167_), .Y(_169_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_163_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_164_) );
OAI21X1 OAI21X1_34 ( .A(_163_), .B(_164_), .C(rca_inst_fa_1__o_carry), .Y(_165_) );
NAND2X1 NAND2X1_38 ( .A(_165_), .B(_169_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_35 ( .A(_166_), .B(_163_), .C(_168_), .Y(rca_inst_fa3_i_carry) );
INVX1 INVX1_32 ( .A(i_add_term2[0]), .Y(_170_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term1[0]), .B(_170_), .Y(_171_) );
INVX1 INVX1_33 ( .A(i_add_term1[0]), .Y(_172_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[0]), .B(_172_), .Y(_173_) );
INVX1 INVX1_34 ( .A(i_add_term1[1]), .Y(_174_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[1]), .B(_174_), .Y(_175_) );
INVX1 INVX1_35 ( .A(i_add_term2[1]), .Y(_176_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term1[1]), .B(_176_), .Y(_177_) );
OAI22X1 OAI22X1_4 ( .A(_171_), .B(_173_), .C(_175_), .D(_177_), .Y(_178_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_179_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_180_) );
NOR2X1 NOR2X1_43 ( .A(_179_), .B(_180_), .Y(_181_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_182_) );
NAND2X1 NAND2X1_39 ( .A(_181_), .B(_182_), .Y(_183_) );
NOR2X1 NOR2X1_44 ( .A(_178_), .B(_183_), .Y(skip0_P) );
INVX1 INVX1_36 ( .A(cout0), .Y(_184_) );
NAND2X1 NAND2X1_40 ( .A(1'b0), .B(skip0_P), .Y(_185_) );
OAI21X1 OAI21X1_36 ( .A(skip0_P), .B(_184_), .C(_185_), .Y(skip0_cin_next) );
BUFX2 BUFX2_18 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_19 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_20 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_21 ( .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_22 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
