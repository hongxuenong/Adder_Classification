module csa_25bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_6_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(csa_inst_mux0_sum_y), .Y(sum[24]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_31_) );
NAND2X1 NAND2X1_1 ( .A(_2_), .B(rca_inst_cout), .Y(_32_) );
OAI21X1 OAI21X1_1 ( .A(rca_inst_cout), .B(_31_), .C(_32_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3__2_), .Y(_33_) );
NAND2X1 NAND2X1_2 ( .A(_4__2_), .B(rca_inst_cout), .Y(_34_) );
OAI21X1 OAI21X1_2 ( .A(rca_inst_cout), .B(_33_), .C(_34_), .Y(_0__6_) );
INVX1 INVX1_3 ( .A(_3__3_), .Y(_35_) );
NAND2X1 NAND2X1_3 ( .A(rca_inst_cout), .B(_4__3_), .Y(_36_) );
OAI21X1 OAI21X1_3 ( .A(rca_inst_cout), .B(_35_), .C(_36_), .Y(_0__7_) );
INVX1 INVX1_4 ( .A(_3__0_), .Y(_37_) );
NAND2X1 NAND2X1_4 ( .A(rca_inst_cout), .B(_4__0_), .Y(_38_) );
OAI21X1 OAI21X1_4 ( .A(rca_inst_cout), .B(_37_), .C(_38_), .Y(_0__4_) );
INVX1 INVX1_5 ( .A(_3__1_), .Y(_39_) );
NAND2X1 NAND2X1_5 ( .A(rca_inst_cout), .B(_4__1_), .Y(_40_) );
OAI21X1 OAI21X1_5 ( .A(rca_inst_cout), .B(_39_), .C(_40_), .Y(_0__5_) );
INVX1 INVX1_6 ( .A(1'b0), .Y(_44_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_45_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_46_) );
NAND3X1 NAND3X1_1 ( .A(_44_), .B(_46_), .C(_45_), .Y(_47_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_41_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_42_) );
OAI21X1 OAI21X1_6 ( .A(_41_), .B(_42_), .C(1'b0), .Y(_43_) );
NAND2X1 NAND2X1_7 ( .A(_43_), .B(_47_), .Y(_3__0_) );
OAI21X1 OAI21X1_7 ( .A(_44_), .B(_41_), .C(_46_), .Y(_5__1_) );
INVX1 INVX1_7 ( .A(_5__3_), .Y(_51_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_52_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_53_) );
NAND3X1 NAND3X1_2 ( .A(_51_), .B(_53_), .C(_52_), .Y(_54_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_48_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_49_) );
OAI21X1 OAI21X1_8 ( .A(_48_), .B(_49_), .C(_5__3_), .Y(_50_) );
NAND2X1 NAND2X1_9 ( .A(_50_), .B(_54_), .Y(_3__3_) );
OAI21X1 OAI21X1_9 ( .A(_51_), .B(_48_), .C(_53_), .Y(_1_) );
INVX1 INVX1_8 ( .A(_5__1_), .Y(_58_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_59_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_60_) );
NAND3X1 NAND3X1_3 ( .A(_58_), .B(_60_), .C(_59_), .Y(_61_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_55_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_56_) );
OAI21X1 OAI21X1_10 ( .A(_55_), .B(_56_), .C(_5__1_), .Y(_57_) );
NAND2X1 NAND2X1_11 ( .A(_57_), .B(_61_), .Y(_3__1_) );
OAI21X1 OAI21X1_11 ( .A(_58_), .B(_55_), .C(_60_), .Y(_5__2_) );
INVX1 INVX1_9 ( .A(_5__2_), .Y(_65_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_66_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_67_) );
NAND3X1 NAND3X1_4 ( .A(_65_), .B(_67_), .C(_66_), .Y(_68_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_62_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_63_) );
OAI21X1 OAI21X1_12 ( .A(_62_), .B(_63_), .C(_5__2_), .Y(_64_) );
NAND2X1 NAND2X1_13 ( .A(_64_), .B(_68_), .Y(_3__2_) );
OAI21X1 OAI21X1_13 ( .A(_65_), .B(_62_), .C(_67_), .Y(_5__3_) );
INVX1 INVX1_10 ( .A(1'b1), .Y(_72_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_73_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_74_) );
NAND3X1 NAND3X1_5 ( .A(_72_), .B(_74_), .C(_73_), .Y(_75_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_69_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_70_) );
OAI21X1 OAI21X1_14 ( .A(_69_), .B(_70_), .C(1'b1), .Y(_71_) );
NAND2X1 NAND2X1_15 ( .A(_71_), .B(_75_), .Y(_4__0_) );
OAI21X1 OAI21X1_15 ( .A(_72_), .B(_69_), .C(_74_), .Y(_6__1_) );
INVX1 INVX1_11 ( .A(_6__3_), .Y(_79_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_80_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_81_) );
NAND3X1 NAND3X1_6 ( .A(_79_), .B(_81_), .C(_80_), .Y(_82_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_76_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_77_) );
OAI21X1 OAI21X1_16 ( .A(_76_), .B(_77_), .C(_6__3_), .Y(_78_) );
NAND2X1 NAND2X1_17 ( .A(_78_), .B(_82_), .Y(_4__3_) );
OAI21X1 OAI21X1_17 ( .A(_79_), .B(_76_), .C(_81_), .Y(_2_) );
INVX1 INVX1_12 ( .A(_6__1_), .Y(_86_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_87_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_88_) );
NAND3X1 NAND3X1_7 ( .A(_86_), .B(_88_), .C(_87_), .Y(_89_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_83_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_84_) );
OAI21X1 OAI21X1_18 ( .A(_83_), .B(_84_), .C(_6__1_), .Y(_85_) );
NAND2X1 NAND2X1_19 ( .A(_85_), .B(_89_), .Y(_4__1_) );
OAI21X1 OAI21X1_19 ( .A(_86_), .B(_83_), .C(_88_), .Y(_6__2_) );
INVX1 INVX1_13 ( .A(_6__2_), .Y(_93_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_94_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_95_) );
NAND3X1 NAND3X1_8 ( .A(_93_), .B(_95_), .C(_94_), .Y(_96_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_90_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_91_) );
OAI21X1 OAI21X1_20 ( .A(_90_), .B(_91_), .C(_6__2_), .Y(_92_) );
NAND2X1 NAND2X1_21 ( .A(_92_), .B(_96_), .Y(_4__2_) );
OAI21X1 OAI21X1_21 ( .A(_93_), .B(_90_), .C(_95_), .Y(_6__3_) );
INVX1 INVX1_14 ( .A(_7_), .Y(_97_) );
NAND2X1 NAND2X1_22 ( .A(_8_), .B(w_cout_1_), .Y(_98_) );
OAI21X1 OAI21X1_22 ( .A(w_cout_1_), .B(_97_), .C(_98_), .Y(w_cout_2_) );
INVX1 INVX1_15 ( .A(_9__2_), .Y(_99_) );
NAND2X1 NAND2X1_23 ( .A(_10__2_), .B(w_cout_1_), .Y(_100_) );
OAI21X1 OAI21X1_23 ( .A(w_cout_1_), .B(_99_), .C(_100_), .Y(_0__10_) );
INVX1 INVX1_16 ( .A(_9__3_), .Y(_101_) );
NAND2X1 NAND2X1_24 ( .A(w_cout_1_), .B(_10__3_), .Y(_102_) );
OAI21X1 OAI21X1_24 ( .A(w_cout_1_), .B(_101_), .C(_102_), .Y(_0__11_) );
INVX1 INVX1_17 ( .A(_9__0_), .Y(_103_) );
NAND2X1 NAND2X1_25 ( .A(w_cout_1_), .B(_10__0_), .Y(_104_) );
OAI21X1 OAI21X1_25 ( .A(w_cout_1_), .B(_103_), .C(_104_), .Y(_0__8_) );
INVX1 INVX1_18 ( .A(_9__1_), .Y(_105_) );
NAND2X1 NAND2X1_26 ( .A(w_cout_1_), .B(_10__1_), .Y(_106_) );
OAI21X1 OAI21X1_26 ( .A(w_cout_1_), .B(_105_), .C(_106_), .Y(_0__9_) );
INVX1 INVX1_19 ( .A(1'b0), .Y(_110_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_111_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_112_) );
NAND3X1 NAND3X1_9 ( .A(_110_), .B(_112_), .C(_111_), .Y(_113_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_107_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_108_) );
OAI21X1 OAI21X1_27 ( .A(_107_), .B(_108_), .C(1'b0), .Y(_109_) );
NAND2X1 NAND2X1_28 ( .A(_109_), .B(_113_), .Y(_9__0_) );
OAI21X1 OAI21X1_28 ( .A(_110_), .B(_107_), .C(_112_), .Y(_11__1_) );
INVX1 INVX1_20 ( .A(_11__3_), .Y(_117_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_118_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_119_) );
NAND3X1 NAND3X1_10 ( .A(_117_), .B(_119_), .C(_118_), .Y(_120_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_114_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_115_) );
OAI21X1 OAI21X1_29 ( .A(_114_), .B(_115_), .C(_11__3_), .Y(_116_) );
NAND2X1 NAND2X1_30 ( .A(_116_), .B(_120_), .Y(_9__3_) );
OAI21X1 OAI21X1_30 ( .A(_117_), .B(_114_), .C(_119_), .Y(_7_) );
INVX1 INVX1_21 ( .A(_11__1_), .Y(_124_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_125_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_126_) );
NAND3X1 NAND3X1_11 ( .A(_124_), .B(_126_), .C(_125_), .Y(_127_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_121_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_122_) );
OAI21X1 OAI21X1_31 ( .A(_121_), .B(_122_), .C(_11__1_), .Y(_123_) );
NAND2X1 NAND2X1_32 ( .A(_123_), .B(_127_), .Y(_9__1_) );
OAI21X1 OAI21X1_32 ( .A(_124_), .B(_121_), .C(_126_), .Y(_11__2_) );
INVX1 INVX1_22 ( .A(_11__2_), .Y(_131_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_132_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_133_) );
NAND3X1 NAND3X1_12 ( .A(_131_), .B(_133_), .C(_132_), .Y(_134_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_128_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_129_) );
OAI21X1 OAI21X1_33 ( .A(_128_), .B(_129_), .C(_11__2_), .Y(_130_) );
NAND2X1 NAND2X1_34 ( .A(_130_), .B(_134_), .Y(_9__2_) );
OAI21X1 OAI21X1_34 ( .A(_131_), .B(_128_), .C(_133_), .Y(_11__3_) );
INVX1 INVX1_23 ( .A(1'b1), .Y(_138_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_139_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_140_) );
NAND3X1 NAND3X1_13 ( .A(_138_), .B(_140_), .C(_139_), .Y(_141_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_135_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_136_) );
OAI21X1 OAI21X1_35 ( .A(_135_), .B(_136_), .C(1'b1), .Y(_137_) );
NAND2X1 NAND2X1_36 ( .A(_137_), .B(_141_), .Y(_10__0_) );
OAI21X1 OAI21X1_36 ( .A(_138_), .B(_135_), .C(_140_), .Y(_12__1_) );
INVX1 INVX1_24 ( .A(_12__3_), .Y(_145_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_146_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_147_) );
NAND3X1 NAND3X1_14 ( .A(_145_), .B(_147_), .C(_146_), .Y(_148_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_142_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_143_) );
OAI21X1 OAI21X1_37 ( .A(_142_), .B(_143_), .C(_12__3_), .Y(_144_) );
NAND2X1 NAND2X1_38 ( .A(_144_), .B(_148_), .Y(_10__3_) );
OAI21X1 OAI21X1_38 ( .A(_145_), .B(_142_), .C(_147_), .Y(_8_) );
INVX1 INVX1_25 ( .A(_12__1_), .Y(_152_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_153_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_154_) );
NAND3X1 NAND3X1_15 ( .A(_152_), .B(_154_), .C(_153_), .Y(_155_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_149_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_150_) );
OAI21X1 OAI21X1_39 ( .A(_149_), .B(_150_), .C(_12__1_), .Y(_151_) );
NAND2X1 NAND2X1_40 ( .A(_151_), .B(_155_), .Y(_10__1_) );
OAI21X1 OAI21X1_40 ( .A(_152_), .B(_149_), .C(_154_), .Y(_12__2_) );
INVX1 INVX1_26 ( .A(_12__2_), .Y(_159_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_160_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_161_) );
NAND3X1 NAND3X1_16 ( .A(_159_), .B(_161_), .C(_160_), .Y(_162_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_156_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_157_) );
OAI21X1 OAI21X1_41 ( .A(_156_), .B(_157_), .C(_12__2_), .Y(_158_) );
NAND2X1 NAND2X1_42 ( .A(_158_), .B(_162_), .Y(_10__2_) );
OAI21X1 OAI21X1_42 ( .A(_159_), .B(_156_), .C(_161_), .Y(_12__3_) );
INVX1 INVX1_27 ( .A(_13_), .Y(_163_) );
NAND2X1 NAND2X1_43 ( .A(_14_), .B(w_cout_2_), .Y(_164_) );
OAI21X1 OAI21X1_43 ( .A(w_cout_2_), .B(_163_), .C(_164_), .Y(w_cout_3_) );
INVX1 INVX1_28 ( .A(_15__2_), .Y(_165_) );
NAND2X1 NAND2X1_44 ( .A(_16__2_), .B(w_cout_2_), .Y(_166_) );
OAI21X1 OAI21X1_44 ( .A(w_cout_2_), .B(_165_), .C(_166_), .Y(_0__14_) );
INVX1 INVX1_29 ( .A(_15__3_), .Y(_167_) );
NAND2X1 NAND2X1_45 ( .A(w_cout_2_), .B(_16__3_), .Y(_168_) );
OAI21X1 OAI21X1_45 ( .A(w_cout_2_), .B(_167_), .C(_168_), .Y(_0__15_) );
INVX1 INVX1_30 ( .A(_15__0_), .Y(_169_) );
NAND2X1 NAND2X1_46 ( .A(w_cout_2_), .B(_16__0_), .Y(_170_) );
OAI21X1 OAI21X1_46 ( .A(w_cout_2_), .B(_169_), .C(_170_), .Y(_0__12_) );
INVX1 INVX1_31 ( .A(_15__1_), .Y(_171_) );
NAND2X1 NAND2X1_47 ( .A(w_cout_2_), .B(_16__1_), .Y(_172_) );
OAI21X1 OAI21X1_47 ( .A(w_cout_2_), .B(_171_), .C(_172_), .Y(_0__13_) );
INVX1 INVX1_32 ( .A(1'b0), .Y(_176_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_177_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_178_) );
NAND3X1 NAND3X1_17 ( .A(_176_), .B(_178_), .C(_177_), .Y(_179_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_173_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_174_) );
OAI21X1 OAI21X1_48 ( .A(_173_), .B(_174_), .C(1'b0), .Y(_175_) );
NAND2X1 NAND2X1_49 ( .A(_175_), .B(_179_), .Y(_15__0_) );
OAI21X1 OAI21X1_49 ( .A(_176_), .B(_173_), .C(_178_), .Y(_17__1_) );
INVX1 INVX1_33 ( .A(_17__3_), .Y(_183_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_184_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_185_) );
NAND3X1 NAND3X1_18 ( .A(_183_), .B(_185_), .C(_184_), .Y(_186_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_180_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_181_) );
OAI21X1 OAI21X1_50 ( .A(_180_), .B(_181_), .C(_17__3_), .Y(_182_) );
NAND2X1 NAND2X1_51 ( .A(_182_), .B(_186_), .Y(_15__3_) );
OAI21X1 OAI21X1_51 ( .A(_183_), .B(_180_), .C(_185_), .Y(_13_) );
INVX1 INVX1_34 ( .A(_17__1_), .Y(_190_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_191_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_192_) );
NAND3X1 NAND3X1_19 ( .A(_190_), .B(_192_), .C(_191_), .Y(_193_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_187_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_188_) );
OAI21X1 OAI21X1_52 ( .A(_187_), .B(_188_), .C(_17__1_), .Y(_189_) );
NAND2X1 NAND2X1_53 ( .A(_189_), .B(_193_), .Y(_15__1_) );
OAI21X1 OAI21X1_53 ( .A(_190_), .B(_187_), .C(_192_), .Y(_17__2_) );
INVX1 INVX1_35 ( .A(_17__2_), .Y(_197_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_198_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_199_) );
NAND3X1 NAND3X1_20 ( .A(_197_), .B(_199_), .C(_198_), .Y(_200_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_194_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_195_) );
OAI21X1 OAI21X1_54 ( .A(_194_), .B(_195_), .C(_17__2_), .Y(_196_) );
NAND2X1 NAND2X1_55 ( .A(_196_), .B(_200_), .Y(_15__2_) );
OAI21X1 OAI21X1_55 ( .A(_197_), .B(_194_), .C(_199_), .Y(_17__3_) );
INVX1 INVX1_36 ( .A(1'b1), .Y(_204_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_205_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_206_) );
NAND3X1 NAND3X1_21 ( .A(_204_), .B(_206_), .C(_205_), .Y(_207_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_201_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_202_) );
OAI21X1 OAI21X1_56 ( .A(_201_), .B(_202_), .C(1'b1), .Y(_203_) );
NAND2X1 NAND2X1_57 ( .A(_203_), .B(_207_), .Y(_16__0_) );
OAI21X1 OAI21X1_57 ( .A(_204_), .B(_201_), .C(_206_), .Y(_18__1_) );
INVX1 INVX1_37 ( .A(_18__3_), .Y(_211_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_212_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_213_) );
NAND3X1 NAND3X1_22 ( .A(_211_), .B(_213_), .C(_212_), .Y(_214_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_208_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_209_) );
OAI21X1 OAI21X1_58 ( .A(_208_), .B(_209_), .C(_18__3_), .Y(_210_) );
NAND2X1 NAND2X1_59 ( .A(_210_), .B(_214_), .Y(_16__3_) );
OAI21X1 OAI21X1_59 ( .A(_211_), .B(_208_), .C(_213_), .Y(_14_) );
INVX1 INVX1_38 ( .A(_18__1_), .Y(_218_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_219_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_220_) );
NAND3X1 NAND3X1_23 ( .A(_218_), .B(_220_), .C(_219_), .Y(_221_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_215_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_216_) );
OAI21X1 OAI21X1_60 ( .A(_215_), .B(_216_), .C(_18__1_), .Y(_217_) );
NAND2X1 NAND2X1_61 ( .A(_217_), .B(_221_), .Y(_16__1_) );
OAI21X1 OAI21X1_61 ( .A(_218_), .B(_215_), .C(_220_), .Y(_18__2_) );
INVX1 INVX1_39 ( .A(_18__2_), .Y(_225_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_226_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_227_) );
NAND3X1 NAND3X1_24 ( .A(_225_), .B(_227_), .C(_226_), .Y(_228_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_222_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_223_) );
OAI21X1 OAI21X1_62 ( .A(_222_), .B(_223_), .C(_18__2_), .Y(_224_) );
NAND2X1 NAND2X1_63 ( .A(_224_), .B(_228_), .Y(_16__2_) );
OAI21X1 OAI21X1_63 ( .A(_225_), .B(_222_), .C(_227_), .Y(_18__3_) );
INVX1 INVX1_40 ( .A(_19_), .Y(_229_) );
NAND2X1 NAND2X1_64 ( .A(_20_), .B(w_cout_3_), .Y(_230_) );
OAI21X1 OAI21X1_64 ( .A(w_cout_3_), .B(_229_), .C(_230_), .Y(w_cout_4_) );
INVX1 INVX1_41 ( .A(_21__2_), .Y(_231_) );
NAND2X1 NAND2X1_65 ( .A(_22__2_), .B(w_cout_3_), .Y(_232_) );
OAI21X1 OAI21X1_65 ( .A(w_cout_3_), .B(_231_), .C(_232_), .Y(_0__18_) );
INVX1 INVX1_42 ( .A(_21__3_), .Y(_233_) );
NAND2X1 NAND2X1_66 ( .A(w_cout_3_), .B(_22__3_), .Y(_234_) );
OAI21X1 OAI21X1_66 ( .A(w_cout_3_), .B(_233_), .C(_234_), .Y(_0__19_) );
INVX1 INVX1_43 ( .A(_21__0_), .Y(_235_) );
NAND2X1 NAND2X1_67 ( .A(w_cout_3_), .B(_22__0_), .Y(_236_) );
OAI21X1 OAI21X1_67 ( .A(w_cout_3_), .B(_235_), .C(_236_), .Y(_0__16_) );
INVX1 INVX1_44 ( .A(_21__1_), .Y(_237_) );
NAND2X1 NAND2X1_68 ( .A(w_cout_3_), .B(_22__1_), .Y(_238_) );
OAI21X1 OAI21X1_68 ( .A(w_cout_3_), .B(_237_), .C(_238_), .Y(_0__17_) );
INVX1 INVX1_45 ( .A(1'b0), .Y(_242_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_243_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_244_) );
NAND3X1 NAND3X1_25 ( .A(_242_), .B(_244_), .C(_243_), .Y(_245_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_239_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_240_) );
OAI21X1 OAI21X1_69 ( .A(_239_), .B(_240_), .C(1'b0), .Y(_241_) );
NAND2X1 NAND2X1_70 ( .A(_241_), .B(_245_), .Y(_21__0_) );
OAI21X1 OAI21X1_70 ( .A(_242_), .B(_239_), .C(_244_), .Y(_23__1_) );
INVX1 INVX1_46 ( .A(_23__3_), .Y(_249_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_250_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_251_) );
NAND3X1 NAND3X1_26 ( .A(_249_), .B(_251_), .C(_250_), .Y(_252_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_246_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_247_) );
OAI21X1 OAI21X1_71 ( .A(_246_), .B(_247_), .C(_23__3_), .Y(_248_) );
NAND2X1 NAND2X1_72 ( .A(_248_), .B(_252_), .Y(_21__3_) );
OAI21X1 OAI21X1_72 ( .A(_249_), .B(_246_), .C(_251_), .Y(_19_) );
INVX1 INVX1_47 ( .A(_23__1_), .Y(_256_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_257_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_258_) );
NAND3X1 NAND3X1_27 ( .A(_256_), .B(_258_), .C(_257_), .Y(_259_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_253_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_254_) );
OAI21X1 OAI21X1_73 ( .A(_253_), .B(_254_), .C(_23__1_), .Y(_255_) );
NAND2X1 NAND2X1_74 ( .A(_255_), .B(_259_), .Y(_21__1_) );
OAI21X1 OAI21X1_74 ( .A(_256_), .B(_253_), .C(_258_), .Y(_23__2_) );
INVX1 INVX1_48 ( .A(_23__2_), .Y(_263_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_264_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_265_) );
NAND3X1 NAND3X1_28 ( .A(_263_), .B(_265_), .C(_264_), .Y(_266_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_260_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_261_) );
OAI21X1 OAI21X1_75 ( .A(_260_), .B(_261_), .C(_23__2_), .Y(_262_) );
NAND2X1 NAND2X1_76 ( .A(_262_), .B(_266_), .Y(_21__2_) );
OAI21X1 OAI21X1_76 ( .A(_263_), .B(_260_), .C(_265_), .Y(_23__3_) );
INVX1 INVX1_49 ( .A(1'b1), .Y(_270_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_271_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_272_) );
NAND3X1 NAND3X1_29 ( .A(_270_), .B(_272_), .C(_271_), .Y(_273_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_267_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_268_) );
OAI21X1 OAI21X1_77 ( .A(_267_), .B(_268_), .C(1'b1), .Y(_269_) );
NAND2X1 NAND2X1_78 ( .A(_269_), .B(_273_), .Y(_22__0_) );
OAI21X1 OAI21X1_78 ( .A(_270_), .B(_267_), .C(_272_), .Y(_24__1_) );
INVX1 INVX1_50 ( .A(_24__3_), .Y(_277_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_278_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_279_) );
NAND3X1 NAND3X1_30 ( .A(_277_), .B(_279_), .C(_278_), .Y(_280_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_274_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_275_) );
OAI21X1 OAI21X1_79 ( .A(_274_), .B(_275_), .C(_24__3_), .Y(_276_) );
NAND2X1 NAND2X1_80 ( .A(_276_), .B(_280_), .Y(_22__3_) );
OAI21X1 OAI21X1_80 ( .A(_277_), .B(_274_), .C(_279_), .Y(_20_) );
INVX1 INVX1_51 ( .A(_24__1_), .Y(_284_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_285_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_286_) );
NAND3X1 NAND3X1_31 ( .A(_284_), .B(_286_), .C(_285_), .Y(_287_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_281_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_282_) );
OAI21X1 OAI21X1_81 ( .A(_281_), .B(_282_), .C(_24__1_), .Y(_283_) );
NAND2X1 NAND2X1_82 ( .A(_283_), .B(_287_), .Y(_22__1_) );
OAI21X1 OAI21X1_82 ( .A(_284_), .B(_281_), .C(_286_), .Y(_24__2_) );
INVX1 INVX1_52 ( .A(_24__2_), .Y(_291_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_292_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_293_) );
NAND3X1 NAND3X1_32 ( .A(_291_), .B(_293_), .C(_292_), .Y(_294_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_288_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_289_) );
OAI21X1 OAI21X1_83 ( .A(_288_), .B(_289_), .C(_24__2_), .Y(_290_) );
NAND2X1 NAND2X1_84 ( .A(_290_), .B(_294_), .Y(_22__2_) );
OAI21X1 OAI21X1_84 ( .A(_291_), .B(_288_), .C(_293_), .Y(_24__3_) );
INVX1 INVX1_53 ( .A(_25_), .Y(_295_) );
NAND2X1 NAND2X1_85 ( .A(_26_), .B(w_cout_4_), .Y(_296_) );
OAI21X1 OAI21X1_85 ( .A(w_cout_4_), .B(_295_), .C(_296_), .Y(csa_inst_cin) );
INVX1 INVX1_54 ( .A(_27__2_), .Y(_297_) );
NAND2X1 NAND2X1_86 ( .A(_28__2_), .B(w_cout_4_), .Y(_298_) );
OAI21X1 OAI21X1_86 ( .A(w_cout_4_), .B(_297_), .C(_298_), .Y(_0__22_) );
INVX1 INVX1_55 ( .A(_27__3_), .Y(_299_) );
NAND2X1 NAND2X1_87 ( .A(w_cout_4_), .B(_28__3_), .Y(_300_) );
OAI21X1 OAI21X1_87 ( .A(w_cout_4_), .B(_299_), .C(_300_), .Y(_0__23_) );
INVX1 INVX1_56 ( .A(_27__0_), .Y(_301_) );
NAND2X1 NAND2X1_88 ( .A(w_cout_4_), .B(_28__0_), .Y(_302_) );
OAI21X1 OAI21X1_88 ( .A(w_cout_4_), .B(_301_), .C(_302_), .Y(_0__20_) );
INVX1 INVX1_57 ( .A(_27__1_), .Y(_303_) );
NAND2X1 NAND2X1_89 ( .A(w_cout_4_), .B(_28__1_), .Y(_304_) );
OAI21X1 OAI21X1_89 ( .A(w_cout_4_), .B(_303_), .C(_304_), .Y(_0__21_) );
INVX1 INVX1_58 ( .A(1'b0), .Y(_308_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_309_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_310_) );
NAND3X1 NAND3X1_33 ( .A(_308_), .B(_310_), .C(_309_), .Y(_311_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_305_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_306_) );
OAI21X1 OAI21X1_90 ( .A(_305_), .B(_306_), .C(1'b0), .Y(_307_) );
NAND2X1 NAND2X1_91 ( .A(_307_), .B(_311_), .Y(_27__0_) );
OAI21X1 OAI21X1_91 ( .A(_308_), .B(_305_), .C(_310_), .Y(_29__1_) );
INVX1 INVX1_59 ( .A(_29__3_), .Y(_315_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_316_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_317_) );
NAND3X1 NAND3X1_34 ( .A(_315_), .B(_317_), .C(_316_), .Y(_318_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_312_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_313_) );
OAI21X1 OAI21X1_92 ( .A(_312_), .B(_313_), .C(_29__3_), .Y(_314_) );
NAND2X1 NAND2X1_93 ( .A(_314_), .B(_318_), .Y(_27__3_) );
OAI21X1 OAI21X1_93 ( .A(_315_), .B(_312_), .C(_317_), .Y(_25_) );
INVX1 INVX1_60 ( .A(_29__1_), .Y(_322_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_323_) );
NAND2X1 NAND2X1_94 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_324_) );
NAND3X1 NAND3X1_35 ( .A(_322_), .B(_324_), .C(_323_), .Y(_325_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_319_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_320_) );
OAI21X1 OAI21X1_94 ( .A(_319_), .B(_320_), .C(_29__1_), .Y(_321_) );
NAND2X1 NAND2X1_95 ( .A(_321_), .B(_325_), .Y(_27__1_) );
OAI21X1 OAI21X1_95 ( .A(_322_), .B(_319_), .C(_324_), .Y(_29__2_) );
INVX1 INVX1_61 ( .A(_29__2_), .Y(_329_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_330_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_331_) );
NAND3X1 NAND3X1_36 ( .A(_329_), .B(_331_), .C(_330_), .Y(_332_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_326_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_327_) );
OAI21X1 OAI21X1_96 ( .A(_326_), .B(_327_), .C(_29__2_), .Y(_328_) );
NAND2X1 NAND2X1_97 ( .A(_328_), .B(_332_), .Y(_27__2_) );
OAI21X1 OAI21X1_97 ( .A(_329_), .B(_326_), .C(_331_), .Y(_29__3_) );
INVX1 INVX1_62 ( .A(1'b1), .Y(_336_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_337_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_338_) );
NAND3X1 NAND3X1_37 ( .A(_336_), .B(_338_), .C(_337_), .Y(_339_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_333_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_334_) );
OAI21X1 OAI21X1_98 ( .A(_333_), .B(_334_), .C(1'b1), .Y(_335_) );
NAND2X1 NAND2X1_99 ( .A(_335_), .B(_339_), .Y(_28__0_) );
OAI21X1 OAI21X1_99 ( .A(_336_), .B(_333_), .C(_338_), .Y(_30__1_) );
INVX1 INVX1_63 ( .A(_30__3_), .Y(_343_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_344_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_345_) );
NAND3X1 NAND3X1_38 ( .A(_343_), .B(_345_), .C(_344_), .Y(_346_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_340_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_341_) );
OAI21X1 OAI21X1_100 ( .A(_340_), .B(_341_), .C(_30__3_), .Y(_342_) );
NAND2X1 NAND2X1_101 ( .A(_342_), .B(_346_), .Y(_28__3_) );
OAI21X1 OAI21X1_101 ( .A(_343_), .B(_340_), .C(_345_), .Y(_26_) );
INVX1 INVX1_64 ( .A(_30__1_), .Y(_350_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_351_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_352_) );
NAND3X1 NAND3X1_39 ( .A(_350_), .B(_352_), .C(_351_), .Y(_353_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_347_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_348_) );
OAI21X1 OAI21X1_102 ( .A(_347_), .B(_348_), .C(_30__1_), .Y(_349_) );
NAND2X1 NAND2X1_103 ( .A(_349_), .B(_353_), .Y(_28__1_) );
OAI21X1 OAI21X1_103 ( .A(_350_), .B(_347_), .C(_352_), .Y(_30__2_) );
INVX1 INVX1_65 ( .A(_30__2_), .Y(_357_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_358_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_359_) );
NAND3X1 NAND3X1_40 ( .A(_357_), .B(_359_), .C(_358_), .Y(_360_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_354_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_355_) );
OAI21X1 OAI21X1_104 ( .A(_354_), .B(_355_), .C(_30__2_), .Y(_356_) );
NAND2X1 NAND2X1_105 ( .A(_356_), .B(_360_), .Y(_28__2_) );
OAI21X1 OAI21X1_105 ( .A(_357_), .B(_354_), .C(_359_), .Y(_30__3_) );
INVX1 INVX1_66 ( .A(csa_inst_cout0_0), .Y(_361_) );
NAND2X1 NAND2X1_106 ( .A(csa_inst_cout0_1), .B(csa_inst_cin), .Y(_362_) );
OAI21X1 OAI21X1_106 ( .A(csa_inst_cin), .B(_361_), .C(_362_), .Y(w_cout_6_) );
INVX1 INVX1_67 ( .A(csa_inst_mux0_sum_i0), .Y(_363_) );
NAND2X1 NAND2X1_107 ( .A(csa_inst_mux0_sum_i1), .B(csa_inst_cin), .Y(_364_) );
OAI21X1 OAI21X1_107 ( .A(csa_inst_cin), .B(_363_), .C(_364_), .Y(csa_inst_mux0_sum_y) );
INVX1 INVX1_68 ( .A(1'b0), .Y(_368_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_369_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_370_) );
NAND3X1 NAND3X1_41 ( .A(_368_), .B(_370_), .C(_369_), .Y(_371_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_365_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_366_) );
OAI21X1 OAI21X1_108 ( .A(_365_), .B(_366_), .C(1'b0), .Y(_367_) );
NAND2X1 NAND2X1_109 ( .A(_367_), .B(_371_), .Y(csa_inst_mux0_sum_i0) );
OAI21X1 OAI21X1_109 ( .A(_368_), .B(_365_), .C(_370_), .Y(csa_inst_cout0_0) );
INVX1 INVX1_69 ( .A(1'b1), .Y(_375_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_376_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_377_) );
NAND3X1 NAND3X1_42 ( .A(_375_), .B(_377_), .C(_376_), .Y(_378_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_372_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_373_) );
OAI21X1 OAI21X1_110 ( .A(_372_), .B(_373_), .C(1'b1), .Y(_374_) );
NAND2X1 NAND2X1_111 ( .A(_374_), .B(_378_), .Y(csa_inst_mux0_sum_i1) );
OAI21X1 OAI21X1_111 ( .A(_375_), .B(_372_), .C(_377_), .Y(csa_inst_cout0_1) );
INVX1 INVX1_70 ( .A(1'b0), .Y(_382_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_383_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_384_) );
NAND3X1 NAND3X1_43 ( .A(_382_), .B(_384_), .C(_383_), .Y(_385_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_379_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_380_) );
OAI21X1 OAI21X1_112 ( .A(_379_), .B(_380_), .C(1'b0), .Y(_381_) );
NAND2X1 NAND2X1_113 ( .A(_381_), .B(_385_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_113 ( .A(_382_), .B(_379_), .C(_384_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_71 ( .A(rca_inst_fa3_i_carry), .Y(_389_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_390_) );
NAND2X1 NAND2X1_114 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_391_) );
NAND3X1 NAND3X1_44 ( .A(_389_), .B(_391_), .C(_390_), .Y(_392_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_386_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_387_) );
OAI21X1 OAI21X1_114 ( .A(_386_), .B(_387_), .C(rca_inst_fa3_i_carry), .Y(_388_) );
NAND2X1 NAND2X1_115 ( .A(_388_), .B(_392_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_115 ( .A(_389_), .B(_386_), .C(_391_), .Y(rca_inst_cout) );
INVX1 INVX1_72 ( .A(rca_inst_fa0_o_carry), .Y(_396_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_397_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_398_) );
NAND3X1 NAND3X1_45 ( .A(_396_), .B(_398_), .C(_397_), .Y(_399_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_393_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_394_) );
OAI21X1 OAI21X1_116 ( .A(_393_), .B(_394_), .C(rca_inst_fa0_o_carry), .Y(_395_) );
NAND2X1 NAND2X1_117 ( .A(_395_), .B(_399_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_117 ( .A(_396_), .B(_393_), .C(_398_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_73 ( .A(rca_inst_fa_1__o_carry), .Y(_403_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_404_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_405_) );
NAND3X1 NAND3X1_46 ( .A(_403_), .B(_405_), .C(_404_), .Y(_406_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_400_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_401_) );
OAI21X1 OAI21X1_118 ( .A(_400_), .B(_401_), .C(rca_inst_fa_1__o_carry), .Y(_402_) );
NAND2X1 NAND2X1_119 ( .A(_402_), .B(_406_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_119 ( .A(_403_), .B(_400_), .C(_405_), .Y(rca_inst_fa3_i_carry) );
BUFX2 BUFX2_27 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_28 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_29 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_30 ( .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_31 ( .A(csa_inst_mux0_sum_y), .Y(_0__24_) );
BUFX2 BUFX2_32 ( .A(rca_inst_cout), .Y(w_cout_0_) );
BUFX2 BUFX2_33 ( .A(csa_inst_cin), .Y(w_cout_5_) );
endmodule
