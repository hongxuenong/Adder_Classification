module csa_38bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output cout;

OR2X2 OR2X2_1 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_275_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_276_) );
NAND3X1 NAND3X1_1 ( .A(_274_), .B(_276_), .C(_275_), .Y(_277_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_271_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_272_) );
OAI21X1 OAI21X1_1 ( .A(_271_), .B(_272_), .C(_17__2_), .Y(_273_) );
NAND2X1 NAND2X1_2 ( .A(_273_), .B(_277_), .Y(_15__2_) );
OAI21X1 OAI21X1_2 ( .A(_274_), .B(_271_), .C(_276_), .Y(_17__3_) );
INVX1 INVX1_1 ( .A(_17__3_), .Y(_281_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_282_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_283_) );
NAND3X1 NAND3X1_2 ( .A(_281_), .B(_283_), .C(_282_), .Y(_284_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_278_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_279_) );
OAI21X1 OAI21X1_3 ( .A(_278_), .B(_279_), .C(_17__3_), .Y(_280_) );
NAND2X1 NAND2X1_4 ( .A(_280_), .B(_284_), .Y(_15__3_) );
OAI21X1 OAI21X1_4 ( .A(_281_), .B(_278_), .C(_283_), .Y(_13_) );
INVX1 INVX1_2 ( .A(1'b1), .Y(_288_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_289_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_290_) );
NAND3X1 NAND3X1_3 ( .A(_288_), .B(_290_), .C(_289_), .Y(_291_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_285_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_286_) );
OAI21X1 OAI21X1_5 ( .A(_285_), .B(_286_), .C(1'b1), .Y(_287_) );
NAND2X1 NAND2X1_6 ( .A(_287_), .B(_291_), .Y(_16__0_) );
OAI21X1 OAI21X1_6 ( .A(_288_), .B(_285_), .C(_290_), .Y(_18__1_) );
INVX1 INVX1_3 ( .A(_18__1_), .Y(_295_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_296_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_297_) );
NAND3X1 NAND3X1_4 ( .A(_295_), .B(_297_), .C(_296_), .Y(_298_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_292_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_293_) );
OAI21X1 OAI21X1_7 ( .A(_292_), .B(_293_), .C(_18__1_), .Y(_294_) );
NAND2X1 NAND2X1_8 ( .A(_294_), .B(_298_), .Y(_16__1_) );
OAI21X1 OAI21X1_8 ( .A(_295_), .B(_292_), .C(_297_), .Y(_18__2_) );
INVX1 INVX1_4 ( .A(_18__2_), .Y(_302_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_303_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_304_) );
NAND3X1 NAND3X1_5 ( .A(_302_), .B(_304_), .C(_303_), .Y(_305_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_299_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_300_) );
OAI21X1 OAI21X1_9 ( .A(_299_), .B(_300_), .C(_18__2_), .Y(_301_) );
NAND2X1 NAND2X1_10 ( .A(_301_), .B(_305_), .Y(_16__2_) );
OAI21X1 OAI21X1_10 ( .A(_302_), .B(_299_), .C(_304_), .Y(_18__3_) );
INVX1 INVX1_5 ( .A(_18__3_), .Y(_309_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_310_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_311_) );
NAND3X1 NAND3X1_6 ( .A(_309_), .B(_311_), .C(_310_), .Y(_312_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_306_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_307_) );
OAI21X1 OAI21X1_11 ( .A(_306_), .B(_307_), .C(_18__3_), .Y(_308_) );
NAND2X1 NAND2X1_12 ( .A(_308_), .B(_312_), .Y(_16__3_) );
OAI21X1 OAI21X1_12 ( .A(_309_), .B(_306_), .C(_311_), .Y(_14_) );
INVX1 INVX1_6 ( .A(1'b0), .Y(_316_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_317_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_318_) );
NAND3X1 NAND3X1_7 ( .A(_316_), .B(_318_), .C(_317_), .Y(_319_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_313_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_314_) );
OAI21X1 OAI21X1_13 ( .A(_313_), .B(_314_), .C(1'b0), .Y(_315_) );
NAND2X1 NAND2X1_14 ( .A(_315_), .B(_319_), .Y(_21__0_) );
OAI21X1 OAI21X1_14 ( .A(_316_), .B(_313_), .C(_318_), .Y(_23__1_) );
INVX1 INVX1_7 ( .A(_23__1_), .Y(_323_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_324_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_325_) );
NAND3X1 NAND3X1_8 ( .A(_323_), .B(_325_), .C(_324_), .Y(_326_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_320_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_321_) );
OAI21X1 OAI21X1_15 ( .A(_320_), .B(_321_), .C(_23__1_), .Y(_322_) );
NAND2X1 NAND2X1_16 ( .A(_322_), .B(_326_), .Y(_21__1_) );
OAI21X1 OAI21X1_16 ( .A(_323_), .B(_320_), .C(_325_), .Y(_23__2_) );
INVX1 INVX1_8 ( .A(_23__2_), .Y(_330_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_331_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_332_) );
NAND3X1 NAND3X1_9 ( .A(_330_), .B(_332_), .C(_331_), .Y(_333_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_327_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_328_) );
OAI21X1 OAI21X1_17 ( .A(_327_), .B(_328_), .C(_23__2_), .Y(_329_) );
NAND2X1 NAND2X1_18 ( .A(_329_), .B(_333_), .Y(_21__2_) );
OAI21X1 OAI21X1_18 ( .A(_330_), .B(_327_), .C(_332_), .Y(_23__3_) );
INVX1 INVX1_9 ( .A(_23__3_), .Y(_337_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_338_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_339_) );
NAND3X1 NAND3X1_10 ( .A(_337_), .B(_339_), .C(_338_), .Y(_340_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_334_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_335_) );
OAI21X1 OAI21X1_19 ( .A(_334_), .B(_335_), .C(_23__3_), .Y(_336_) );
NAND2X1 NAND2X1_20 ( .A(_336_), .B(_340_), .Y(_21__3_) );
OAI21X1 OAI21X1_20 ( .A(_337_), .B(_334_), .C(_339_), .Y(_19_) );
INVX1 INVX1_10 ( .A(1'b1), .Y(_344_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_345_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_346_) );
NAND3X1 NAND3X1_11 ( .A(_344_), .B(_346_), .C(_345_), .Y(_347_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_341_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_342_) );
OAI21X1 OAI21X1_21 ( .A(_341_), .B(_342_), .C(1'b1), .Y(_343_) );
NAND2X1 NAND2X1_22 ( .A(_343_), .B(_347_), .Y(_22__0_) );
OAI21X1 OAI21X1_22 ( .A(_344_), .B(_341_), .C(_346_), .Y(_24__1_) );
INVX1 INVX1_11 ( .A(_24__1_), .Y(_351_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_352_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_353_) );
NAND3X1 NAND3X1_12 ( .A(_351_), .B(_353_), .C(_352_), .Y(_354_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_348_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_349_) );
OAI21X1 OAI21X1_23 ( .A(_348_), .B(_349_), .C(_24__1_), .Y(_350_) );
NAND2X1 NAND2X1_24 ( .A(_350_), .B(_354_), .Y(_22__1_) );
OAI21X1 OAI21X1_24 ( .A(_351_), .B(_348_), .C(_353_), .Y(_24__2_) );
INVX1 INVX1_12 ( .A(_24__2_), .Y(_358_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_359_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_360_) );
NAND3X1 NAND3X1_13 ( .A(_358_), .B(_360_), .C(_359_), .Y(_361_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_355_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_356_) );
OAI21X1 OAI21X1_25 ( .A(_355_), .B(_356_), .C(_24__2_), .Y(_357_) );
NAND2X1 NAND2X1_26 ( .A(_357_), .B(_361_), .Y(_22__2_) );
OAI21X1 OAI21X1_26 ( .A(_358_), .B(_355_), .C(_360_), .Y(_24__3_) );
INVX1 INVX1_13 ( .A(_24__3_), .Y(_365_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_366_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_367_) );
NAND3X1 NAND3X1_14 ( .A(_365_), .B(_367_), .C(_366_), .Y(_368_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_362_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_363_) );
OAI21X1 OAI21X1_27 ( .A(_362_), .B(_363_), .C(_24__3_), .Y(_364_) );
NAND2X1 NAND2X1_28 ( .A(_364_), .B(_368_), .Y(_22__3_) );
OAI21X1 OAI21X1_28 ( .A(_365_), .B(_362_), .C(_367_), .Y(_20_) );
INVX1 INVX1_14 ( .A(1'b0), .Y(_372_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_373_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_374_) );
NAND3X1 NAND3X1_15 ( .A(_372_), .B(_374_), .C(_373_), .Y(_375_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_369_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_370_) );
OAI21X1 OAI21X1_29 ( .A(_369_), .B(_370_), .C(1'b0), .Y(_371_) );
NAND2X1 NAND2X1_30 ( .A(_371_), .B(_375_), .Y(_27__0_) );
OAI21X1 OAI21X1_30 ( .A(_372_), .B(_369_), .C(_374_), .Y(_29__1_) );
INVX1 INVX1_15 ( .A(_29__1_), .Y(_379_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_380_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_381_) );
NAND3X1 NAND3X1_16 ( .A(_379_), .B(_381_), .C(_380_), .Y(_382_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_376_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_377_) );
OAI21X1 OAI21X1_31 ( .A(_376_), .B(_377_), .C(_29__1_), .Y(_378_) );
NAND2X1 NAND2X1_32 ( .A(_378_), .B(_382_), .Y(_27__1_) );
OAI21X1 OAI21X1_32 ( .A(_379_), .B(_376_), .C(_381_), .Y(_29__2_) );
INVX1 INVX1_16 ( .A(_29__2_), .Y(_386_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_387_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_388_) );
NAND3X1 NAND3X1_17 ( .A(_386_), .B(_388_), .C(_387_), .Y(_389_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_383_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_384_) );
OAI21X1 OAI21X1_33 ( .A(_383_), .B(_384_), .C(_29__2_), .Y(_385_) );
NAND2X1 NAND2X1_34 ( .A(_385_), .B(_389_), .Y(_27__2_) );
OAI21X1 OAI21X1_34 ( .A(_386_), .B(_383_), .C(_388_), .Y(_29__3_) );
INVX1 INVX1_17 ( .A(_29__3_), .Y(_393_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_394_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_395_) );
NAND3X1 NAND3X1_18 ( .A(_393_), .B(_395_), .C(_394_), .Y(_396_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_390_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_391_) );
OAI21X1 OAI21X1_35 ( .A(_390_), .B(_391_), .C(_29__3_), .Y(_392_) );
NAND2X1 NAND2X1_36 ( .A(_392_), .B(_396_), .Y(_27__3_) );
OAI21X1 OAI21X1_36 ( .A(_393_), .B(_390_), .C(_395_), .Y(_25_) );
INVX1 INVX1_18 ( .A(1'b1), .Y(_400_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_401_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_402_) );
NAND3X1 NAND3X1_19 ( .A(_400_), .B(_402_), .C(_401_), .Y(_403_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_397_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_398_) );
OAI21X1 OAI21X1_37 ( .A(_397_), .B(_398_), .C(1'b1), .Y(_399_) );
NAND2X1 NAND2X1_38 ( .A(_399_), .B(_403_), .Y(_28__0_) );
OAI21X1 OAI21X1_38 ( .A(_400_), .B(_397_), .C(_402_), .Y(_30__1_) );
INVX1 INVX1_19 ( .A(_30__1_), .Y(_407_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_408_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_409_) );
NAND3X1 NAND3X1_20 ( .A(_407_), .B(_409_), .C(_408_), .Y(_410_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_404_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_405_) );
OAI21X1 OAI21X1_39 ( .A(_404_), .B(_405_), .C(_30__1_), .Y(_406_) );
NAND2X1 NAND2X1_40 ( .A(_406_), .B(_410_), .Y(_28__1_) );
OAI21X1 OAI21X1_40 ( .A(_407_), .B(_404_), .C(_409_), .Y(_30__2_) );
INVX1 INVX1_20 ( .A(_30__2_), .Y(_414_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_415_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_416_) );
NAND3X1 NAND3X1_21 ( .A(_414_), .B(_416_), .C(_415_), .Y(_417_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_411_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_412_) );
OAI21X1 OAI21X1_41 ( .A(_411_), .B(_412_), .C(_30__2_), .Y(_413_) );
NAND2X1 NAND2X1_42 ( .A(_413_), .B(_417_), .Y(_28__2_) );
OAI21X1 OAI21X1_42 ( .A(_414_), .B(_411_), .C(_416_), .Y(_30__3_) );
INVX1 INVX1_21 ( .A(_30__3_), .Y(_421_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_422_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_423_) );
NAND3X1 NAND3X1_22 ( .A(_421_), .B(_423_), .C(_422_), .Y(_424_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_418_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_419_) );
OAI21X1 OAI21X1_43 ( .A(_418_), .B(_419_), .C(_30__3_), .Y(_420_) );
NAND2X1 NAND2X1_44 ( .A(_420_), .B(_424_), .Y(_28__3_) );
OAI21X1 OAI21X1_44 ( .A(_421_), .B(_418_), .C(_423_), .Y(_26_) );
INVX1 INVX1_22 ( .A(1'b0), .Y(_428_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_429_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_430_) );
NAND3X1 NAND3X1_23 ( .A(_428_), .B(_430_), .C(_429_), .Y(_431_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_425_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_426_) );
OAI21X1 OAI21X1_45 ( .A(_425_), .B(_426_), .C(1'b0), .Y(_427_) );
NAND2X1 NAND2X1_46 ( .A(_427_), .B(_431_), .Y(_33__0_) );
OAI21X1 OAI21X1_46 ( .A(_428_), .B(_425_), .C(_430_), .Y(_35__1_) );
INVX1 INVX1_23 ( .A(_35__1_), .Y(_435_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_436_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_437_) );
NAND3X1 NAND3X1_24 ( .A(_435_), .B(_437_), .C(_436_), .Y(_438_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_432_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_433_) );
OAI21X1 OAI21X1_47 ( .A(_432_), .B(_433_), .C(_35__1_), .Y(_434_) );
NAND2X1 NAND2X1_48 ( .A(_434_), .B(_438_), .Y(_33__1_) );
OAI21X1 OAI21X1_48 ( .A(_435_), .B(_432_), .C(_437_), .Y(_35__2_) );
INVX1 INVX1_24 ( .A(_35__2_), .Y(_442_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_443_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_444_) );
NAND3X1 NAND3X1_25 ( .A(_442_), .B(_444_), .C(_443_), .Y(_445_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_439_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_440_) );
OAI21X1 OAI21X1_49 ( .A(_439_), .B(_440_), .C(_35__2_), .Y(_441_) );
NAND2X1 NAND2X1_50 ( .A(_441_), .B(_445_), .Y(_33__2_) );
OAI21X1 OAI21X1_50 ( .A(_442_), .B(_439_), .C(_444_), .Y(_35__3_) );
INVX1 INVX1_25 ( .A(_35__3_), .Y(_449_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_450_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_451_) );
NAND3X1 NAND3X1_26 ( .A(_449_), .B(_451_), .C(_450_), .Y(_452_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_446_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_447_) );
OAI21X1 OAI21X1_51 ( .A(_446_), .B(_447_), .C(_35__3_), .Y(_448_) );
NAND2X1 NAND2X1_52 ( .A(_448_), .B(_452_), .Y(_33__3_) );
OAI21X1 OAI21X1_52 ( .A(_449_), .B(_446_), .C(_451_), .Y(_31_) );
INVX1 INVX1_26 ( .A(1'b1), .Y(_456_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_457_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_458_) );
NAND3X1 NAND3X1_27 ( .A(_456_), .B(_458_), .C(_457_), .Y(_459_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_453_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_454_) );
OAI21X1 OAI21X1_53 ( .A(_453_), .B(_454_), .C(1'b1), .Y(_455_) );
NAND2X1 NAND2X1_54 ( .A(_455_), .B(_459_), .Y(_34__0_) );
OAI21X1 OAI21X1_54 ( .A(_456_), .B(_453_), .C(_458_), .Y(_36__1_) );
INVX1 INVX1_27 ( .A(_36__1_), .Y(_463_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_464_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_465_) );
NAND3X1 NAND3X1_28 ( .A(_463_), .B(_465_), .C(_464_), .Y(_466_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_460_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_461_) );
OAI21X1 OAI21X1_55 ( .A(_460_), .B(_461_), .C(_36__1_), .Y(_462_) );
NAND2X1 NAND2X1_56 ( .A(_462_), .B(_466_), .Y(_34__1_) );
OAI21X1 OAI21X1_56 ( .A(_463_), .B(_460_), .C(_465_), .Y(_36__2_) );
INVX1 INVX1_28 ( .A(_36__2_), .Y(_470_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_471_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_472_) );
NAND3X1 NAND3X1_29 ( .A(_470_), .B(_472_), .C(_471_), .Y(_473_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_467_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_468_) );
OAI21X1 OAI21X1_57 ( .A(_467_), .B(_468_), .C(_36__2_), .Y(_469_) );
NAND2X1 NAND2X1_58 ( .A(_469_), .B(_473_), .Y(_34__2_) );
OAI21X1 OAI21X1_58 ( .A(_470_), .B(_467_), .C(_472_), .Y(_36__3_) );
INVX1 INVX1_29 ( .A(_36__3_), .Y(_477_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_478_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_479_) );
NAND3X1 NAND3X1_30 ( .A(_477_), .B(_479_), .C(_478_), .Y(_480_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_474_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_475_) );
OAI21X1 OAI21X1_59 ( .A(_474_), .B(_475_), .C(_36__3_), .Y(_476_) );
NAND2X1 NAND2X1_60 ( .A(_476_), .B(_480_), .Y(_34__3_) );
OAI21X1 OAI21X1_60 ( .A(_477_), .B(_474_), .C(_479_), .Y(_32_) );
INVX1 INVX1_30 ( .A(1'b0), .Y(_484_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_485_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_486_) );
NAND3X1 NAND3X1_31 ( .A(_484_), .B(_486_), .C(_485_), .Y(_487_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_481_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_482_) );
OAI21X1 OAI21X1_61 ( .A(_481_), .B(_482_), .C(1'b0), .Y(_483_) );
NAND2X1 NAND2X1_62 ( .A(_483_), .B(_487_), .Y(_39__0_) );
OAI21X1 OAI21X1_62 ( .A(_484_), .B(_481_), .C(_486_), .Y(_41__1_) );
INVX1 INVX1_31 ( .A(_41__1_), .Y(_491_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_492_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_493_) );
NAND3X1 NAND3X1_32 ( .A(_491_), .B(_493_), .C(_492_), .Y(_494_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_488_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_489_) );
OAI21X1 OAI21X1_63 ( .A(_488_), .B(_489_), .C(_41__1_), .Y(_490_) );
NAND2X1 NAND2X1_64 ( .A(_490_), .B(_494_), .Y(_39__1_) );
OAI21X1 OAI21X1_64 ( .A(_491_), .B(_488_), .C(_493_), .Y(_41__2_) );
INVX1 INVX1_32 ( .A(_41__2_), .Y(_498_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_499_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_500_) );
NAND3X1 NAND3X1_33 ( .A(_498_), .B(_500_), .C(_499_), .Y(_501_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_495_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_496_) );
OAI21X1 OAI21X1_65 ( .A(_495_), .B(_496_), .C(_41__2_), .Y(_497_) );
NAND2X1 NAND2X1_66 ( .A(_497_), .B(_501_), .Y(_39__2_) );
OAI21X1 OAI21X1_66 ( .A(_498_), .B(_495_), .C(_500_), .Y(_41__3_) );
INVX1 INVX1_33 ( .A(_41__3_), .Y(_505_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_506_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_507_) );
NAND3X1 NAND3X1_34 ( .A(_505_), .B(_507_), .C(_506_), .Y(_508_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_502_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_503_) );
OAI21X1 OAI21X1_67 ( .A(_502_), .B(_503_), .C(_41__3_), .Y(_504_) );
NAND2X1 NAND2X1_68 ( .A(_504_), .B(_508_), .Y(_39__3_) );
OAI21X1 OAI21X1_68 ( .A(_505_), .B(_502_), .C(_507_), .Y(_37_) );
INVX1 INVX1_34 ( .A(1'b1), .Y(_512_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_513_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_514_) );
NAND3X1 NAND3X1_35 ( .A(_512_), .B(_514_), .C(_513_), .Y(_515_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_509_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_510_) );
OAI21X1 OAI21X1_69 ( .A(_509_), .B(_510_), .C(1'b1), .Y(_511_) );
NAND2X1 NAND2X1_70 ( .A(_511_), .B(_515_), .Y(_40__0_) );
OAI21X1 OAI21X1_70 ( .A(_512_), .B(_509_), .C(_514_), .Y(_42__1_) );
INVX1 INVX1_35 ( .A(_42__1_), .Y(_519_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_520_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_521_) );
NAND3X1 NAND3X1_36 ( .A(_519_), .B(_521_), .C(_520_), .Y(_522_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_516_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_517_) );
OAI21X1 OAI21X1_71 ( .A(_516_), .B(_517_), .C(_42__1_), .Y(_518_) );
NAND2X1 NAND2X1_72 ( .A(_518_), .B(_522_), .Y(_40__1_) );
OAI21X1 OAI21X1_72 ( .A(_519_), .B(_516_), .C(_521_), .Y(_42__2_) );
INVX1 INVX1_36 ( .A(_42__2_), .Y(_526_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_527_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_528_) );
NAND3X1 NAND3X1_37 ( .A(_526_), .B(_528_), .C(_527_), .Y(_529_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_523_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_524_) );
OAI21X1 OAI21X1_73 ( .A(_523_), .B(_524_), .C(_42__2_), .Y(_525_) );
NAND2X1 NAND2X1_74 ( .A(_525_), .B(_529_), .Y(_40__2_) );
OAI21X1 OAI21X1_74 ( .A(_526_), .B(_523_), .C(_528_), .Y(_42__3_) );
INVX1 INVX1_37 ( .A(_42__3_), .Y(_533_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_534_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_535_) );
NAND3X1 NAND3X1_38 ( .A(_533_), .B(_535_), .C(_534_), .Y(_536_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_530_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_531_) );
OAI21X1 OAI21X1_75 ( .A(_530_), .B(_531_), .C(_42__3_), .Y(_532_) );
NAND2X1 NAND2X1_76 ( .A(_532_), .B(_536_), .Y(_40__3_) );
OAI21X1 OAI21X1_76 ( .A(_533_), .B(_530_), .C(_535_), .Y(_38_) );
INVX1 INVX1_38 ( .A(1'b0), .Y(_540_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_541_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_542_) );
NAND3X1 NAND3X1_39 ( .A(_540_), .B(_542_), .C(_541_), .Y(_543_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_537_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_538_) );
OAI21X1 OAI21X1_77 ( .A(_537_), .B(_538_), .C(1'b0), .Y(_539_) );
NAND2X1 NAND2X1_78 ( .A(_539_), .B(_543_), .Y(_45__0_) );
OAI21X1 OAI21X1_78 ( .A(_540_), .B(_537_), .C(_542_), .Y(_47__1_) );
INVX1 INVX1_39 ( .A(_47__1_), .Y(_547_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_548_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_549_) );
NAND3X1 NAND3X1_40 ( .A(_547_), .B(_549_), .C(_548_), .Y(_550_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_544_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_545_) );
OAI21X1 OAI21X1_79 ( .A(_544_), .B(_545_), .C(_47__1_), .Y(_546_) );
NAND2X1 NAND2X1_80 ( .A(_546_), .B(_550_), .Y(_45__1_) );
OAI21X1 OAI21X1_80 ( .A(_547_), .B(_544_), .C(_549_), .Y(_47__2_) );
INVX1 INVX1_40 ( .A(_47__2_), .Y(_554_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_555_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_556_) );
NAND3X1 NAND3X1_41 ( .A(_554_), .B(_556_), .C(_555_), .Y(_557_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_551_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_552_) );
OAI21X1 OAI21X1_81 ( .A(_551_), .B(_552_), .C(_47__2_), .Y(_553_) );
NAND2X1 NAND2X1_82 ( .A(_553_), .B(_557_), .Y(_45__2_) );
OAI21X1 OAI21X1_82 ( .A(_554_), .B(_551_), .C(_556_), .Y(_47__3_) );
INVX1 INVX1_41 ( .A(_47__3_), .Y(_561_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_562_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_563_) );
NAND3X1 NAND3X1_42 ( .A(_561_), .B(_563_), .C(_562_), .Y(_564_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_558_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_559_) );
OAI21X1 OAI21X1_83 ( .A(_558_), .B(_559_), .C(_47__3_), .Y(_560_) );
NAND2X1 NAND2X1_84 ( .A(_560_), .B(_564_), .Y(_45__3_) );
OAI21X1 OAI21X1_84 ( .A(_561_), .B(_558_), .C(_563_), .Y(_43_) );
INVX1 INVX1_42 ( .A(1'b1), .Y(_568_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_569_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_570_) );
NAND3X1 NAND3X1_43 ( .A(_568_), .B(_570_), .C(_569_), .Y(_571_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_565_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_566_) );
OAI21X1 OAI21X1_85 ( .A(_565_), .B(_566_), .C(1'b1), .Y(_567_) );
NAND2X1 NAND2X1_86 ( .A(_567_), .B(_571_), .Y(_46__0_) );
OAI21X1 OAI21X1_86 ( .A(_568_), .B(_565_), .C(_570_), .Y(_48__1_) );
INVX1 INVX1_43 ( .A(_48__1_), .Y(_575_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_576_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_577_) );
NAND3X1 NAND3X1_44 ( .A(_575_), .B(_577_), .C(_576_), .Y(_578_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_572_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_573_) );
OAI21X1 OAI21X1_87 ( .A(_572_), .B(_573_), .C(_48__1_), .Y(_574_) );
NAND2X1 NAND2X1_88 ( .A(_574_), .B(_578_), .Y(_46__1_) );
OAI21X1 OAI21X1_88 ( .A(_575_), .B(_572_), .C(_577_), .Y(_48__2_) );
INVX1 INVX1_44 ( .A(_48__2_), .Y(_582_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_583_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_584_) );
NAND3X1 NAND3X1_45 ( .A(_582_), .B(_584_), .C(_583_), .Y(_585_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_579_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_580_) );
OAI21X1 OAI21X1_89 ( .A(_579_), .B(_580_), .C(_48__2_), .Y(_581_) );
NAND2X1 NAND2X1_90 ( .A(_581_), .B(_585_), .Y(_46__2_) );
OAI21X1 OAI21X1_90 ( .A(_582_), .B(_579_), .C(_584_), .Y(_48__3_) );
INVX1 INVX1_45 ( .A(_48__3_), .Y(_589_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_590_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_591_) );
NAND3X1 NAND3X1_46 ( .A(_589_), .B(_591_), .C(_590_), .Y(_592_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_586_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_587_) );
OAI21X1 OAI21X1_91 ( .A(_586_), .B(_587_), .C(_48__3_), .Y(_588_) );
NAND2X1 NAND2X1_92 ( .A(_588_), .B(_592_), .Y(_46__3_) );
OAI21X1 OAI21X1_92 ( .A(_589_), .B(_586_), .C(_591_), .Y(_44_) );
INVX1 INVX1_46 ( .A(1'b0), .Y(_596_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_597_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_598_) );
NAND3X1 NAND3X1_47 ( .A(_596_), .B(_598_), .C(_597_), .Y(_599_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_593_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_594_) );
OAI21X1 OAI21X1_93 ( .A(_593_), .B(_594_), .C(1'b0), .Y(_595_) );
NAND2X1 NAND2X1_94 ( .A(_595_), .B(_599_), .Y(_51__0_) );
OAI21X1 OAI21X1_94 ( .A(_596_), .B(_593_), .C(_598_), .Y(_53__1_) );
INVX1 INVX1_47 ( .A(_53__1_), .Y(_603_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_604_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_605_) );
NAND3X1 NAND3X1_48 ( .A(_603_), .B(_605_), .C(_604_), .Y(_606_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_600_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_601_) );
OAI21X1 OAI21X1_95 ( .A(_600_), .B(_601_), .C(_53__1_), .Y(_602_) );
NAND2X1 NAND2X1_96 ( .A(_602_), .B(_606_), .Y(_51__1_) );
OAI21X1 OAI21X1_96 ( .A(_603_), .B(_600_), .C(_605_), .Y(_53__2_) );
INVX1 INVX1_48 ( .A(_53__2_), .Y(_610_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_611_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_612_) );
NAND3X1 NAND3X1_49 ( .A(_610_), .B(_612_), .C(_611_), .Y(_613_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_607_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_608_) );
OAI21X1 OAI21X1_97 ( .A(_607_), .B(_608_), .C(_53__2_), .Y(_609_) );
NAND2X1 NAND2X1_98 ( .A(_609_), .B(_613_), .Y(_51__2_) );
OAI21X1 OAI21X1_98 ( .A(_610_), .B(_607_), .C(_612_), .Y(_53__3_) );
INVX1 INVX1_49 ( .A(_53__3_), .Y(_617_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_618_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_619_) );
NAND3X1 NAND3X1_50 ( .A(_617_), .B(_619_), .C(_618_), .Y(_620_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_614_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_615_) );
OAI21X1 OAI21X1_99 ( .A(_614_), .B(_615_), .C(_53__3_), .Y(_616_) );
NAND2X1 NAND2X1_100 ( .A(_616_), .B(_620_), .Y(_51__3_) );
OAI21X1 OAI21X1_100 ( .A(_617_), .B(_614_), .C(_619_), .Y(_49_) );
INVX1 INVX1_50 ( .A(1'b1), .Y(_624_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_625_) );
NAND2X1 NAND2X1_101 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_626_) );
NAND3X1 NAND3X1_51 ( .A(_624_), .B(_626_), .C(_625_), .Y(_627_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_621_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_622_) );
OAI21X1 OAI21X1_101 ( .A(_621_), .B(_622_), .C(1'b1), .Y(_623_) );
NAND2X1 NAND2X1_102 ( .A(_623_), .B(_627_), .Y(_52__0_) );
OAI21X1 OAI21X1_102 ( .A(_624_), .B(_621_), .C(_626_), .Y(_54__1_) );
INVX1 INVX1_51 ( .A(_54__1_), .Y(_631_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_632_) );
NAND2X1 NAND2X1_103 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_633_) );
NAND3X1 NAND3X1_52 ( .A(_631_), .B(_633_), .C(_632_), .Y(_634_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_628_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_629_) );
OAI21X1 OAI21X1_103 ( .A(_628_), .B(_629_), .C(_54__1_), .Y(_630_) );
NAND2X1 NAND2X1_104 ( .A(_630_), .B(_634_), .Y(_52__1_) );
OAI21X1 OAI21X1_104 ( .A(_631_), .B(_628_), .C(_633_), .Y(_54__2_) );
INVX1 INVX1_52 ( .A(_54__2_), .Y(_638_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_639_) );
NAND2X1 NAND2X1_105 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_640_) );
NAND3X1 NAND3X1_53 ( .A(_638_), .B(_640_), .C(_639_), .Y(_641_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_635_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_636_) );
OAI21X1 OAI21X1_105 ( .A(_635_), .B(_636_), .C(_54__2_), .Y(_637_) );
NAND2X1 NAND2X1_106 ( .A(_637_), .B(_641_), .Y(_52__2_) );
OAI21X1 OAI21X1_106 ( .A(_638_), .B(_635_), .C(_640_), .Y(_54__3_) );
INVX1 INVX1_53 ( .A(_54__3_), .Y(_645_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_646_) );
NAND2X1 NAND2X1_107 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_647_) );
NAND3X1 NAND3X1_54 ( .A(_645_), .B(_647_), .C(_646_), .Y(_648_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_642_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_643_) );
OAI21X1 OAI21X1_107 ( .A(_642_), .B(_643_), .C(_54__3_), .Y(_644_) );
NAND2X1 NAND2X1_108 ( .A(_644_), .B(_648_), .Y(_52__3_) );
OAI21X1 OAI21X1_108 ( .A(_645_), .B(_642_), .C(_647_), .Y(_50_) );
INVX1 INVX1_54 ( .A(1'b0), .Y(_652_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_653_) );
NAND2X1 NAND2X1_109 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_654_) );
NAND3X1 NAND3X1_55 ( .A(_652_), .B(_654_), .C(_653_), .Y(_655_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_649_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_650_) );
OAI21X1 OAI21X1_109 ( .A(_649_), .B(_650_), .C(1'b0), .Y(_651_) );
NAND2X1 NAND2X1_110 ( .A(_651_), .B(_655_), .Y(_0__0_) );
OAI21X1 OAI21X1_110 ( .A(_652_), .B(_649_), .C(_654_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_55 ( .A(rca_inst_w_CARRY_1_), .Y(_659_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_660_) );
NAND2X1 NAND2X1_111 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_661_) );
NAND3X1 NAND3X1_56 ( .A(_659_), .B(_661_), .C(_660_), .Y(_662_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_656_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_657_) );
OAI21X1 OAI21X1_111 ( .A(_656_), .B(_657_), .C(rca_inst_w_CARRY_1_), .Y(_658_) );
NAND2X1 NAND2X1_112 ( .A(_658_), .B(_662_), .Y(_0__1_) );
BUFX2 BUFX2_1 ( .A(w_cout_9_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
INVX1 INVX1_56 ( .A(_1_), .Y(_55_) );
NAND2X1 NAND2X1_113 ( .A(_2_), .B(1'b0), .Y(_56_) );
OAI21X1 OAI21X1_112 ( .A(1'b0), .B(_55_), .C(_56_), .Y(w_cout_1_) );
INVX1 INVX1_57 ( .A(_3__0_), .Y(_57_) );
NAND2X1 NAND2X1_114 ( .A(_4__0_), .B(1'b0), .Y(_58_) );
OAI21X1 OAI21X1_113 ( .A(1'b0), .B(_57_), .C(_58_), .Y(_0__2_) );
INVX1 INVX1_58 ( .A(_3__1_), .Y(_59_) );
NAND2X1 NAND2X1_115 ( .A(1'b0), .B(_4__1_), .Y(_60_) );
OAI21X1 OAI21X1_114 ( .A(1'b0), .B(_59_), .C(_60_), .Y(_0__3_) );
INVX1 INVX1_59 ( .A(_3__2_), .Y(_61_) );
NAND2X1 NAND2X1_116 ( .A(1'b0), .B(_4__2_), .Y(_62_) );
OAI21X1 OAI21X1_115 ( .A(1'b0), .B(_61_), .C(_62_), .Y(_0__4_) );
INVX1 INVX1_60 ( .A(_3__3_), .Y(_63_) );
NAND2X1 NAND2X1_117 ( .A(1'b0), .B(_4__3_), .Y(_64_) );
OAI21X1 OAI21X1_116 ( .A(1'b0), .B(_63_), .C(_64_), .Y(_0__5_) );
INVX1 INVX1_61 ( .A(_7_), .Y(_65_) );
NAND2X1 NAND2X1_118 ( .A(_8_), .B(w_cout_1_), .Y(_66_) );
OAI21X1 OAI21X1_117 ( .A(w_cout_1_), .B(_65_), .C(_66_), .Y(w_cout_2_) );
INVX1 INVX1_62 ( .A(_9__0_), .Y(_67_) );
NAND2X1 NAND2X1_119 ( .A(_10__0_), .B(w_cout_1_), .Y(_68_) );
OAI21X1 OAI21X1_118 ( .A(w_cout_1_), .B(_67_), .C(_68_), .Y(_0__6_) );
INVX1 INVX1_63 ( .A(_9__1_), .Y(_69_) );
NAND2X1 NAND2X1_120 ( .A(w_cout_1_), .B(_10__1_), .Y(_70_) );
OAI21X1 OAI21X1_119 ( .A(w_cout_1_), .B(_69_), .C(_70_), .Y(_0__7_) );
INVX1 INVX1_64 ( .A(_9__2_), .Y(_71_) );
NAND2X1 NAND2X1_121 ( .A(w_cout_1_), .B(_10__2_), .Y(_72_) );
OAI21X1 OAI21X1_120 ( .A(w_cout_1_), .B(_71_), .C(_72_), .Y(_0__8_) );
INVX1 INVX1_65 ( .A(_9__3_), .Y(_73_) );
NAND2X1 NAND2X1_122 ( .A(w_cout_1_), .B(_10__3_), .Y(_74_) );
OAI21X1 OAI21X1_121 ( .A(w_cout_1_), .B(_73_), .C(_74_), .Y(_0__9_) );
INVX1 INVX1_66 ( .A(_13_), .Y(_75_) );
NAND2X1 NAND2X1_123 ( .A(_14_), .B(w_cout_2_), .Y(_76_) );
OAI21X1 OAI21X1_122 ( .A(w_cout_2_), .B(_75_), .C(_76_), .Y(w_cout_3_) );
INVX1 INVX1_67 ( .A(_15__0_), .Y(_77_) );
NAND2X1 NAND2X1_124 ( .A(_16__0_), .B(w_cout_2_), .Y(_78_) );
OAI21X1 OAI21X1_123 ( .A(w_cout_2_), .B(_77_), .C(_78_), .Y(_0__10_) );
INVX1 INVX1_68 ( .A(_15__1_), .Y(_79_) );
NAND2X1 NAND2X1_125 ( .A(w_cout_2_), .B(_16__1_), .Y(_80_) );
OAI21X1 OAI21X1_124 ( .A(w_cout_2_), .B(_79_), .C(_80_), .Y(_0__11_) );
INVX1 INVX1_69 ( .A(_15__2_), .Y(_81_) );
NAND2X1 NAND2X1_126 ( .A(w_cout_2_), .B(_16__2_), .Y(_82_) );
OAI21X1 OAI21X1_125 ( .A(w_cout_2_), .B(_81_), .C(_82_), .Y(_0__12_) );
INVX1 INVX1_70 ( .A(_15__3_), .Y(_83_) );
NAND2X1 NAND2X1_127 ( .A(w_cout_2_), .B(_16__3_), .Y(_84_) );
OAI21X1 OAI21X1_126 ( .A(w_cout_2_), .B(_83_), .C(_84_), .Y(_0__13_) );
INVX1 INVX1_71 ( .A(_19_), .Y(_85_) );
NAND2X1 NAND2X1_128 ( .A(_20_), .B(w_cout_3_), .Y(_86_) );
OAI21X1 OAI21X1_127 ( .A(w_cout_3_), .B(_85_), .C(_86_), .Y(w_cout_4_) );
INVX1 INVX1_72 ( .A(_21__0_), .Y(_87_) );
NAND2X1 NAND2X1_129 ( .A(_22__0_), .B(w_cout_3_), .Y(_88_) );
OAI21X1 OAI21X1_128 ( .A(w_cout_3_), .B(_87_), .C(_88_), .Y(_0__14_) );
INVX1 INVX1_73 ( .A(_21__1_), .Y(_89_) );
NAND2X1 NAND2X1_130 ( .A(w_cout_3_), .B(_22__1_), .Y(_90_) );
OAI21X1 OAI21X1_129 ( .A(w_cout_3_), .B(_89_), .C(_90_), .Y(_0__15_) );
INVX1 INVX1_74 ( .A(_21__2_), .Y(_91_) );
NAND2X1 NAND2X1_131 ( .A(w_cout_3_), .B(_22__2_), .Y(_92_) );
OAI21X1 OAI21X1_130 ( .A(w_cout_3_), .B(_91_), .C(_92_), .Y(_0__16_) );
INVX1 INVX1_75 ( .A(_21__3_), .Y(_93_) );
NAND2X1 NAND2X1_132 ( .A(w_cout_3_), .B(_22__3_), .Y(_94_) );
OAI21X1 OAI21X1_131 ( .A(w_cout_3_), .B(_93_), .C(_94_), .Y(_0__17_) );
INVX1 INVX1_76 ( .A(_25_), .Y(_95_) );
NAND2X1 NAND2X1_133 ( .A(_26_), .B(w_cout_4_), .Y(_96_) );
OAI21X1 OAI21X1_132 ( .A(w_cout_4_), .B(_95_), .C(_96_), .Y(w_cout_5_) );
INVX1 INVX1_77 ( .A(_27__0_), .Y(_97_) );
NAND2X1 NAND2X1_134 ( .A(_28__0_), .B(w_cout_4_), .Y(_98_) );
OAI21X1 OAI21X1_133 ( .A(w_cout_4_), .B(_97_), .C(_98_), .Y(_0__18_) );
INVX1 INVX1_78 ( .A(_27__1_), .Y(_99_) );
NAND2X1 NAND2X1_135 ( .A(w_cout_4_), .B(_28__1_), .Y(_100_) );
OAI21X1 OAI21X1_134 ( .A(w_cout_4_), .B(_99_), .C(_100_), .Y(_0__19_) );
INVX1 INVX1_79 ( .A(_27__2_), .Y(_101_) );
NAND2X1 NAND2X1_136 ( .A(w_cout_4_), .B(_28__2_), .Y(_102_) );
OAI21X1 OAI21X1_135 ( .A(w_cout_4_), .B(_101_), .C(_102_), .Y(_0__20_) );
INVX1 INVX1_80 ( .A(_27__3_), .Y(_103_) );
NAND2X1 NAND2X1_137 ( .A(w_cout_4_), .B(_28__3_), .Y(_104_) );
OAI21X1 OAI21X1_136 ( .A(w_cout_4_), .B(_103_), .C(_104_), .Y(_0__21_) );
INVX1 INVX1_81 ( .A(_31_), .Y(_105_) );
NAND2X1 NAND2X1_138 ( .A(_32_), .B(w_cout_5_), .Y(_106_) );
OAI21X1 OAI21X1_137 ( .A(w_cout_5_), .B(_105_), .C(_106_), .Y(w_cout_6_) );
INVX1 INVX1_82 ( .A(_33__0_), .Y(_107_) );
NAND2X1 NAND2X1_139 ( .A(_34__0_), .B(w_cout_5_), .Y(_108_) );
OAI21X1 OAI21X1_138 ( .A(w_cout_5_), .B(_107_), .C(_108_), .Y(_0__22_) );
INVX1 INVX1_83 ( .A(_33__1_), .Y(_109_) );
NAND2X1 NAND2X1_140 ( .A(w_cout_5_), .B(_34__1_), .Y(_110_) );
OAI21X1 OAI21X1_139 ( .A(w_cout_5_), .B(_109_), .C(_110_), .Y(_0__23_) );
INVX1 INVX1_84 ( .A(_33__2_), .Y(_111_) );
NAND2X1 NAND2X1_141 ( .A(w_cout_5_), .B(_34__2_), .Y(_112_) );
OAI21X1 OAI21X1_140 ( .A(w_cout_5_), .B(_111_), .C(_112_), .Y(_0__24_) );
INVX1 INVX1_85 ( .A(_33__3_), .Y(_113_) );
NAND2X1 NAND2X1_142 ( .A(w_cout_5_), .B(_34__3_), .Y(_114_) );
OAI21X1 OAI21X1_141 ( .A(w_cout_5_), .B(_113_), .C(_114_), .Y(_0__25_) );
INVX1 INVX1_86 ( .A(_37_), .Y(_115_) );
NAND2X1 NAND2X1_143 ( .A(_38_), .B(w_cout_6_), .Y(_116_) );
OAI21X1 OAI21X1_142 ( .A(w_cout_6_), .B(_115_), .C(_116_), .Y(w_cout_7_) );
INVX1 INVX1_87 ( .A(_39__0_), .Y(_117_) );
NAND2X1 NAND2X1_144 ( .A(_40__0_), .B(w_cout_6_), .Y(_118_) );
OAI21X1 OAI21X1_143 ( .A(w_cout_6_), .B(_117_), .C(_118_), .Y(_0__26_) );
INVX1 INVX1_88 ( .A(_39__1_), .Y(_119_) );
NAND2X1 NAND2X1_145 ( .A(w_cout_6_), .B(_40__1_), .Y(_120_) );
OAI21X1 OAI21X1_144 ( .A(w_cout_6_), .B(_119_), .C(_120_), .Y(_0__27_) );
INVX1 INVX1_89 ( .A(_39__2_), .Y(_121_) );
NAND2X1 NAND2X1_146 ( .A(w_cout_6_), .B(_40__2_), .Y(_122_) );
OAI21X1 OAI21X1_145 ( .A(w_cout_6_), .B(_121_), .C(_122_), .Y(_0__28_) );
INVX1 INVX1_90 ( .A(_39__3_), .Y(_123_) );
NAND2X1 NAND2X1_147 ( .A(w_cout_6_), .B(_40__3_), .Y(_124_) );
OAI21X1 OAI21X1_146 ( .A(w_cout_6_), .B(_123_), .C(_124_), .Y(_0__29_) );
INVX1 INVX1_91 ( .A(_43_), .Y(_125_) );
NAND2X1 NAND2X1_148 ( .A(_44_), .B(w_cout_7_), .Y(_126_) );
OAI21X1 OAI21X1_147 ( .A(w_cout_7_), .B(_125_), .C(_126_), .Y(w_cout_8_) );
INVX1 INVX1_92 ( .A(_45__0_), .Y(_127_) );
NAND2X1 NAND2X1_149 ( .A(_46__0_), .B(w_cout_7_), .Y(_128_) );
OAI21X1 OAI21X1_148 ( .A(w_cout_7_), .B(_127_), .C(_128_), .Y(_0__30_) );
INVX1 INVX1_93 ( .A(_45__1_), .Y(_129_) );
NAND2X1 NAND2X1_150 ( .A(w_cout_7_), .B(_46__1_), .Y(_130_) );
OAI21X1 OAI21X1_149 ( .A(w_cout_7_), .B(_129_), .C(_130_), .Y(_0__31_) );
INVX1 INVX1_94 ( .A(_45__2_), .Y(_131_) );
NAND2X1 NAND2X1_151 ( .A(w_cout_7_), .B(_46__2_), .Y(_132_) );
OAI21X1 OAI21X1_150 ( .A(w_cout_7_), .B(_131_), .C(_132_), .Y(_0__32_) );
INVX1 INVX1_95 ( .A(_45__3_), .Y(_133_) );
NAND2X1 NAND2X1_152 ( .A(w_cout_7_), .B(_46__3_), .Y(_134_) );
OAI21X1 OAI21X1_151 ( .A(w_cout_7_), .B(_133_), .C(_134_), .Y(_0__33_) );
INVX1 INVX1_96 ( .A(_49_), .Y(_135_) );
NAND2X1 NAND2X1_153 ( .A(_50_), .B(w_cout_8_), .Y(_136_) );
OAI21X1 OAI21X1_152 ( .A(w_cout_8_), .B(_135_), .C(_136_), .Y(w_cout_9_) );
INVX1 INVX1_97 ( .A(_51__0_), .Y(_137_) );
NAND2X1 NAND2X1_154 ( .A(_52__0_), .B(w_cout_8_), .Y(_138_) );
OAI21X1 OAI21X1_153 ( .A(w_cout_8_), .B(_137_), .C(_138_), .Y(_0__34_) );
INVX1 INVX1_98 ( .A(_51__1_), .Y(_139_) );
NAND2X1 NAND2X1_155 ( .A(w_cout_8_), .B(_52__1_), .Y(_140_) );
OAI21X1 OAI21X1_154 ( .A(w_cout_8_), .B(_139_), .C(_140_), .Y(_0__35_) );
INVX1 INVX1_99 ( .A(_51__2_), .Y(_141_) );
NAND2X1 NAND2X1_156 ( .A(w_cout_8_), .B(_52__2_), .Y(_142_) );
OAI21X1 OAI21X1_155 ( .A(w_cout_8_), .B(_141_), .C(_142_), .Y(_0__36_) );
INVX1 INVX1_100 ( .A(_51__3_), .Y(_143_) );
NAND2X1 NAND2X1_157 ( .A(w_cout_8_), .B(_52__3_), .Y(_144_) );
OAI21X1 OAI21X1_156 ( .A(w_cout_8_), .B(_143_), .C(_144_), .Y(_0__37_) );
INVX1 INVX1_101 ( .A(1'b0), .Y(_148_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_149_) );
NAND2X1 NAND2X1_158 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_150_) );
NAND3X1 NAND3X1_57 ( .A(_148_), .B(_150_), .C(_149_), .Y(_151_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_145_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_146_) );
OAI21X1 OAI21X1_157 ( .A(_145_), .B(_146_), .C(1'b0), .Y(_147_) );
NAND2X1 NAND2X1_159 ( .A(_147_), .B(_151_), .Y(_3__0_) );
OAI21X1 OAI21X1_158 ( .A(_148_), .B(_145_), .C(_150_), .Y(_5__1_) );
INVX1 INVX1_102 ( .A(_5__1_), .Y(_155_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_156_) );
NAND2X1 NAND2X1_160 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_157_) );
NAND3X1 NAND3X1_58 ( .A(_155_), .B(_157_), .C(_156_), .Y(_158_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_152_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_153_) );
OAI21X1 OAI21X1_159 ( .A(_152_), .B(_153_), .C(_5__1_), .Y(_154_) );
NAND2X1 NAND2X1_161 ( .A(_154_), .B(_158_), .Y(_3__1_) );
OAI21X1 OAI21X1_160 ( .A(_155_), .B(_152_), .C(_157_), .Y(_5__2_) );
INVX1 INVX1_103 ( .A(_5__2_), .Y(_162_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_163_) );
NAND2X1 NAND2X1_162 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_164_) );
NAND3X1 NAND3X1_59 ( .A(_162_), .B(_164_), .C(_163_), .Y(_165_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_159_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_160_) );
OAI21X1 OAI21X1_161 ( .A(_159_), .B(_160_), .C(_5__2_), .Y(_161_) );
NAND2X1 NAND2X1_163 ( .A(_161_), .B(_165_), .Y(_3__2_) );
OAI21X1 OAI21X1_162 ( .A(_162_), .B(_159_), .C(_164_), .Y(_5__3_) );
INVX1 INVX1_104 ( .A(_5__3_), .Y(_169_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_170_) );
NAND2X1 NAND2X1_164 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_171_) );
NAND3X1 NAND3X1_60 ( .A(_169_), .B(_171_), .C(_170_), .Y(_172_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_166_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_167_) );
OAI21X1 OAI21X1_163 ( .A(_166_), .B(_167_), .C(_5__3_), .Y(_168_) );
NAND2X1 NAND2X1_165 ( .A(_168_), .B(_172_), .Y(_3__3_) );
OAI21X1 OAI21X1_164 ( .A(_169_), .B(_166_), .C(_171_), .Y(_1_) );
INVX1 INVX1_105 ( .A(1'b1), .Y(_176_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_177_) );
NAND2X1 NAND2X1_166 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_178_) );
NAND3X1 NAND3X1_61 ( .A(_176_), .B(_178_), .C(_177_), .Y(_179_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_173_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_174_) );
OAI21X1 OAI21X1_165 ( .A(_173_), .B(_174_), .C(1'b1), .Y(_175_) );
NAND2X1 NAND2X1_167 ( .A(_175_), .B(_179_), .Y(_4__0_) );
OAI21X1 OAI21X1_166 ( .A(_176_), .B(_173_), .C(_178_), .Y(_6__1_) );
INVX1 INVX1_106 ( .A(_6__1_), .Y(_183_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_184_) );
NAND2X1 NAND2X1_168 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_185_) );
NAND3X1 NAND3X1_62 ( .A(_183_), .B(_185_), .C(_184_), .Y(_186_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_180_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_181_) );
OAI21X1 OAI21X1_167 ( .A(_180_), .B(_181_), .C(_6__1_), .Y(_182_) );
NAND2X1 NAND2X1_169 ( .A(_182_), .B(_186_), .Y(_4__1_) );
OAI21X1 OAI21X1_168 ( .A(_183_), .B(_180_), .C(_185_), .Y(_6__2_) );
INVX1 INVX1_107 ( .A(_6__2_), .Y(_190_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_191_) );
NAND2X1 NAND2X1_170 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_192_) );
NAND3X1 NAND3X1_63 ( .A(_190_), .B(_192_), .C(_191_), .Y(_193_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_187_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_188_) );
OAI21X1 OAI21X1_169 ( .A(_187_), .B(_188_), .C(_6__2_), .Y(_189_) );
NAND2X1 NAND2X1_171 ( .A(_189_), .B(_193_), .Y(_4__2_) );
OAI21X1 OAI21X1_170 ( .A(_190_), .B(_187_), .C(_192_), .Y(_6__3_) );
INVX1 INVX1_108 ( .A(_6__3_), .Y(_197_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_198_) );
NAND2X1 NAND2X1_172 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_199_) );
NAND3X1 NAND3X1_64 ( .A(_197_), .B(_199_), .C(_198_), .Y(_200_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_194_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_195_) );
OAI21X1 OAI21X1_171 ( .A(_194_), .B(_195_), .C(_6__3_), .Y(_196_) );
NAND2X1 NAND2X1_173 ( .A(_196_), .B(_200_), .Y(_4__3_) );
OAI21X1 OAI21X1_172 ( .A(_197_), .B(_194_), .C(_199_), .Y(_2_) );
INVX1 INVX1_109 ( .A(1'b0), .Y(_204_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_205_) );
NAND2X1 NAND2X1_174 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_206_) );
NAND3X1 NAND3X1_65 ( .A(_204_), .B(_206_), .C(_205_), .Y(_207_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_201_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_202_) );
OAI21X1 OAI21X1_173 ( .A(_201_), .B(_202_), .C(1'b0), .Y(_203_) );
NAND2X1 NAND2X1_175 ( .A(_203_), .B(_207_), .Y(_9__0_) );
OAI21X1 OAI21X1_174 ( .A(_204_), .B(_201_), .C(_206_), .Y(_11__1_) );
INVX1 INVX1_110 ( .A(_11__1_), .Y(_211_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_212_) );
NAND2X1 NAND2X1_176 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_213_) );
NAND3X1 NAND3X1_66 ( .A(_211_), .B(_213_), .C(_212_), .Y(_214_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_208_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_209_) );
OAI21X1 OAI21X1_175 ( .A(_208_), .B(_209_), .C(_11__1_), .Y(_210_) );
NAND2X1 NAND2X1_177 ( .A(_210_), .B(_214_), .Y(_9__1_) );
OAI21X1 OAI21X1_176 ( .A(_211_), .B(_208_), .C(_213_), .Y(_11__2_) );
INVX1 INVX1_111 ( .A(_11__2_), .Y(_218_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_219_) );
NAND2X1 NAND2X1_178 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_220_) );
NAND3X1 NAND3X1_67 ( .A(_218_), .B(_220_), .C(_219_), .Y(_221_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_215_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_216_) );
OAI21X1 OAI21X1_177 ( .A(_215_), .B(_216_), .C(_11__2_), .Y(_217_) );
NAND2X1 NAND2X1_179 ( .A(_217_), .B(_221_), .Y(_9__2_) );
OAI21X1 OAI21X1_178 ( .A(_218_), .B(_215_), .C(_220_), .Y(_11__3_) );
INVX1 INVX1_112 ( .A(_11__3_), .Y(_225_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_226_) );
NAND2X1 NAND2X1_180 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_227_) );
NAND3X1 NAND3X1_68 ( .A(_225_), .B(_227_), .C(_226_), .Y(_228_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_222_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_223_) );
OAI21X1 OAI21X1_179 ( .A(_222_), .B(_223_), .C(_11__3_), .Y(_224_) );
NAND2X1 NAND2X1_181 ( .A(_224_), .B(_228_), .Y(_9__3_) );
OAI21X1 OAI21X1_180 ( .A(_225_), .B(_222_), .C(_227_), .Y(_7_) );
INVX1 INVX1_113 ( .A(1'b1), .Y(_232_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_233_) );
NAND2X1 NAND2X1_182 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_234_) );
NAND3X1 NAND3X1_69 ( .A(_232_), .B(_234_), .C(_233_), .Y(_235_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_229_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_230_) );
OAI21X1 OAI21X1_181 ( .A(_229_), .B(_230_), .C(1'b1), .Y(_231_) );
NAND2X1 NAND2X1_183 ( .A(_231_), .B(_235_), .Y(_10__0_) );
OAI21X1 OAI21X1_182 ( .A(_232_), .B(_229_), .C(_234_), .Y(_12__1_) );
INVX1 INVX1_114 ( .A(_12__1_), .Y(_239_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_240_) );
NAND2X1 NAND2X1_184 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_241_) );
NAND3X1 NAND3X1_70 ( .A(_239_), .B(_241_), .C(_240_), .Y(_242_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_236_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_237_) );
OAI21X1 OAI21X1_183 ( .A(_236_), .B(_237_), .C(_12__1_), .Y(_238_) );
NAND2X1 NAND2X1_185 ( .A(_238_), .B(_242_), .Y(_10__1_) );
OAI21X1 OAI21X1_184 ( .A(_239_), .B(_236_), .C(_241_), .Y(_12__2_) );
INVX1 INVX1_115 ( .A(_12__2_), .Y(_246_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_247_) );
NAND2X1 NAND2X1_186 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_248_) );
NAND3X1 NAND3X1_71 ( .A(_246_), .B(_248_), .C(_247_), .Y(_249_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_243_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_244_) );
OAI21X1 OAI21X1_185 ( .A(_243_), .B(_244_), .C(_12__2_), .Y(_245_) );
NAND2X1 NAND2X1_187 ( .A(_245_), .B(_249_), .Y(_10__2_) );
OAI21X1 OAI21X1_186 ( .A(_246_), .B(_243_), .C(_248_), .Y(_12__3_) );
INVX1 INVX1_116 ( .A(_12__3_), .Y(_253_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_254_) );
NAND2X1 NAND2X1_188 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_255_) );
NAND3X1 NAND3X1_72 ( .A(_253_), .B(_255_), .C(_254_), .Y(_256_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_250_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_251_) );
OAI21X1 OAI21X1_187 ( .A(_250_), .B(_251_), .C(_12__3_), .Y(_252_) );
NAND2X1 NAND2X1_189 ( .A(_252_), .B(_256_), .Y(_10__3_) );
OAI21X1 OAI21X1_188 ( .A(_253_), .B(_250_), .C(_255_), .Y(_8_) );
INVX1 INVX1_117 ( .A(1'b0), .Y(_260_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_261_) );
NAND2X1 NAND2X1_190 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_262_) );
NAND3X1 NAND3X1_73 ( .A(_260_), .B(_262_), .C(_261_), .Y(_263_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_257_) );
AND2X2 AND2X2_73 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_258_) );
OAI21X1 OAI21X1_189 ( .A(_257_), .B(_258_), .C(1'b0), .Y(_259_) );
NAND2X1 NAND2X1_191 ( .A(_259_), .B(_263_), .Y(_15__0_) );
OAI21X1 OAI21X1_190 ( .A(_260_), .B(_257_), .C(_262_), .Y(_17__1_) );
INVX1 INVX1_118 ( .A(_17__1_), .Y(_267_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_268_) );
NAND2X1 NAND2X1_192 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_269_) );
NAND3X1 NAND3X1_74 ( .A(_267_), .B(_269_), .C(_268_), .Y(_270_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_264_) );
AND2X2 AND2X2_74 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_265_) );
OAI21X1 OAI21X1_191 ( .A(_264_), .B(_265_), .C(_17__1_), .Y(_266_) );
NAND2X1 NAND2X1_193 ( .A(_266_), .B(_270_), .Y(_15__1_) );
OAI21X1 OAI21X1_192 ( .A(_267_), .B(_264_), .C(_269_), .Y(_17__2_) );
INVX1 INVX1_119 ( .A(_17__2_), .Y(_274_) );
BUFX2 BUFX2_40 ( .A(1'b0), .Y(_5__0_) );
BUFX2 BUFX2_41 ( .A(_1_), .Y(_5__4_) );
BUFX2 BUFX2_42 ( .A(1'b1), .Y(_6__0_) );
BUFX2 BUFX2_43 ( .A(_2_), .Y(_6__4_) );
BUFX2 BUFX2_44 ( .A(1'b0), .Y(_11__0_) );
BUFX2 BUFX2_45 ( .A(_7_), .Y(_11__4_) );
BUFX2 BUFX2_46 ( .A(1'b1), .Y(_12__0_) );
BUFX2 BUFX2_47 ( .A(_8_), .Y(_12__4_) );
BUFX2 BUFX2_48 ( .A(1'b0), .Y(_17__0_) );
BUFX2 BUFX2_49 ( .A(_13_), .Y(_17__4_) );
BUFX2 BUFX2_50 ( .A(1'b1), .Y(_18__0_) );
BUFX2 BUFX2_51 ( .A(_14_), .Y(_18__4_) );
BUFX2 BUFX2_52 ( .A(1'b0), .Y(_23__0_) );
BUFX2 BUFX2_53 ( .A(_19_), .Y(_23__4_) );
BUFX2 BUFX2_54 ( .A(1'b1), .Y(_24__0_) );
BUFX2 BUFX2_55 ( .A(_20_), .Y(_24__4_) );
BUFX2 BUFX2_56 ( .A(1'b0), .Y(_29__0_) );
BUFX2 BUFX2_57 ( .A(_25_), .Y(_29__4_) );
BUFX2 BUFX2_58 ( .A(1'b1), .Y(_30__0_) );
BUFX2 BUFX2_59 ( .A(_26_), .Y(_30__4_) );
BUFX2 BUFX2_60 ( .A(1'b0), .Y(_35__0_) );
BUFX2 BUFX2_61 ( .A(_31_), .Y(_35__4_) );
BUFX2 BUFX2_62 ( .A(1'b1), .Y(_36__0_) );
BUFX2 BUFX2_63 ( .A(_32_), .Y(_36__4_) );
BUFX2 BUFX2_64 ( .A(1'b0), .Y(_41__0_) );
BUFX2 BUFX2_65 ( .A(_37_), .Y(_41__4_) );
BUFX2 BUFX2_66 ( .A(1'b1), .Y(_42__0_) );
BUFX2 BUFX2_67 ( .A(_38_), .Y(_42__4_) );
BUFX2 BUFX2_68 ( .A(1'b0), .Y(_47__0_) );
BUFX2 BUFX2_69 ( .A(_43_), .Y(_47__4_) );
BUFX2 BUFX2_70 ( .A(1'b1), .Y(_48__0_) );
BUFX2 BUFX2_71 ( .A(_44_), .Y(_48__4_) );
BUFX2 BUFX2_72 ( .A(1'b0), .Y(_53__0_) );
BUFX2 BUFX2_73 ( .A(_49_), .Y(_53__4_) );
BUFX2 BUFX2_74 ( .A(1'b1), .Y(_54__0_) );
BUFX2 BUFX2_75 ( .A(_50_), .Y(_54__4_) );
BUFX2 BUFX2_76 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_77 ( .A(1'b0), .Y(w_cout_0_) );
endmodule
