module CSkipA_36bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_8_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
INVX1 INVX1_1 ( .A(skip0_cin_next), .Y(_28_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_29_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_30_) );
NAND3X1 NAND3X1_1 ( .A(_28_), .B(_30_), .C(_29_), .Y(_31_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_25_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_26_) );
OAI21X1 OAI21X1_1 ( .A(_25_), .B(_26_), .C(skip0_cin_next), .Y(_27_) );
NAND2X1 NAND2X1_2 ( .A(_27_), .B(_31_), .Y(_0__4_) );
OAI21X1 OAI21X1_2 ( .A(_28_), .B(_25_), .C(_30_), .Y(_2__1_) );
INVX1 INVX1_2 ( .A(_2__3_), .Y(_35_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_36_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_37_) );
NAND3X1 NAND3X1_2 ( .A(_35_), .B(_37_), .C(_36_), .Y(_38_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_32_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_33_) );
OAI21X1 OAI21X1_3 ( .A(_32_), .B(_33_), .C(_2__3_), .Y(_34_) );
NAND2X1 NAND2X1_4 ( .A(_34_), .B(_38_), .Y(_0__7_) );
OAI21X1 OAI21X1_4 ( .A(_35_), .B(_32_), .C(_37_), .Y(_1_) );
INVX1 INVX1_3 ( .A(_2__1_), .Y(_42_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_43_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_44_) );
NAND3X1 NAND3X1_3 ( .A(_42_), .B(_44_), .C(_43_), .Y(_45_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_39_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_40_) );
OAI21X1 OAI21X1_5 ( .A(_39_), .B(_40_), .C(_2__1_), .Y(_41_) );
NAND2X1 NAND2X1_6 ( .A(_41_), .B(_45_), .Y(_0__5_) );
OAI21X1 OAI21X1_6 ( .A(_42_), .B(_39_), .C(_44_), .Y(_2__2_) );
INVX1 INVX1_4 ( .A(_2__2_), .Y(_49_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_50_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_51_) );
NAND3X1 NAND3X1_4 ( .A(_49_), .B(_51_), .C(_50_), .Y(_52_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_46_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_47_) );
OAI21X1 OAI21X1_7 ( .A(_46_), .B(_47_), .C(_2__2_), .Y(_48_) );
NAND2X1 NAND2X1_8 ( .A(_48_), .B(_52_), .Y(_0__6_) );
OAI21X1 OAI21X1_8 ( .A(_49_), .B(_46_), .C(_51_), .Y(_2__3_) );
INVX1 INVX1_5 ( .A(i_add_term1[4]), .Y(_53_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[4]), .B(_53_), .Y(_54_) );
INVX1 INVX1_6 ( .A(i_add_term2[4]), .Y(_55_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term1[4]), .B(_55_), .Y(_56_) );
INVX1 INVX1_7 ( .A(i_add_term1[5]), .Y(_57_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[5]), .B(_57_), .Y(_58_) );
INVX1 INVX1_8 ( .A(i_add_term2[5]), .Y(_59_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term1[5]), .B(_59_), .Y(_60_) );
OAI22X1 OAI22X1_1 ( .A(_54_), .B(_56_), .C(_58_), .D(_60_), .Y(_61_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_62_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_63_) );
NOR2X1 NOR2X1_10 ( .A(_62_), .B(_63_), .Y(_64_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_65_) );
NAND2X1 NAND2X1_9 ( .A(_64_), .B(_65_), .Y(_66_) );
NOR2X1 NOR2X1_11 ( .A(_61_), .B(_66_), .Y(_3_) );
INVX1 INVX1_9 ( .A(_1_), .Y(_67_) );
NAND2X1 NAND2X1_10 ( .A(1'b0), .B(_3_), .Y(_68_) );
OAI21X1 OAI21X1_9 ( .A(_3_), .B(_67_), .C(_68_), .Y(w_cout_1_) );
INVX1 INVX1_10 ( .A(w_cout_1_), .Y(_72_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_73_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_74_) );
NAND3X1 NAND3X1_5 ( .A(_72_), .B(_74_), .C(_73_), .Y(_75_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_69_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_70_) );
OAI21X1 OAI21X1_10 ( .A(_69_), .B(_70_), .C(w_cout_1_), .Y(_71_) );
NAND2X1 NAND2X1_12 ( .A(_71_), .B(_75_), .Y(_0__8_) );
OAI21X1 OAI21X1_11 ( .A(_72_), .B(_69_), .C(_74_), .Y(_5__1_) );
INVX1 INVX1_11 ( .A(_5__3_), .Y(_79_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_80_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_81_) );
NAND3X1 NAND3X1_6 ( .A(_79_), .B(_81_), .C(_80_), .Y(_82_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_76_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_77_) );
OAI21X1 OAI21X1_12 ( .A(_76_), .B(_77_), .C(_5__3_), .Y(_78_) );
NAND2X1 NAND2X1_14 ( .A(_78_), .B(_82_), .Y(_0__11_) );
OAI21X1 OAI21X1_13 ( .A(_79_), .B(_76_), .C(_81_), .Y(_4_) );
INVX1 INVX1_12 ( .A(_5__1_), .Y(_86_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_87_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_88_) );
NAND3X1 NAND3X1_7 ( .A(_86_), .B(_88_), .C(_87_), .Y(_89_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_83_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_84_) );
OAI21X1 OAI21X1_14 ( .A(_83_), .B(_84_), .C(_5__1_), .Y(_85_) );
NAND2X1 NAND2X1_16 ( .A(_85_), .B(_89_), .Y(_0__9_) );
OAI21X1 OAI21X1_15 ( .A(_86_), .B(_83_), .C(_88_), .Y(_5__2_) );
INVX1 INVX1_13 ( .A(_5__2_), .Y(_93_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_94_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_95_) );
NAND3X1 NAND3X1_8 ( .A(_93_), .B(_95_), .C(_94_), .Y(_96_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_90_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_91_) );
OAI21X1 OAI21X1_16 ( .A(_90_), .B(_91_), .C(_5__2_), .Y(_92_) );
NAND2X1 NAND2X1_18 ( .A(_92_), .B(_96_), .Y(_0__10_) );
OAI21X1 OAI21X1_17 ( .A(_93_), .B(_90_), .C(_95_), .Y(_5__3_) );
INVX1 INVX1_14 ( .A(i_add_term1[8]), .Y(_97_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[8]), .B(_97_), .Y(_98_) );
INVX1 INVX1_15 ( .A(i_add_term2[8]), .Y(_99_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term1[8]), .B(_99_), .Y(_100_) );
INVX1 INVX1_16 ( .A(i_add_term1[9]), .Y(_101_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[9]), .B(_101_), .Y(_102_) );
INVX1 INVX1_17 ( .A(i_add_term2[9]), .Y(_103_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term1[9]), .B(_103_), .Y(_104_) );
OAI22X1 OAI22X1_2 ( .A(_98_), .B(_100_), .C(_102_), .D(_104_), .Y(_105_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_106_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_107_) );
NOR2X1 NOR2X1_21 ( .A(_106_), .B(_107_), .Y(_108_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_109_) );
NAND2X1 NAND2X1_19 ( .A(_108_), .B(_109_), .Y(_110_) );
NOR2X1 NOR2X1_22 ( .A(_105_), .B(_110_), .Y(_6_) );
INVX1 INVX1_18 ( .A(_4_), .Y(_111_) );
NAND2X1 NAND2X1_20 ( .A(1'b0), .B(_6_), .Y(_112_) );
OAI21X1 OAI21X1_18 ( .A(_6_), .B(_111_), .C(_112_), .Y(w_cout_2_) );
INVX1 INVX1_19 ( .A(w_cout_2_), .Y(_116_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_117_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_118_) );
NAND3X1 NAND3X1_9 ( .A(_116_), .B(_118_), .C(_117_), .Y(_119_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_113_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_114_) );
OAI21X1 OAI21X1_19 ( .A(_113_), .B(_114_), .C(w_cout_2_), .Y(_115_) );
NAND2X1 NAND2X1_22 ( .A(_115_), .B(_119_), .Y(_0__12_) );
OAI21X1 OAI21X1_20 ( .A(_116_), .B(_113_), .C(_118_), .Y(_8__1_) );
INVX1 INVX1_20 ( .A(_8__3_), .Y(_123_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_124_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_125_) );
NAND3X1 NAND3X1_10 ( .A(_123_), .B(_125_), .C(_124_), .Y(_126_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_120_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_121_) );
OAI21X1 OAI21X1_21 ( .A(_120_), .B(_121_), .C(_8__3_), .Y(_122_) );
NAND2X1 NAND2X1_24 ( .A(_122_), .B(_126_), .Y(_0__15_) );
OAI21X1 OAI21X1_22 ( .A(_123_), .B(_120_), .C(_125_), .Y(_7_) );
INVX1 INVX1_21 ( .A(_8__1_), .Y(_130_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_131_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_132_) );
NAND3X1 NAND3X1_11 ( .A(_130_), .B(_132_), .C(_131_), .Y(_133_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_127_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_128_) );
OAI21X1 OAI21X1_23 ( .A(_127_), .B(_128_), .C(_8__1_), .Y(_129_) );
NAND2X1 NAND2X1_26 ( .A(_129_), .B(_133_), .Y(_0__13_) );
OAI21X1 OAI21X1_24 ( .A(_130_), .B(_127_), .C(_132_), .Y(_8__2_) );
INVX1 INVX1_22 ( .A(_8__2_), .Y(_137_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_138_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_139_) );
NAND3X1 NAND3X1_12 ( .A(_137_), .B(_139_), .C(_138_), .Y(_140_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_134_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_135_) );
OAI21X1 OAI21X1_25 ( .A(_134_), .B(_135_), .C(_8__2_), .Y(_136_) );
NAND2X1 NAND2X1_28 ( .A(_136_), .B(_140_), .Y(_0__14_) );
OAI21X1 OAI21X1_26 ( .A(_137_), .B(_134_), .C(_139_), .Y(_8__3_) );
INVX1 INVX1_23 ( .A(i_add_term1[12]), .Y(_141_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[12]), .B(_141_), .Y(_142_) );
INVX1 INVX1_24 ( .A(i_add_term2[12]), .Y(_143_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term1[12]), .B(_143_), .Y(_144_) );
INVX1 INVX1_25 ( .A(i_add_term1[13]), .Y(_145_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[13]), .B(_145_), .Y(_146_) );
INVX1 INVX1_26 ( .A(i_add_term2[13]), .Y(_147_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term1[13]), .B(_147_), .Y(_148_) );
OAI22X1 OAI22X1_3 ( .A(_142_), .B(_144_), .C(_146_), .D(_148_), .Y(_149_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_150_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_151_) );
NOR2X1 NOR2X1_32 ( .A(_150_), .B(_151_), .Y(_152_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_153_) );
NAND2X1 NAND2X1_29 ( .A(_152_), .B(_153_), .Y(_154_) );
NOR2X1 NOR2X1_33 ( .A(_149_), .B(_154_), .Y(_9_) );
INVX1 INVX1_27 ( .A(_7_), .Y(_155_) );
NAND2X1 NAND2X1_30 ( .A(1'b0), .B(_9_), .Y(_156_) );
OAI21X1 OAI21X1_27 ( .A(_9_), .B(_155_), .C(_156_), .Y(w_cout_3_) );
INVX1 INVX1_28 ( .A(w_cout_3_), .Y(_160_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_161_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_162_) );
NAND3X1 NAND3X1_13 ( .A(_160_), .B(_162_), .C(_161_), .Y(_163_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_157_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_158_) );
OAI21X1 OAI21X1_28 ( .A(_157_), .B(_158_), .C(w_cout_3_), .Y(_159_) );
NAND2X1 NAND2X1_32 ( .A(_159_), .B(_163_), .Y(_0__16_) );
OAI21X1 OAI21X1_29 ( .A(_160_), .B(_157_), .C(_162_), .Y(_11__1_) );
INVX1 INVX1_29 ( .A(_11__3_), .Y(_167_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_168_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_169_) );
NAND3X1 NAND3X1_14 ( .A(_167_), .B(_169_), .C(_168_), .Y(_170_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_164_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_165_) );
OAI21X1 OAI21X1_30 ( .A(_164_), .B(_165_), .C(_11__3_), .Y(_166_) );
NAND2X1 NAND2X1_34 ( .A(_166_), .B(_170_), .Y(_0__19_) );
OAI21X1 OAI21X1_31 ( .A(_167_), .B(_164_), .C(_169_), .Y(_10_) );
INVX1 INVX1_30 ( .A(_11__1_), .Y(_174_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_175_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_176_) );
NAND3X1 NAND3X1_15 ( .A(_174_), .B(_176_), .C(_175_), .Y(_177_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_171_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_172_) );
OAI21X1 OAI21X1_32 ( .A(_171_), .B(_172_), .C(_11__1_), .Y(_173_) );
NAND2X1 NAND2X1_36 ( .A(_173_), .B(_177_), .Y(_0__17_) );
OAI21X1 OAI21X1_33 ( .A(_174_), .B(_171_), .C(_176_), .Y(_11__2_) );
INVX1 INVX1_31 ( .A(_11__2_), .Y(_181_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_182_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_183_) );
NAND3X1 NAND3X1_16 ( .A(_181_), .B(_183_), .C(_182_), .Y(_184_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_178_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_179_) );
OAI21X1 OAI21X1_34 ( .A(_178_), .B(_179_), .C(_11__2_), .Y(_180_) );
NAND2X1 NAND2X1_38 ( .A(_180_), .B(_184_), .Y(_0__18_) );
OAI21X1 OAI21X1_35 ( .A(_181_), .B(_178_), .C(_183_), .Y(_11__3_) );
INVX1 INVX1_32 ( .A(i_add_term1[16]), .Y(_185_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[16]), .B(_185_), .Y(_186_) );
INVX1 INVX1_33 ( .A(i_add_term2[16]), .Y(_187_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term1[16]), .B(_187_), .Y(_188_) );
INVX1 INVX1_34 ( .A(i_add_term1[17]), .Y(_189_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[17]), .B(_189_), .Y(_190_) );
INVX1 INVX1_35 ( .A(i_add_term2[17]), .Y(_191_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term1[17]), .B(_191_), .Y(_192_) );
OAI22X1 OAI22X1_4 ( .A(_186_), .B(_188_), .C(_190_), .D(_192_), .Y(_193_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_194_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_195_) );
NOR2X1 NOR2X1_43 ( .A(_194_), .B(_195_), .Y(_196_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_197_) );
NAND2X1 NAND2X1_39 ( .A(_196_), .B(_197_), .Y(_198_) );
NOR2X1 NOR2X1_44 ( .A(_193_), .B(_198_), .Y(_12_) );
INVX1 INVX1_36 ( .A(_10_), .Y(_199_) );
NAND2X1 NAND2X1_40 ( .A(1'b0), .B(_12_), .Y(_200_) );
OAI21X1 OAI21X1_36 ( .A(_12_), .B(_199_), .C(_200_), .Y(w_cout_4_) );
INVX1 INVX1_37 ( .A(w_cout_4_), .Y(_204_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_205_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_206_) );
NAND3X1 NAND3X1_17 ( .A(_204_), .B(_206_), .C(_205_), .Y(_207_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_201_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_202_) );
OAI21X1 OAI21X1_37 ( .A(_201_), .B(_202_), .C(w_cout_4_), .Y(_203_) );
NAND2X1 NAND2X1_42 ( .A(_203_), .B(_207_), .Y(_0__20_) );
OAI21X1 OAI21X1_38 ( .A(_204_), .B(_201_), .C(_206_), .Y(_14__1_) );
INVX1 INVX1_38 ( .A(_14__3_), .Y(_211_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_212_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_213_) );
NAND3X1 NAND3X1_18 ( .A(_211_), .B(_213_), .C(_212_), .Y(_214_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_208_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_209_) );
OAI21X1 OAI21X1_39 ( .A(_208_), .B(_209_), .C(_14__3_), .Y(_210_) );
NAND2X1 NAND2X1_44 ( .A(_210_), .B(_214_), .Y(_0__23_) );
OAI21X1 OAI21X1_40 ( .A(_211_), .B(_208_), .C(_213_), .Y(_13_) );
INVX1 INVX1_39 ( .A(_14__1_), .Y(_218_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_219_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_220_) );
NAND3X1 NAND3X1_19 ( .A(_218_), .B(_220_), .C(_219_), .Y(_221_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_215_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_216_) );
OAI21X1 OAI21X1_41 ( .A(_215_), .B(_216_), .C(_14__1_), .Y(_217_) );
NAND2X1 NAND2X1_46 ( .A(_217_), .B(_221_), .Y(_0__21_) );
OAI21X1 OAI21X1_42 ( .A(_218_), .B(_215_), .C(_220_), .Y(_14__2_) );
INVX1 INVX1_40 ( .A(_14__2_), .Y(_225_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_226_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_227_) );
NAND3X1 NAND3X1_20 ( .A(_225_), .B(_227_), .C(_226_), .Y(_228_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_222_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_223_) );
OAI21X1 OAI21X1_43 ( .A(_222_), .B(_223_), .C(_14__2_), .Y(_224_) );
NAND2X1 NAND2X1_48 ( .A(_224_), .B(_228_), .Y(_0__22_) );
OAI21X1 OAI21X1_44 ( .A(_225_), .B(_222_), .C(_227_), .Y(_14__3_) );
INVX1 INVX1_41 ( .A(i_add_term1[20]), .Y(_229_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[20]), .B(_229_), .Y(_230_) );
INVX1 INVX1_42 ( .A(i_add_term2[20]), .Y(_231_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term1[20]), .B(_231_), .Y(_232_) );
INVX1 INVX1_43 ( .A(i_add_term1[21]), .Y(_233_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[21]), .B(_233_), .Y(_234_) );
INVX1 INVX1_44 ( .A(i_add_term2[21]), .Y(_235_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term1[21]), .B(_235_), .Y(_236_) );
OAI22X1 OAI22X1_5 ( .A(_230_), .B(_232_), .C(_234_), .D(_236_), .Y(_237_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_238_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_239_) );
NOR2X1 NOR2X1_54 ( .A(_238_), .B(_239_), .Y(_240_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_241_) );
NAND2X1 NAND2X1_49 ( .A(_240_), .B(_241_), .Y(_242_) );
NOR2X1 NOR2X1_55 ( .A(_237_), .B(_242_), .Y(_15_) );
INVX1 INVX1_45 ( .A(_13_), .Y(_243_) );
NAND2X1 NAND2X1_50 ( .A(1'b0), .B(_15_), .Y(_244_) );
OAI21X1 OAI21X1_45 ( .A(_15_), .B(_243_), .C(_244_), .Y(w_cout_5_) );
INVX1 INVX1_46 ( .A(w_cout_5_), .Y(_248_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_249_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_250_) );
NAND3X1 NAND3X1_21 ( .A(_248_), .B(_250_), .C(_249_), .Y(_251_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_245_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_246_) );
OAI21X1 OAI21X1_46 ( .A(_245_), .B(_246_), .C(w_cout_5_), .Y(_247_) );
NAND2X1 NAND2X1_52 ( .A(_247_), .B(_251_), .Y(_0__24_) );
OAI21X1 OAI21X1_47 ( .A(_248_), .B(_245_), .C(_250_), .Y(_17__1_) );
INVX1 INVX1_47 ( .A(_17__3_), .Y(_255_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_256_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_257_) );
NAND3X1 NAND3X1_22 ( .A(_255_), .B(_257_), .C(_256_), .Y(_258_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_252_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_253_) );
OAI21X1 OAI21X1_48 ( .A(_252_), .B(_253_), .C(_17__3_), .Y(_254_) );
NAND2X1 NAND2X1_54 ( .A(_254_), .B(_258_), .Y(_0__27_) );
OAI21X1 OAI21X1_49 ( .A(_255_), .B(_252_), .C(_257_), .Y(_16_) );
INVX1 INVX1_48 ( .A(_17__1_), .Y(_262_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_263_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_264_) );
NAND3X1 NAND3X1_23 ( .A(_262_), .B(_264_), .C(_263_), .Y(_265_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_259_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_260_) );
OAI21X1 OAI21X1_50 ( .A(_259_), .B(_260_), .C(_17__1_), .Y(_261_) );
NAND2X1 NAND2X1_56 ( .A(_261_), .B(_265_), .Y(_0__25_) );
OAI21X1 OAI21X1_51 ( .A(_262_), .B(_259_), .C(_264_), .Y(_17__2_) );
INVX1 INVX1_49 ( .A(_17__2_), .Y(_269_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_270_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_271_) );
NAND3X1 NAND3X1_24 ( .A(_269_), .B(_271_), .C(_270_), .Y(_272_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_266_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_267_) );
OAI21X1 OAI21X1_52 ( .A(_266_), .B(_267_), .C(_17__2_), .Y(_268_) );
NAND2X1 NAND2X1_58 ( .A(_268_), .B(_272_), .Y(_0__26_) );
OAI21X1 OAI21X1_53 ( .A(_269_), .B(_266_), .C(_271_), .Y(_17__3_) );
INVX1 INVX1_50 ( .A(i_add_term1[24]), .Y(_273_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[24]), .B(_273_), .Y(_274_) );
INVX1 INVX1_51 ( .A(i_add_term2[24]), .Y(_275_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term1[24]), .B(_275_), .Y(_276_) );
INVX1 INVX1_52 ( .A(i_add_term1[25]), .Y(_277_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[25]), .B(_277_), .Y(_278_) );
INVX1 INVX1_53 ( .A(i_add_term2[25]), .Y(_279_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term1[25]), .B(_279_), .Y(_280_) );
OAI22X1 OAI22X1_6 ( .A(_274_), .B(_276_), .C(_278_), .D(_280_), .Y(_281_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_282_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_283_) );
NOR2X1 NOR2X1_65 ( .A(_282_), .B(_283_), .Y(_284_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_285_) );
NAND2X1 NAND2X1_59 ( .A(_284_), .B(_285_), .Y(_286_) );
NOR2X1 NOR2X1_66 ( .A(_281_), .B(_286_), .Y(_18_) );
INVX1 INVX1_54 ( .A(_16_), .Y(_287_) );
NAND2X1 NAND2X1_60 ( .A(1'b0), .B(_18_), .Y(_288_) );
OAI21X1 OAI21X1_54 ( .A(_18_), .B(_287_), .C(_288_), .Y(w_cout_6_) );
INVX1 INVX1_55 ( .A(w_cout_6_), .Y(_292_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_293_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_294_) );
NAND3X1 NAND3X1_25 ( .A(_292_), .B(_294_), .C(_293_), .Y(_295_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_289_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_290_) );
OAI21X1 OAI21X1_55 ( .A(_289_), .B(_290_), .C(w_cout_6_), .Y(_291_) );
NAND2X1 NAND2X1_62 ( .A(_291_), .B(_295_), .Y(_0__28_) );
OAI21X1 OAI21X1_56 ( .A(_292_), .B(_289_), .C(_294_), .Y(_20__1_) );
INVX1 INVX1_56 ( .A(_20__3_), .Y(_299_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_300_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_301_) );
NAND3X1 NAND3X1_26 ( .A(_299_), .B(_301_), .C(_300_), .Y(_302_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_296_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_297_) );
OAI21X1 OAI21X1_57 ( .A(_296_), .B(_297_), .C(_20__3_), .Y(_298_) );
NAND2X1 NAND2X1_64 ( .A(_298_), .B(_302_), .Y(_0__31_) );
OAI21X1 OAI21X1_58 ( .A(_299_), .B(_296_), .C(_301_), .Y(_19_) );
INVX1 INVX1_57 ( .A(_20__1_), .Y(_306_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_307_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_308_) );
NAND3X1 NAND3X1_27 ( .A(_306_), .B(_308_), .C(_307_), .Y(_309_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_303_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_304_) );
OAI21X1 OAI21X1_59 ( .A(_303_), .B(_304_), .C(_20__1_), .Y(_305_) );
NAND2X1 NAND2X1_66 ( .A(_305_), .B(_309_), .Y(_0__29_) );
OAI21X1 OAI21X1_60 ( .A(_306_), .B(_303_), .C(_308_), .Y(_20__2_) );
INVX1 INVX1_58 ( .A(_20__2_), .Y(_313_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_314_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_315_) );
NAND3X1 NAND3X1_28 ( .A(_313_), .B(_315_), .C(_314_), .Y(_316_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_310_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_311_) );
OAI21X1 OAI21X1_61 ( .A(_310_), .B(_311_), .C(_20__2_), .Y(_312_) );
NAND2X1 NAND2X1_68 ( .A(_312_), .B(_316_), .Y(_0__30_) );
OAI21X1 OAI21X1_62 ( .A(_313_), .B(_310_), .C(_315_), .Y(_20__3_) );
INVX1 INVX1_59 ( .A(i_add_term1[28]), .Y(_317_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[28]), .B(_317_), .Y(_318_) );
INVX1 INVX1_60 ( .A(i_add_term2[28]), .Y(_319_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term1[28]), .B(_319_), .Y(_320_) );
INVX1 INVX1_61 ( .A(i_add_term1[29]), .Y(_321_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[29]), .B(_321_), .Y(_322_) );
INVX1 INVX1_62 ( .A(i_add_term2[29]), .Y(_323_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term1[29]), .B(_323_), .Y(_324_) );
OAI22X1 OAI22X1_7 ( .A(_318_), .B(_320_), .C(_322_), .D(_324_), .Y(_325_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_326_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_327_) );
NOR2X1 NOR2X1_76 ( .A(_326_), .B(_327_), .Y(_328_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_329_) );
NAND2X1 NAND2X1_69 ( .A(_328_), .B(_329_), .Y(_330_) );
NOR2X1 NOR2X1_77 ( .A(_325_), .B(_330_), .Y(_21_) );
INVX1 INVX1_63 ( .A(_19_), .Y(_331_) );
NAND2X1 NAND2X1_70 ( .A(1'b0), .B(_21_), .Y(_332_) );
OAI21X1 OAI21X1_63 ( .A(_21_), .B(_331_), .C(_332_), .Y(w_cout_7_) );
INVX1 INVX1_64 ( .A(w_cout_7_), .Y(_336_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_337_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_338_) );
NAND3X1 NAND3X1_29 ( .A(_336_), .B(_338_), .C(_337_), .Y(_339_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_333_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_334_) );
OAI21X1 OAI21X1_64 ( .A(_333_), .B(_334_), .C(w_cout_7_), .Y(_335_) );
NAND2X1 NAND2X1_72 ( .A(_335_), .B(_339_), .Y(_0__32_) );
OAI21X1 OAI21X1_65 ( .A(_336_), .B(_333_), .C(_338_), .Y(_23__1_) );
INVX1 INVX1_65 ( .A(_23__3_), .Y(_343_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_344_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_345_) );
NAND3X1 NAND3X1_30 ( .A(_343_), .B(_345_), .C(_344_), .Y(_346_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_340_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_341_) );
OAI21X1 OAI21X1_66 ( .A(_340_), .B(_341_), .C(_23__3_), .Y(_342_) );
NAND2X1 NAND2X1_74 ( .A(_342_), .B(_346_), .Y(_0__35_) );
OAI21X1 OAI21X1_67 ( .A(_343_), .B(_340_), .C(_345_), .Y(_22_) );
INVX1 INVX1_66 ( .A(_23__1_), .Y(_350_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_351_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_352_) );
NAND3X1 NAND3X1_31 ( .A(_350_), .B(_352_), .C(_351_), .Y(_353_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_347_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_348_) );
OAI21X1 OAI21X1_68 ( .A(_347_), .B(_348_), .C(_23__1_), .Y(_349_) );
NAND2X1 NAND2X1_76 ( .A(_349_), .B(_353_), .Y(_0__33_) );
OAI21X1 OAI21X1_69 ( .A(_350_), .B(_347_), .C(_352_), .Y(_23__2_) );
INVX1 INVX1_67 ( .A(_23__2_), .Y(_357_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_358_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_359_) );
NAND3X1 NAND3X1_32 ( .A(_357_), .B(_359_), .C(_358_), .Y(_360_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_354_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_355_) );
OAI21X1 OAI21X1_70 ( .A(_354_), .B(_355_), .C(_23__2_), .Y(_356_) );
NAND2X1 NAND2X1_78 ( .A(_356_), .B(_360_), .Y(_0__34_) );
OAI21X1 OAI21X1_71 ( .A(_357_), .B(_354_), .C(_359_), .Y(_23__3_) );
INVX1 INVX1_68 ( .A(i_add_term1[32]), .Y(_361_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[32]), .B(_361_), .Y(_362_) );
INVX1 INVX1_69 ( .A(i_add_term2[32]), .Y(_363_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term1[32]), .B(_363_), .Y(_364_) );
INVX1 INVX1_70 ( .A(i_add_term1[33]), .Y(_365_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[33]), .B(_365_), .Y(_366_) );
INVX1 INVX1_71 ( .A(i_add_term2[33]), .Y(_367_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term1[33]), .B(_367_), .Y(_368_) );
OAI22X1 OAI22X1_8 ( .A(_362_), .B(_364_), .C(_366_), .D(_368_), .Y(_369_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_370_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_371_) );
NOR2X1 NOR2X1_87 ( .A(_370_), .B(_371_), .Y(_372_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_373_) );
NAND2X1 NAND2X1_79 ( .A(_372_), .B(_373_), .Y(_374_) );
NOR2X1 NOR2X1_88 ( .A(_369_), .B(_374_), .Y(_24_) );
INVX1 INVX1_72 ( .A(_22_), .Y(_375_) );
NAND2X1 NAND2X1_80 ( .A(1'b0), .B(_24_), .Y(_376_) );
OAI21X1 OAI21X1_72 ( .A(_24_), .B(_375_), .C(_376_), .Y(w_cout_8_) );
INVX1 INVX1_73 ( .A(1'b0), .Y(_380_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_381_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_382_) );
NAND3X1 NAND3X1_33 ( .A(_380_), .B(_382_), .C(_381_), .Y(_383_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_377_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_378_) );
OAI21X1 OAI21X1_73 ( .A(_377_), .B(_378_), .C(1'b0), .Y(_379_) );
NAND2X1 NAND2X1_82 ( .A(_379_), .B(_383_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_74 ( .A(_380_), .B(_377_), .C(_382_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_74 ( .A(rca_inst_fa3_i_carry), .Y(_387_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_388_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_389_) );
NAND3X1 NAND3X1_34 ( .A(_387_), .B(_389_), .C(_388_), .Y(_390_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_384_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_385_) );
OAI21X1 OAI21X1_75 ( .A(_384_), .B(_385_), .C(rca_inst_fa3_i_carry), .Y(_386_) );
NAND2X1 NAND2X1_84 ( .A(_386_), .B(_390_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_76 ( .A(_387_), .B(_384_), .C(_389_), .Y(cout0) );
INVX1 INVX1_75 ( .A(rca_inst_fa0_o_carry), .Y(_394_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_395_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_396_) );
NAND3X1 NAND3X1_35 ( .A(_394_), .B(_396_), .C(_395_), .Y(_397_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_391_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_392_) );
OAI21X1 OAI21X1_77 ( .A(_391_), .B(_392_), .C(rca_inst_fa0_o_carry), .Y(_393_) );
NAND2X1 NAND2X1_86 ( .A(_393_), .B(_397_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_78 ( .A(_394_), .B(_391_), .C(_396_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_76 ( .A(rca_inst_fa_1__o_carry), .Y(_401_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_402_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_403_) );
NAND3X1 NAND3X1_36 ( .A(_401_), .B(_403_), .C(_402_), .Y(_404_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_398_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_399_) );
OAI21X1 OAI21X1_79 ( .A(_398_), .B(_399_), .C(rca_inst_fa_1__o_carry), .Y(_400_) );
NAND2X1 NAND2X1_88 ( .A(_400_), .B(_404_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_80 ( .A(_401_), .B(_398_), .C(_403_), .Y(rca_inst_fa3_i_carry) );
INVX1 INVX1_77 ( .A(i_add_term1[0]), .Y(_405_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[0]), .B(_405_), .Y(_406_) );
INVX1 INVX1_78 ( .A(i_add_term2[0]), .Y(_407_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term1[0]), .B(_407_), .Y(_408_) );
INVX1 INVX1_79 ( .A(i_add_term1[1]), .Y(_409_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[1]), .B(_409_), .Y(_410_) );
INVX1 INVX1_80 ( .A(i_add_term2[1]), .Y(_411_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term1[1]), .B(_411_), .Y(_412_) );
OAI22X1 OAI22X1_9 ( .A(_406_), .B(_408_), .C(_410_), .D(_412_), .Y(_413_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_414_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_415_) );
NOR2X1 NOR2X1_98 ( .A(_414_), .B(_415_), .Y(_416_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_417_) );
NAND2X1 NAND2X1_89 ( .A(_416_), .B(_417_), .Y(_418_) );
NOR2X1 NOR2X1_99 ( .A(_413_), .B(_418_), .Y(skip0_P) );
INVX1 INVX1_81 ( .A(cout0), .Y(_419_) );
NAND2X1 NAND2X1_90 ( .A(1'b0), .B(skip0_P), .Y(_420_) );
OAI21X1 OAI21X1_81 ( .A(skip0_P), .B(_419_), .C(_420_), .Y(skip0_cin_next) );
BUFX2 BUFX2_38 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_39 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_40 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_41 ( .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_42 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
