module cla_64bit (i_add1, i_add2, o_result);

input [63:0] i_add1;
input [63:0] i_add2;
output [64:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

NAND3X1 NAND3X1_1 ( .A(_139_), .B(_147_), .C(_144_), .Y(_148_) );
OAI21X1 OAI21X1_1 ( .A(i_add2[24]), .B(i_add1[24]), .C(_148_), .Y(_149_) );
INVX1 INVX1_1 ( .A(_149_), .Y(w_C_25_) );
INVX1 INVX1_2 ( .A(i_add2[25]), .Y(_150_) );
INVX1 INVX1_3 ( .A(i_add1[25]), .Y(_151_) );
NOR2X1 NOR2X1_1 ( .A(_150_), .B(_151_), .Y(_152_) );
INVX1 INVX1_4 ( .A(_152_), .Y(_153_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_154_) );
INVX1 INVX1_5 ( .A(_154_), .Y(_155_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_156_) );
INVX1 INVX1_6 ( .A(_156_), .Y(_157_) );
NAND3X1 NAND3X1_2 ( .A(_155_), .B(_157_), .C(_148_), .Y(_158_) );
AND2X2 AND2X2_1 ( .A(_158_), .B(_153_), .Y(_159_) );
INVX1 INVX1_7 ( .A(_159_), .Y(w_C_26_) );
AND2X2 AND2X2_2 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_160_) );
INVX1 INVX1_8 ( .A(_160_), .Y(_161_) );
NAND3X1 NAND3X1_3 ( .A(_153_), .B(_161_), .C(_158_), .Y(_162_) );
OAI21X1 OAI21X1_2 ( .A(i_add2[26]), .B(i_add1[26]), .C(_162_), .Y(_163_) );
INVX1 INVX1_9 ( .A(_163_), .Y(w_C_27_) );
INVX1 INVX1_10 ( .A(i_add2[27]), .Y(_164_) );
INVX1 INVX1_11 ( .A(i_add1[27]), .Y(_165_) );
NOR2X1 NOR2X1_4 ( .A(_164_), .B(_165_), .Y(_166_) );
INVX1 INVX1_12 ( .A(_166_), .Y(_167_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_168_) );
INVX1 INVX1_13 ( .A(_168_), .Y(_169_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_170_) );
INVX1 INVX1_14 ( .A(_170_), .Y(_171_) );
NAND3X1 NAND3X1_4 ( .A(_169_), .B(_171_), .C(_162_), .Y(_172_) );
AND2X2 AND2X2_3 ( .A(_172_), .B(_167_), .Y(_173_) );
INVX1 INVX1_15 ( .A(_173_), .Y(w_C_28_) );
AND2X2 AND2X2_4 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_174_) );
INVX1 INVX1_16 ( .A(_174_), .Y(_175_) );
NAND3X1 NAND3X1_5 ( .A(_167_), .B(_175_), .C(_172_), .Y(_176_) );
OAI21X1 OAI21X1_3 ( .A(i_add2[28]), .B(i_add1[28]), .C(_176_), .Y(_177_) );
INVX1 INVX1_17 ( .A(_177_), .Y(w_C_29_) );
INVX1 INVX1_18 ( .A(i_add2[29]), .Y(_178_) );
INVX1 INVX1_19 ( .A(i_add1[29]), .Y(_179_) );
NOR2X1 NOR2X1_7 ( .A(_178_), .B(_179_), .Y(_180_) );
INVX1 INVX1_20 ( .A(_180_), .Y(_181_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_182_) );
INVX1 INVX1_21 ( .A(_182_), .Y(_183_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_184_) );
INVX1 INVX1_22 ( .A(_184_), .Y(_185_) );
NAND3X1 NAND3X1_6 ( .A(_183_), .B(_185_), .C(_176_), .Y(_186_) );
AND2X2 AND2X2_5 ( .A(_186_), .B(_181_), .Y(_187_) );
INVX1 INVX1_23 ( .A(_187_), .Y(w_C_30_) );
AND2X2 AND2X2_6 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_188_) );
INVX1 INVX1_24 ( .A(_188_), .Y(_189_) );
NAND3X1 NAND3X1_7 ( .A(_181_), .B(_189_), .C(_186_), .Y(_190_) );
OAI21X1 OAI21X1_4 ( .A(i_add2[30]), .B(i_add1[30]), .C(_190_), .Y(_191_) );
INVX1 INVX1_25 ( .A(_191_), .Y(w_C_31_) );
INVX1 INVX1_26 ( .A(i_add2[31]), .Y(_192_) );
INVX1 INVX1_27 ( .A(i_add1[31]), .Y(_193_) );
NOR2X1 NOR2X1_10 ( .A(_192_), .B(_193_), .Y(_194_) );
INVX1 INVX1_28 ( .A(_194_), .Y(_195_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_196_) );
INVX1 INVX1_29 ( .A(_196_), .Y(_197_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_198_) );
INVX1 INVX1_30 ( .A(_198_), .Y(_199_) );
NAND3X1 NAND3X1_8 ( .A(_197_), .B(_199_), .C(_190_), .Y(_200_) );
AND2X2 AND2X2_7 ( .A(_200_), .B(_195_), .Y(_201_) );
INVX1 INVX1_31 ( .A(_201_), .Y(w_C_32_) );
AND2X2 AND2X2_8 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_202_) );
INVX1 INVX1_32 ( .A(_202_), .Y(_203_) );
NAND3X1 NAND3X1_9 ( .A(_195_), .B(_203_), .C(_200_), .Y(_204_) );
OAI21X1 OAI21X1_5 ( .A(i_add2[32]), .B(i_add1[32]), .C(_204_), .Y(_205_) );
INVX1 INVX1_33 ( .A(_205_), .Y(w_C_33_) );
INVX1 INVX1_34 ( .A(i_add2[33]), .Y(_206_) );
INVX1 INVX1_35 ( .A(i_add1[33]), .Y(_207_) );
NOR2X1 NOR2X1_13 ( .A(_206_), .B(_207_), .Y(_208_) );
INVX1 INVX1_36 ( .A(_208_), .Y(_209_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_210_) );
INVX1 INVX1_37 ( .A(_210_), .Y(_211_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_212_) );
INVX1 INVX1_38 ( .A(_212_), .Y(_213_) );
NAND3X1 NAND3X1_10 ( .A(_211_), .B(_213_), .C(_204_), .Y(_214_) );
AND2X2 AND2X2_9 ( .A(_214_), .B(_209_), .Y(_215_) );
INVX1 INVX1_39 ( .A(_215_), .Y(w_C_34_) );
AND2X2 AND2X2_10 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_216_) );
INVX1 INVX1_40 ( .A(_216_), .Y(_217_) );
NAND3X1 NAND3X1_11 ( .A(_209_), .B(_217_), .C(_214_), .Y(_218_) );
OAI21X1 OAI21X1_6 ( .A(i_add2[34]), .B(i_add1[34]), .C(_218_), .Y(_219_) );
INVX1 INVX1_41 ( .A(_219_), .Y(w_C_35_) );
INVX1 INVX1_42 ( .A(i_add2[35]), .Y(_220_) );
INVX1 INVX1_43 ( .A(i_add1[35]), .Y(_221_) );
NOR2X1 NOR2X1_16 ( .A(_220_), .B(_221_), .Y(_222_) );
INVX1 INVX1_44 ( .A(_222_), .Y(_223_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_224_) );
INVX1 INVX1_45 ( .A(_224_), .Y(_225_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_226_) );
INVX1 INVX1_46 ( .A(_226_), .Y(_227_) );
NAND3X1 NAND3X1_12 ( .A(_225_), .B(_227_), .C(_218_), .Y(_228_) );
AND2X2 AND2X2_11 ( .A(_228_), .B(_223_), .Y(_229_) );
INVX1 INVX1_47 ( .A(_229_), .Y(w_C_36_) );
AND2X2 AND2X2_12 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_230_) );
INVX1 INVX1_48 ( .A(_230_), .Y(_231_) );
NAND3X1 NAND3X1_13 ( .A(_223_), .B(_231_), .C(_228_), .Y(_232_) );
OAI21X1 OAI21X1_7 ( .A(i_add2[36]), .B(i_add1[36]), .C(_232_), .Y(_233_) );
INVX1 INVX1_49 ( .A(_233_), .Y(w_C_37_) );
INVX1 INVX1_50 ( .A(i_add2[37]), .Y(_234_) );
INVX1 INVX1_51 ( .A(i_add1[37]), .Y(_235_) );
NOR2X1 NOR2X1_19 ( .A(_234_), .B(_235_), .Y(_236_) );
INVX1 INVX1_52 ( .A(_236_), .Y(_237_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_238_) );
INVX1 INVX1_53 ( .A(_238_), .Y(_239_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_240_) );
INVX1 INVX1_54 ( .A(_240_), .Y(_241_) );
NAND3X1 NAND3X1_14 ( .A(_239_), .B(_241_), .C(_232_), .Y(_242_) );
AND2X2 AND2X2_13 ( .A(_242_), .B(_237_), .Y(_243_) );
INVX1 INVX1_55 ( .A(_243_), .Y(w_C_38_) );
AND2X2 AND2X2_14 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_244_) );
INVX1 INVX1_56 ( .A(_244_), .Y(_245_) );
NAND3X1 NAND3X1_15 ( .A(_237_), .B(_245_), .C(_242_), .Y(_246_) );
OAI21X1 OAI21X1_8 ( .A(i_add2[38]), .B(i_add1[38]), .C(_246_), .Y(_247_) );
INVX1 INVX1_57 ( .A(_247_), .Y(w_C_39_) );
INVX1 INVX1_58 ( .A(i_add2[39]), .Y(_248_) );
INVX1 INVX1_59 ( .A(i_add1[39]), .Y(_249_) );
NOR2X1 NOR2X1_22 ( .A(_248_), .B(_249_), .Y(_250_) );
INVX1 INVX1_60 ( .A(_250_), .Y(_251_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_252_) );
INVX1 INVX1_61 ( .A(_252_), .Y(_253_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_254_) );
INVX1 INVX1_62 ( .A(_254_), .Y(_255_) );
NAND3X1 NAND3X1_16 ( .A(_253_), .B(_255_), .C(_246_), .Y(_256_) );
AND2X2 AND2X2_15 ( .A(_256_), .B(_251_), .Y(_257_) );
INVX1 INVX1_63 ( .A(_257_), .Y(w_C_40_) );
AND2X2 AND2X2_16 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_258_) );
INVX1 INVX1_64 ( .A(_258_), .Y(_259_) );
NAND3X1 NAND3X1_17 ( .A(_251_), .B(_259_), .C(_256_), .Y(_260_) );
OAI21X1 OAI21X1_9 ( .A(i_add2[40]), .B(i_add1[40]), .C(_260_), .Y(_261_) );
INVX1 INVX1_65 ( .A(_261_), .Y(w_C_41_) );
INVX1 INVX1_66 ( .A(i_add2[41]), .Y(_262_) );
INVX1 INVX1_67 ( .A(i_add1[41]), .Y(_263_) );
NOR2X1 NOR2X1_25 ( .A(_262_), .B(_263_), .Y(_264_) );
INVX1 INVX1_68 ( .A(_264_), .Y(_265_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_266_) );
INVX1 INVX1_69 ( .A(_266_), .Y(_267_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_268_) );
INVX1 INVX1_70 ( .A(_268_), .Y(_269_) );
NAND3X1 NAND3X1_18 ( .A(_267_), .B(_269_), .C(_260_), .Y(_270_) );
AND2X2 AND2X2_17 ( .A(_270_), .B(_265_), .Y(_271_) );
INVX1 INVX1_71 ( .A(_271_), .Y(w_C_42_) );
AND2X2 AND2X2_18 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_272_) );
INVX1 INVX1_72 ( .A(_272_), .Y(_273_) );
NAND3X1 NAND3X1_19 ( .A(_265_), .B(_273_), .C(_270_), .Y(_274_) );
OAI21X1 OAI21X1_10 ( .A(i_add2[42]), .B(i_add1[42]), .C(_274_), .Y(_275_) );
INVX1 INVX1_73 ( .A(_275_), .Y(w_C_43_) );
INVX1 INVX1_74 ( .A(i_add2[43]), .Y(_276_) );
INVX1 INVX1_75 ( .A(i_add1[43]), .Y(_277_) );
NOR2X1 NOR2X1_28 ( .A(_276_), .B(_277_), .Y(_278_) );
INVX1 INVX1_76 ( .A(_278_), .Y(_279_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_280_) );
INVX1 INVX1_77 ( .A(_280_), .Y(_281_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_282_) );
INVX1 INVX1_78 ( .A(_282_), .Y(_283_) );
NAND3X1 NAND3X1_20 ( .A(_281_), .B(_283_), .C(_274_), .Y(_284_) );
AND2X2 AND2X2_19 ( .A(_284_), .B(_279_), .Y(_285_) );
INVX1 INVX1_79 ( .A(_285_), .Y(w_C_44_) );
AND2X2 AND2X2_20 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_286_) );
INVX1 INVX1_80 ( .A(_286_), .Y(_287_) );
NAND3X1 NAND3X1_21 ( .A(_279_), .B(_287_), .C(_284_), .Y(_288_) );
OAI21X1 OAI21X1_11 ( .A(i_add2[44]), .B(i_add1[44]), .C(_288_), .Y(_289_) );
INVX1 INVX1_81 ( .A(_289_), .Y(w_C_45_) );
INVX1 INVX1_82 ( .A(i_add2[45]), .Y(_290_) );
INVX1 INVX1_83 ( .A(i_add1[45]), .Y(_291_) );
NOR2X1 NOR2X1_31 ( .A(_290_), .B(_291_), .Y(_292_) );
INVX1 INVX1_84 ( .A(_292_), .Y(_293_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_294_) );
INVX1 INVX1_85 ( .A(_294_), .Y(_295_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_296_) );
INVX1 INVX1_86 ( .A(_296_), .Y(_297_) );
NAND3X1 NAND3X1_22 ( .A(_295_), .B(_297_), .C(_288_), .Y(_298_) );
AND2X2 AND2X2_21 ( .A(_298_), .B(_293_), .Y(_299_) );
INVX1 INVX1_87 ( .A(_299_), .Y(w_C_46_) );
AND2X2 AND2X2_22 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_300_) );
INVX1 INVX1_88 ( .A(_300_), .Y(_301_) );
NAND3X1 NAND3X1_23 ( .A(_293_), .B(_301_), .C(_298_), .Y(_302_) );
OAI21X1 OAI21X1_12 ( .A(i_add2[46]), .B(i_add1[46]), .C(_302_), .Y(_303_) );
INVX1 INVX1_89 ( .A(_303_), .Y(w_C_47_) );
INVX1 INVX1_90 ( .A(i_add2[47]), .Y(_304_) );
INVX1 INVX1_91 ( .A(i_add1[47]), .Y(_305_) );
NOR2X1 NOR2X1_34 ( .A(_304_), .B(_305_), .Y(_306_) );
INVX1 INVX1_92 ( .A(_306_), .Y(_307_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_308_) );
INVX1 INVX1_93 ( .A(_308_), .Y(_309_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_310_) );
INVX1 INVX1_94 ( .A(_310_), .Y(_311_) );
NAND3X1 NAND3X1_24 ( .A(_309_), .B(_311_), .C(_302_), .Y(_312_) );
AND2X2 AND2X2_23 ( .A(_312_), .B(_307_), .Y(_313_) );
INVX1 INVX1_95 ( .A(_313_), .Y(w_C_48_) );
AND2X2 AND2X2_24 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_314_) );
INVX1 INVX1_96 ( .A(_314_), .Y(_315_) );
NAND3X1 NAND3X1_25 ( .A(_307_), .B(_315_), .C(_312_), .Y(_316_) );
OAI21X1 OAI21X1_13 ( .A(i_add2[48]), .B(i_add1[48]), .C(_316_), .Y(_317_) );
INVX1 INVX1_97 ( .A(_317_), .Y(w_C_49_) );
INVX1 INVX1_98 ( .A(i_add2[49]), .Y(_318_) );
INVX1 INVX1_99 ( .A(i_add1[49]), .Y(_319_) );
NOR2X1 NOR2X1_37 ( .A(_318_), .B(_319_), .Y(_320_) );
INVX1 INVX1_100 ( .A(_320_), .Y(_321_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_322_) );
INVX1 INVX1_101 ( .A(_322_), .Y(_323_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_324_) );
INVX1 INVX1_102 ( .A(_324_), .Y(_325_) );
NAND3X1 NAND3X1_26 ( .A(_323_), .B(_325_), .C(_316_), .Y(_326_) );
AND2X2 AND2X2_25 ( .A(_326_), .B(_321_), .Y(_327_) );
INVX1 INVX1_103 ( .A(_327_), .Y(w_C_50_) );
AND2X2 AND2X2_26 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_328_) );
INVX1 INVX1_104 ( .A(_328_), .Y(_329_) );
NAND3X1 NAND3X1_27 ( .A(_321_), .B(_329_), .C(_326_), .Y(_330_) );
OAI21X1 OAI21X1_14 ( .A(i_add2[50]), .B(i_add1[50]), .C(_330_), .Y(_331_) );
INVX1 INVX1_105 ( .A(_331_), .Y(w_C_51_) );
NAND2X1 NAND2X1_1 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_332_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_333_) );
OAI21X1 OAI21X1_15 ( .A(_333_), .B(_331_), .C(_332_), .Y(w_C_52_) );
OR2X2 OR2X2_1 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_334_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_335_) );
INVX1 INVX1_106 ( .A(_335_), .Y(_336_) );
INVX1 INVX1_107 ( .A(_333_), .Y(_337_) );
NAND3X1 NAND3X1_28 ( .A(_336_), .B(_337_), .C(_330_), .Y(_338_) );
NAND2X1 NAND2X1_2 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_339_) );
NAND3X1 NAND3X1_29 ( .A(_332_), .B(_339_), .C(_338_), .Y(_340_) );
AND2X2 AND2X2_27 ( .A(_340_), .B(_334_), .Y(w_C_53_) );
INVX1 INVX1_108 ( .A(i_add2[53]), .Y(_341_) );
INVX1 INVX1_109 ( .A(i_add1[53]), .Y(_342_) );
NAND2X1 NAND2X1_3 ( .A(_341_), .B(_342_), .Y(_343_) );
NAND3X1 NAND3X1_30 ( .A(_334_), .B(_343_), .C(_340_), .Y(_344_) );
OAI21X1 OAI21X1_16 ( .A(_341_), .B(_342_), .C(_344_), .Y(w_C_54_) );
INVX1 INVX1_110 ( .A(i_add2[54]), .Y(_345_) );
INVX1 INVX1_111 ( .A(i_add1[54]), .Y(_346_) );
NAND2X1 NAND2X1_4 ( .A(_345_), .B(_346_), .Y(_347_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_348_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_349_) );
NAND3X1 NAND3X1_31 ( .A(_348_), .B(_349_), .C(_344_), .Y(_350_) );
AND2X2 AND2X2_28 ( .A(_350_), .B(_347_), .Y(w_C_55_) );
INVX1 INVX1_112 ( .A(i_add2[55]), .Y(_351_) );
INVX1 INVX1_113 ( .A(i_add1[55]), .Y(_352_) );
NAND2X1 NAND2X1_7 ( .A(_351_), .B(_352_), .Y(_353_) );
NAND3X1 NAND3X1_32 ( .A(_347_), .B(_353_), .C(_350_), .Y(_354_) );
OAI21X1 OAI21X1_17 ( .A(_351_), .B(_352_), .C(_354_), .Y(w_C_56_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_355_) );
INVX1 INVX1_114 ( .A(_355_), .Y(_356_) );
NOR2X1 NOR2X1_43 ( .A(_351_), .B(_352_), .Y(_357_) );
INVX1 INVX1_115 ( .A(_357_), .Y(_358_) );
INVX1 INVX1_116 ( .A(i_add2[56]), .Y(_359_) );
INVX1 INVX1_117 ( .A(i_add1[56]), .Y(_360_) );
NOR2X1 NOR2X1_44 ( .A(_359_), .B(_360_), .Y(_361_) );
INVX1 INVX1_118 ( .A(_361_), .Y(_362_) );
NAND3X1 NAND3X1_33 ( .A(_358_), .B(_362_), .C(_354_), .Y(_363_) );
AND2X2 AND2X2_29 ( .A(_363_), .B(_356_), .Y(w_C_57_) );
INVX1 INVX1_119 ( .A(i_add2[57]), .Y(_364_) );
INVX1 INVX1_120 ( .A(i_add1[57]), .Y(_365_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_366_) );
INVX1 INVX1_121 ( .A(_366_), .Y(_367_) );
NAND3X1 NAND3X1_34 ( .A(_356_), .B(_367_), .C(_363_), .Y(_368_) );
OAI21X1 OAI21X1_18 ( .A(_364_), .B(_365_), .C(_368_), .Y(w_C_58_) );
INVX1 INVX1_122 ( .A(i_add2[58]), .Y(_369_) );
INVX1 INVX1_123 ( .A(i_add1[58]), .Y(_370_) );
OAI21X1 OAI21X1_19 ( .A(i_add2[58]), .B(i_add1[58]), .C(w_C_58_), .Y(_371_) );
OAI21X1 OAI21X1_20 ( .A(_369_), .B(_370_), .C(_371_), .Y(w_C_59_) );
NOR2X1 NOR2X1_46 ( .A(_369_), .B(_370_), .Y(_372_) );
INVX1 INVX1_124 ( .A(_372_), .Y(_373_) );
AND2X2 AND2X2_30 ( .A(i_add2[59]), .B(i_add1[59]), .Y(_374_) );
INVX1 INVX1_125 ( .A(_374_), .Y(_375_) );
NAND3X1 NAND3X1_35 ( .A(_373_), .B(_375_), .C(_371_), .Y(_376_) );
OAI21X1 OAI21X1_21 ( .A(i_add2[59]), .B(i_add1[59]), .C(_376_), .Y(_377_) );
INVX1 INVX1_126 ( .A(_377_), .Y(w_C_60_) );
NAND2X1 NAND2X1_8 ( .A(i_add2[60]), .B(i_add1[60]), .Y(_378_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[60]), .B(i_add1[60]), .Y(_379_) );
OAI21X1 OAI21X1_22 ( .A(_379_), .B(_377_), .C(_378_), .Y(w_C_61_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[61]), .B(i_add1[61]), .Y(_380_) );
INVX1 INVX1_127 ( .A(_379_), .Y(_381_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[58]), .B(i_add1[58]), .Y(_382_) );
INVX1 INVX1_128 ( .A(_382_), .Y(_383_) );
NOR2X1 NOR2X1_49 ( .A(_364_), .B(_365_), .Y(_384_) );
INVX1 INVX1_129 ( .A(_384_), .Y(_385_) );
NAND3X1 NAND3X1_36 ( .A(_385_), .B(_373_), .C(_368_), .Y(_386_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[59]), .B(i_add1[59]), .Y(_387_) );
INVX1 INVX1_130 ( .A(_387_), .Y(_388_) );
NAND3X1 NAND3X1_37 ( .A(_383_), .B(_388_), .C(_386_), .Y(_389_) );
NAND3X1 NAND3X1_38 ( .A(_375_), .B(_378_), .C(_389_), .Y(_390_) );
OR2X2 OR2X2_2 ( .A(i_add2[61]), .B(i_add1[61]), .Y(_391_) );
NAND3X1 NAND3X1_39 ( .A(_381_), .B(_391_), .C(_390_), .Y(_392_) );
NAND2X1 NAND2X1_10 ( .A(_380_), .B(_392_), .Y(w_C_62_) );
OR2X2 OR2X2_3 ( .A(i_add2[62]), .B(i_add1[62]), .Y(_393_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[62]), .B(i_add1[62]), .Y(_394_) );
NAND3X1 NAND3X1_40 ( .A(_380_), .B(_394_), .C(_392_), .Y(_395_) );
AND2X2 AND2X2_31 ( .A(_395_), .B(_393_), .Y(w_C_63_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[63]), .B(i_add1[63]), .Y(_396_) );
OR2X2 OR2X2_4 ( .A(i_add2[63]), .B(i_add1[63]), .Y(_397_) );
NAND3X1 NAND3X1_41 ( .A(_393_), .B(_397_), .C(_395_), .Y(_398_) );
NAND2X1 NAND2X1_13 ( .A(_396_), .B(_398_), .Y(w_C_64_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_131 ( .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_52 ( .A(_1_), .B(_2_), .Y(w_C_2_) );
INVX1 INVX1_132 ( .A(i_add2[2]), .Y(_3_) );
INVX1 INVX1_133 ( .A(i_add1[2]), .Y(_4_) );
NAND2X1 NAND2X1_15 ( .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
OAI21X1 OAI21X1_23 ( .A(_1_), .B(_2_), .C(_6_), .Y(_7_) );
AND2X2 AND2X2_32 ( .A(_7_), .B(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
OR2X2 OR2X2_5 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_42 ( .A(_5_), .B(_9_), .C(_7_), .Y(_10_) );
NAND2X1 NAND2X1_18 ( .A(_8_), .B(_10_), .Y(w_C_4_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
NAND3X1 NAND3X1_43 ( .A(_8_), .B(_11_), .C(_10_), .Y(_12_) );
OAI21X1 OAI21X1_24 ( .A(i_add2[4]), .B(i_add1[4]), .C(_12_), .Y(_13_) );
INVX1 INVX1_134 ( .A(_13_), .Y(w_C_5_) );
INVX1 INVX1_135 ( .A(i_add2[5]), .Y(_14_) );
BUFX2 BUFX2_1 ( .A(_399__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_399__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_399__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_399__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_399__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_399__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_399__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_399__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_399__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_399__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_399__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_399__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_399__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_399__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_399__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_399__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_399__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_399__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_399__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_399__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_399__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_399__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_399__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_399__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_399__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_399__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_399__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_399__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_399__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_399__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_399__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_399__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_399__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_399__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_399__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_399__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_399__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(_399__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .A(_399__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .A(_399__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .A(_399__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .A(_399__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .A(_399__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .A(_399__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .A(_399__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .A(_399__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .A(_399__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .A(_399__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .A(_399__48_), .Y(o_result[48]) );
BUFX2 BUFX2_50 ( .A(_399__49_), .Y(o_result[49]) );
BUFX2 BUFX2_51 ( .A(_399__50_), .Y(o_result[50]) );
BUFX2 BUFX2_52 ( .A(_399__51_), .Y(o_result[51]) );
BUFX2 BUFX2_53 ( .A(_399__52_), .Y(o_result[52]) );
BUFX2 BUFX2_54 ( .A(_399__53_), .Y(o_result[53]) );
BUFX2 BUFX2_55 ( .A(_399__54_), .Y(o_result[54]) );
BUFX2 BUFX2_56 ( .A(_399__55_), .Y(o_result[55]) );
BUFX2 BUFX2_57 ( .A(_399__56_), .Y(o_result[56]) );
BUFX2 BUFX2_58 ( .A(_399__57_), .Y(o_result[57]) );
BUFX2 BUFX2_59 ( .A(_399__58_), .Y(o_result[58]) );
BUFX2 BUFX2_60 ( .A(_399__59_), .Y(o_result[59]) );
BUFX2 BUFX2_61 ( .A(_399__60_), .Y(o_result[60]) );
BUFX2 BUFX2_62 ( .A(_399__61_), .Y(o_result[61]) );
BUFX2 BUFX2_63 ( .A(_399__62_), .Y(o_result[62]) );
BUFX2 BUFX2_64 ( .A(_399__63_), .Y(o_result[63]) );
BUFX2 BUFX2_65 ( .A(w_C_64_), .Y(o_result[64]) );
INVX1 INVX1_136 ( .A(w_C_4_), .Y(_403_) );
OR2X2 OR2X2_6 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_404_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_405_) );
NAND3X1 NAND3X1_44 ( .A(_403_), .B(_405_), .C(_404_), .Y(_406_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_400_) );
AND2X2 AND2X2_33 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_401_) );
OAI21X1 OAI21X1_25 ( .A(_400_), .B(_401_), .C(w_C_4_), .Y(_402_) );
NAND2X1 NAND2X1_21 ( .A(_402_), .B(_406_), .Y(_399__4_) );
INVX1 INVX1_137 ( .A(w_C_5_), .Y(_410_) );
OR2X2 OR2X2_7 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_411_) );
NAND2X1 NAND2X1_22 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_412_) );
NAND3X1 NAND3X1_45 ( .A(_410_), .B(_412_), .C(_411_), .Y(_413_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_407_) );
AND2X2 AND2X2_34 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_408_) );
OAI21X1 OAI21X1_26 ( .A(_407_), .B(_408_), .C(w_C_5_), .Y(_409_) );
NAND2X1 NAND2X1_23 ( .A(_409_), .B(_413_), .Y(_399__5_) );
INVX1 INVX1_138 ( .A(w_C_6_), .Y(_417_) );
OR2X2 OR2X2_8 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_418_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_419_) );
NAND3X1 NAND3X1_46 ( .A(_417_), .B(_419_), .C(_418_), .Y(_420_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_414_) );
AND2X2 AND2X2_35 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_415_) );
OAI21X1 OAI21X1_27 ( .A(_414_), .B(_415_), .C(w_C_6_), .Y(_416_) );
NAND2X1 NAND2X1_25 ( .A(_416_), .B(_420_), .Y(_399__6_) );
INVX1 INVX1_139 ( .A(w_C_7_), .Y(_424_) );
OR2X2 OR2X2_9 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_425_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_426_) );
NAND3X1 NAND3X1_47 ( .A(_424_), .B(_426_), .C(_425_), .Y(_427_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_421_) );
AND2X2 AND2X2_36 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_422_) );
OAI21X1 OAI21X1_28 ( .A(_421_), .B(_422_), .C(w_C_7_), .Y(_423_) );
NAND2X1 NAND2X1_27 ( .A(_423_), .B(_427_), .Y(_399__7_) );
INVX1 INVX1_140 ( .A(w_C_8_), .Y(_431_) );
OR2X2 OR2X2_10 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_432_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_433_) );
NAND3X1 NAND3X1_48 ( .A(_431_), .B(_433_), .C(_432_), .Y(_434_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_428_) );
AND2X2 AND2X2_37 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_429_) );
OAI21X1 OAI21X1_29 ( .A(_428_), .B(_429_), .C(w_C_8_), .Y(_430_) );
NAND2X1 NAND2X1_29 ( .A(_430_), .B(_434_), .Y(_399__8_) );
INVX1 INVX1_141 ( .A(w_C_9_), .Y(_438_) );
OR2X2 OR2X2_11 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_439_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_440_) );
NAND3X1 NAND3X1_49 ( .A(_438_), .B(_440_), .C(_439_), .Y(_441_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_435_) );
AND2X2 AND2X2_38 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_436_) );
OAI21X1 OAI21X1_30 ( .A(_435_), .B(_436_), .C(w_C_9_), .Y(_437_) );
NAND2X1 NAND2X1_31 ( .A(_437_), .B(_441_), .Y(_399__9_) );
INVX1 INVX1_142 ( .A(w_C_10_), .Y(_445_) );
OR2X2 OR2X2_12 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_446_) );
NAND2X1 NAND2X1_32 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_447_) );
NAND3X1 NAND3X1_50 ( .A(_445_), .B(_447_), .C(_446_), .Y(_448_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_442_) );
AND2X2 AND2X2_39 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_443_) );
OAI21X1 OAI21X1_31 ( .A(_442_), .B(_443_), .C(w_C_10_), .Y(_444_) );
NAND2X1 NAND2X1_33 ( .A(_444_), .B(_448_), .Y(_399__10_) );
INVX1 INVX1_143 ( .A(w_C_11_), .Y(_452_) );
OR2X2 OR2X2_13 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_453_) );
NAND2X1 NAND2X1_34 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_454_) );
NAND3X1 NAND3X1_51 ( .A(_452_), .B(_454_), .C(_453_), .Y(_455_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_449_) );
AND2X2 AND2X2_40 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_450_) );
OAI21X1 OAI21X1_32 ( .A(_449_), .B(_450_), .C(w_C_11_), .Y(_451_) );
NAND2X1 NAND2X1_35 ( .A(_451_), .B(_455_), .Y(_399__11_) );
INVX1 INVX1_144 ( .A(w_C_12_), .Y(_459_) );
OR2X2 OR2X2_14 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_460_) );
NAND2X1 NAND2X1_36 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_461_) );
NAND3X1 NAND3X1_52 ( .A(_459_), .B(_461_), .C(_460_), .Y(_462_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_456_) );
AND2X2 AND2X2_41 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_457_) );
OAI21X1 OAI21X1_33 ( .A(_456_), .B(_457_), .C(w_C_12_), .Y(_458_) );
NAND2X1 NAND2X1_37 ( .A(_458_), .B(_462_), .Y(_399__12_) );
INVX1 INVX1_145 ( .A(w_C_13_), .Y(_466_) );
OR2X2 OR2X2_15 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_467_) );
NAND2X1 NAND2X1_38 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_468_) );
NAND3X1 NAND3X1_53 ( .A(_466_), .B(_468_), .C(_467_), .Y(_469_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_463_) );
AND2X2 AND2X2_42 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_464_) );
OAI21X1 OAI21X1_34 ( .A(_463_), .B(_464_), .C(w_C_13_), .Y(_465_) );
NAND2X1 NAND2X1_39 ( .A(_465_), .B(_469_), .Y(_399__13_) );
INVX1 INVX1_146 ( .A(w_C_14_), .Y(_473_) );
OR2X2 OR2X2_16 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_474_) );
NAND2X1 NAND2X1_40 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_475_) );
NAND3X1 NAND3X1_54 ( .A(_473_), .B(_475_), .C(_474_), .Y(_476_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_470_) );
AND2X2 AND2X2_43 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_471_) );
OAI21X1 OAI21X1_35 ( .A(_470_), .B(_471_), .C(w_C_14_), .Y(_472_) );
NAND2X1 NAND2X1_41 ( .A(_472_), .B(_476_), .Y(_399__14_) );
INVX1 INVX1_147 ( .A(w_C_15_), .Y(_480_) );
OR2X2 OR2X2_17 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_481_) );
NAND2X1 NAND2X1_42 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_482_) );
NAND3X1 NAND3X1_55 ( .A(_480_), .B(_482_), .C(_481_), .Y(_483_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_477_) );
AND2X2 AND2X2_44 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_478_) );
OAI21X1 OAI21X1_36 ( .A(_477_), .B(_478_), .C(w_C_15_), .Y(_479_) );
NAND2X1 NAND2X1_43 ( .A(_479_), .B(_483_), .Y(_399__15_) );
INVX1 INVX1_148 ( .A(w_C_16_), .Y(_487_) );
OR2X2 OR2X2_18 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_488_) );
NAND2X1 NAND2X1_44 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_489_) );
NAND3X1 NAND3X1_56 ( .A(_487_), .B(_489_), .C(_488_), .Y(_490_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_484_) );
AND2X2 AND2X2_45 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_485_) );
OAI21X1 OAI21X1_37 ( .A(_484_), .B(_485_), .C(w_C_16_), .Y(_486_) );
NAND2X1 NAND2X1_45 ( .A(_486_), .B(_490_), .Y(_399__16_) );
INVX1 INVX1_149 ( .A(w_C_17_), .Y(_494_) );
OR2X2 OR2X2_19 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_495_) );
NAND2X1 NAND2X1_46 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_496_) );
NAND3X1 NAND3X1_57 ( .A(_494_), .B(_496_), .C(_495_), .Y(_497_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_491_) );
AND2X2 AND2X2_46 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_492_) );
OAI21X1 OAI21X1_38 ( .A(_491_), .B(_492_), .C(w_C_17_), .Y(_493_) );
NAND2X1 NAND2X1_47 ( .A(_493_), .B(_497_), .Y(_399__17_) );
INVX1 INVX1_150 ( .A(w_C_18_), .Y(_501_) );
OR2X2 OR2X2_20 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_502_) );
NAND2X1 NAND2X1_48 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_503_) );
NAND3X1 NAND3X1_58 ( .A(_501_), .B(_503_), .C(_502_), .Y(_504_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_498_) );
AND2X2 AND2X2_47 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_499_) );
OAI21X1 OAI21X1_39 ( .A(_498_), .B(_499_), .C(w_C_18_), .Y(_500_) );
NAND2X1 NAND2X1_49 ( .A(_500_), .B(_504_), .Y(_399__18_) );
INVX1 INVX1_151 ( .A(w_C_19_), .Y(_508_) );
OR2X2 OR2X2_21 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_509_) );
NAND2X1 NAND2X1_50 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_510_) );
NAND3X1 NAND3X1_59 ( .A(_508_), .B(_510_), .C(_509_), .Y(_511_) );
NOR2X1 NOR2X1_68 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_505_) );
AND2X2 AND2X2_48 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_506_) );
OAI21X1 OAI21X1_40 ( .A(_505_), .B(_506_), .C(w_C_19_), .Y(_507_) );
NAND2X1 NAND2X1_51 ( .A(_507_), .B(_511_), .Y(_399__19_) );
INVX1 INVX1_152 ( .A(w_C_20_), .Y(_515_) );
OR2X2 OR2X2_22 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_516_) );
NAND2X1 NAND2X1_52 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_517_) );
NAND3X1 NAND3X1_60 ( .A(_515_), .B(_517_), .C(_516_), .Y(_518_) );
NOR2X1 NOR2X1_69 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_512_) );
AND2X2 AND2X2_49 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_513_) );
OAI21X1 OAI21X1_41 ( .A(_512_), .B(_513_), .C(w_C_20_), .Y(_514_) );
NAND2X1 NAND2X1_53 ( .A(_514_), .B(_518_), .Y(_399__20_) );
INVX1 INVX1_153 ( .A(w_C_21_), .Y(_522_) );
OR2X2 OR2X2_23 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_523_) );
NAND2X1 NAND2X1_54 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_524_) );
NAND3X1 NAND3X1_61 ( .A(_522_), .B(_524_), .C(_523_), .Y(_525_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_519_) );
AND2X2 AND2X2_50 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_520_) );
OAI21X1 OAI21X1_42 ( .A(_519_), .B(_520_), .C(w_C_21_), .Y(_521_) );
NAND2X1 NAND2X1_55 ( .A(_521_), .B(_525_), .Y(_399__21_) );
INVX1 INVX1_154 ( .A(w_C_22_), .Y(_529_) );
OR2X2 OR2X2_24 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_530_) );
NAND2X1 NAND2X1_56 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_531_) );
NAND3X1 NAND3X1_62 ( .A(_529_), .B(_531_), .C(_530_), .Y(_532_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_526_) );
AND2X2 AND2X2_51 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_527_) );
OAI21X1 OAI21X1_43 ( .A(_526_), .B(_527_), .C(w_C_22_), .Y(_528_) );
NAND2X1 NAND2X1_57 ( .A(_528_), .B(_532_), .Y(_399__22_) );
INVX1 INVX1_155 ( .A(w_C_23_), .Y(_536_) );
OR2X2 OR2X2_25 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_537_) );
NAND2X1 NAND2X1_58 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_538_) );
NAND3X1 NAND3X1_63 ( .A(_536_), .B(_538_), .C(_537_), .Y(_539_) );
NOR2X1 NOR2X1_72 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_533_) );
AND2X2 AND2X2_52 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_534_) );
OAI21X1 OAI21X1_44 ( .A(_533_), .B(_534_), .C(w_C_23_), .Y(_535_) );
NAND2X1 NAND2X1_59 ( .A(_535_), .B(_539_), .Y(_399__23_) );
INVX1 INVX1_156 ( .A(w_C_24_), .Y(_543_) );
OR2X2 OR2X2_26 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_544_) );
NAND2X1 NAND2X1_60 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_545_) );
NAND3X1 NAND3X1_64 ( .A(_543_), .B(_545_), .C(_544_), .Y(_546_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_540_) );
AND2X2 AND2X2_53 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_541_) );
OAI21X1 OAI21X1_45 ( .A(_540_), .B(_541_), .C(w_C_24_), .Y(_542_) );
NAND2X1 NAND2X1_61 ( .A(_542_), .B(_546_), .Y(_399__24_) );
INVX1 INVX1_157 ( .A(w_C_25_), .Y(_550_) );
OR2X2 OR2X2_27 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_551_) );
NAND2X1 NAND2X1_62 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_552_) );
NAND3X1 NAND3X1_65 ( .A(_550_), .B(_552_), .C(_551_), .Y(_553_) );
NOR2X1 NOR2X1_74 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_547_) );
AND2X2 AND2X2_54 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_548_) );
OAI21X1 OAI21X1_46 ( .A(_547_), .B(_548_), .C(w_C_25_), .Y(_549_) );
NAND2X1 NAND2X1_63 ( .A(_549_), .B(_553_), .Y(_399__25_) );
INVX1 INVX1_158 ( .A(w_C_26_), .Y(_557_) );
OR2X2 OR2X2_28 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_558_) );
NAND2X1 NAND2X1_64 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_559_) );
NAND3X1 NAND3X1_66 ( .A(_557_), .B(_559_), .C(_558_), .Y(_560_) );
NOR2X1 NOR2X1_75 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_554_) );
AND2X2 AND2X2_55 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_555_) );
OAI21X1 OAI21X1_47 ( .A(_554_), .B(_555_), .C(w_C_26_), .Y(_556_) );
NAND2X1 NAND2X1_65 ( .A(_556_), .B(_560_), .Y(_399__26_) );
INVX1 INVX1_159 ( .A(w_C_27_), .Y(_564_) );
OR2X2 OR2X2_29 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_565_) );
NAND2X1 NAND2X1_66 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_566_) );
NAND3X1 NAND3X1_67 ( .A(_564_), .B(_566_), .C(_565_), .Y(_567_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_561_) );
AND2X2 AND2X2_56 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_562_) );
OAI21X1 OAI21X1_48 ( .A(_561_), .B(_562_), .C(w_C_27_), .Y(_563_) );
NAND2X1 NAND2X1_67 ( .A(_563_), .B(_567_), .Y(_399__27_) );
INVX1 INVX1_160 ( .A(w_C_28_), .Y(_571_) );
OR2X2 OR2X2_30 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_572_) );
NAND2X1 NAND2X1_68 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_573_) );
NAND3X1 NAND3X1_68 ( .A(_571_), .B(_573_), .C(_572_), .Y(_574_) );
NOR2X1 NOR2X1_77 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_568_) );
AND2X2 AND2X2_57 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_569_) );
OAI21X1 OAI21X1_49 ( .A(_568_), .B(_569_), .C(w_C_28_), .Y(_570_) );
NAND2X1 NAND2X1_69 ( .A(_570_), .B(_574_), .Y(_399__28_) );
INVX1 INVX1_161 ( .A(w_C_29_), .Y(_578_) );
OR2X2 OR2X2_31 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_579_) );
NAND2X1 NAND2X1_70 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_580_) );
NAND3X1 NAND3X1_69 ( .A(_578_), .B(_580_), .C(_579_), .Y(_581_) );
NOR2X1 NOR2X1_78 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_575_) );
AND2X2 AND2X2_58 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_576_) );
OAI21X1 OAI21X1_50 ( .A(_575_), .B(_576_), .C(w_C_29_), .Y(_577_) );
NAND2X1 NAND2X1_71 ( .A(_577_), .B(_581_), .Y(_399__29_) );
INVX1 INVX1_162 ( .A(w_C_30_), .Y(_585_) );
OR2X2 OR2X2_32 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_586_) );
NAND2X1 NAND2X1_72 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_587_) );
NAND3X1 NAND3X1_70 ( .A(_585_), .B(_587_), .C(_586_), .Y(_588_) );
NOR2X1 NOR2X1_79 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_582_) );
AND2X2 AND2X2_59 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_583_) );
OAI21X1 OAI21X1_51 ( .A(_582_), .B(_583_), .C(w_C_30_), .Y(_584_) );
NAND2X1 NAND2X1_73 ( .A(_584_), .B(_588_), .Y(_399__30_) );
INVX1 INVX1_163 ( .A(w_C_31_), .Y(_592_) );
OR2X2 OR2X2_33 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_593_) );
NAND2X1 NAND2X1_74 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_594_) );
NAND3X1 NAND3X1_71 ( .A(_592_), .B(_594_), .C(_593_), .Y(_595_) );
NOR2X1 NOR2X1_80 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_589_) );
AND2X2 AND2X2_60 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_590_) );
OAI21X1 OAI21X1_52 ( .A(_589_), .B(_590_), .C(w_C_31_), .Y(_591_) );
NAND2X1 NAND2X1_75 ( .A(_591_), .B(_595_), .Y(_399__31_) );
INVX1 INVX1_164 ( .A(w_C_32_), .Y(_599_) );
OR2X2 OR2X2_34 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_600_) );
NAND2X1 NAND2X1_76 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_601_) );
NAND3X1 NAND3X1_72 ( .A(_599_), .B(_601_), .C(_600_), .Y(_602_) );
NOR2X1 NOR2X1_81 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_596_) );
AND2X2 AND2X2_61 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_597_) );
OAI21X1 OAI21X1_53 ( .A(_596_), .B(_597_), .C(w_C_32_), .Y(_598_) );
NAND2X1 NAND2X1_77 ( .A(_598_), .B(_602_), .Y(_399__32_) );
INVX1 INVX1_165 ( .A(w_C_33_), .Y(_606_) );
OR2X2 OR2X2_35 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_607_) );
NAND2X1 NAND2X1_78 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_608_) );
NAND3X1 NAND3X1_73 ( .A(_606_), .B(_608_), .C(_607_), .Y(_609_) );
NOR2X1 NOR2X1_82 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_603_) );
AND2X2 AND2X2_62 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_604_) );
OAI21X1 OAI21X1_54 ( .A(_603_), .B(_604_), .C(w_C_33_), .Y(_605_) );
NAND2X1 NAND2X1_79 ( .A(_605_), .B(_609_), .Y(_399__33_) );
INVX1 INVX1_166 ( .A(w_C_34_), .Y(_613_) );
OR2X2 OR2X2_36 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_614_) );
NAND2X1 NAND2X1_80 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_615_) );
NAND3X1 NAND3X1_74 ( .A(_613_), .B(_615_), .C(_614_), .Y(_616_) );
NOR2X1 NOR2X1_83 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_610_) );
AND2X2 AND2X2_63 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_611_) );
OAI21X1 OAI21X1_55 ( .A(_610_), .B(_611_), .C(w_C_34_), .Y(_612_) );
NAND2X1 NAND2X1_81 ( .A(_612_), .B(_616_), .Y(_399__34_) );
INVX1 INVX1_167 ( .A(w_C_35_), .Y(_620_) );
OR2X2 OR2X2_37 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_621_) );
NAND2X1 NAND2X1_82 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_622_) );
NAND3X1 NAND3X1_75 ( .A(_620_), .B(_622_), .C(_621_), .Y(_623_) );
NOR2X1 NOR2X1_84 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_617_) );
AND2X2 AND2X2_64 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_618_) );
OAI21X1 OAI21X1_56 ( .A(_617_), .B(_618_), .C(w_C_35_), .Y(_619_) );
NAND2X1 NAND2X1_83 ( .A(_619_), .B(_623_), .Y(_399__35_) );
INVX1 INVX1_168 ( .A(w_C_36_), .Y(_627_) );
OR2X2 OR2X2_38 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_628_) );
NAND2X1 NAND2X1_84 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_629_) );
NAND3X1 NAND3X1_76 ( .A(_627_), .B(_629_), .C(_628_), .Y(_630_) );
NOR2X1 NOR2X1_85 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_624_) );
AND2X2 AND2X2_65 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_625_) );
OAI21X1 OAI21X1_57 ( .A(_624_), .B(_625_), .C(w_C_36_), .Y(_626_) );
NAND2X1 NAND2X1_85 ( .A(_626_), .B(_630_), .Y(_399__36_) );
INVX1 INVX1_169 ( .A(w_C_37_), .Y(_634_) );
OR2X2 OR2X2_39 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_635_) );
NAND2X1 NAND2X1_86 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_636_) );
NAND3X1 NAND3X1_77 ( .A(_634_), .B(_636_), .C(_635_), .Y(_637_) );
NOR2X1 NOR2X1_86 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_631_) );
AND2X2 AND2X2_66 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_632_) );
OAI21X1 OAI21X1_58 ( .A(_631_), .B(_632_), .C(w_C_37_), .Y(_633_) );
NAND2X1 NAND2X1_87 ( .A(_633_), .B(_637_), .Y(_399__37_) );
INVX1 INVX1_170 ( .A(w_C_38_), .Y(_641_) );
OR2X2 OR2X2_40 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_642_) );
NAND2X1 NAND2X1_88 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_643_) );
NAND3X1 NAND3X1_78 ( .A(_641_), .B(_643_), .C(_642_), .Y(_644_) );
NOR2X1 NOR2X1_87 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_638_) );
AND2X2 AND2X2_67 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_639_) );
OAI21X1 OAI21X1_59 ( .A(_638_), .B(_639_), .C(w_C_38_), .Y(_640_) );
NAND2X1 NAND2X1_89 ( .A(_640_), .B(_644_), .Y(_399__38_) );
INVX1 INVX1_171 ( .A(w_C_39_), .Y(_648_) );
OR2X2 OR2X2_41 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_649_) );
NAND2X1 NAND2X1_90 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_650_) );
NAND3X1 NAND3X1_79 ( .A(_648_), .B(_650_), .C(_649_), .Y(_651_) );
NOR2X1 NOR2X1_88 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_645_) );
AND2X2 AND2X2_68 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_646_) );
OAI21X1 OAI21X1_60 ( .A(_645_), .B(_646_), .C(w_C_39_), .Y(_647_) );
NAND2X1 NAND2X1_91 ( .A(_647_), .B(_651_), .Y(_399__39_) );
INVX1 INVX1_172 ( .A(w_C_40_), .Y(_655_) );
OR2X2 OR2X2_42 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_656_) );
NAND2X1 NAND2X1_92 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_657_) );
NAND3X1 NAND3X1_80 ( .A(_655_), .B(_657_), .C(_656_), .Y(_658_) );
NOR2X1 NOR2X1_89 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_652_) );
AND2X2 AND2X2_69 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_653_) );
OAI21X1 OAI21X1_61 ( .A(_652_), .B(_653_), .C(w_C_40_), .Y(_654_) );
NAND2X1 NAND2X1_93 ( .A(_654_), .B(_658_), .Y(_399__40_) );
INVX1 INVX1_173 ( .A(w_C_41_), .Y(_662_) );
OR2X2 OR2X2_43 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_663_) );
NAND2X1 NAND2X1_94 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_664_) );
NAND3X1 NAND3X1_81 ( .A(_662_), .B(_664_), .C(_663_), .Y(_665_) );
NOR2X1 NOR2X1_90 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_659_) );
AND2X2 AND2X2_70 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_660_) );
OAI21X1 OAI21X1_62 ( .A(_659_), .B(_660_), .C(w_C_41_), .Y(_661_) );
NAND2X1 NAND2X1_95 ( .A(_661_), .B(_665_), .Y(_399__41_) );
INVX1 INVX1_174 ( .A(w_C_42_), .Y(_669_) );
OR2X2 OR2X2_44 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_670_) );
NAND2X1 NAND2X1_96 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_671_) );
NAND3X1 NAND3X1_82 ( .A(_669_), .B(_671_), .C(_670_), .Y(_672_) );
NOR2X1 NOR2X1_91 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_666_) );
AND2X2 AND2X2_71 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_667_) );
OAI21X1 OAI21X1_63 ( .A(_666_), .B(_667_), .C(w_C_42_), .Y(_668_) );
NAND2X1 NAND2X1_97 ( .A(_668_), .B(_672_), .Y(_399__42_) );
INVX1 INVX1_175 ( .A(w_C_43_), .Y(_676_) );
OR2X2 OR2X2_45 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_677_) );
NAND2X1 NAND2X1_98 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_678_) );
NAND3X1 NAND3X1_83 ( .A(_676_), .B(_678_), .C(_677_), .Y(_679_) );
NOR2X1 NOR2X1_92 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_673_) );
AND2X2 AND2X2_72 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_674_) );
OAI21X1 OAI21X1_64 ( .A(_673_), .B(_674_), .C(w_C_43_), .Y(_675_) );
NAND2X1 NAND2X1_99 ( .A(_675_), .B(_679_), .Y(_399__43_) );
INVX1 INVX1_176 ( .A(w_C_44_), .Y(_683_) );
OR2X2 OR2X2_46 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_684_) );
NAND2X1 NAND2X1_100 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_685_) );
NAND3X1 NAND3X1_84 ( .A(_683_), .B(_685_), .C(_684_), .Y(_686_) );
NOR2X1 NOR2X1_93 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_680_) );
AND2X2 AND2X2_73 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_681_) );
OAI21X1 OAI21X1_65 ( .A(_680_), .B(_681_), .C(w_C_44_), .Y(_682_) );
NAND2X1 NAND2X1_101 ( .A(_682_), .B(_686_), .Y(_399__44_) );
INVX1 INVX1_177 ( .A(w_C_45_), .Y(_690_) );
OR2X2 OR2X2_47 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_691_) );
NAND2X1 NAND2X1_102 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_692_) );
NAND3X1 NAND3X1_85 ( .A(_690_), .B(_692_), .C(_691_), .Y(_693_) );
NOR2X1 NOR2X1_94 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_687_) );
AND2X2 AND2X2_74 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_688_) );
OAI21X1 OAI21X1_66 ( .A(_687_), .B(_688_), .C(w_C_45_), .Y(_689_) );
NAND2X1 NAND2X1_103 ( .A(_689_), .B(_693_), .Y(_399__45_) );
INVX1 INVX1_178 ( .A(w_C_46_), .Y(_697_) );
OR2X2 OR2X2_48 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_698_) );
NAND2X1 NAND2X1_104 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_699_) );
NAND3X1 NAND3X1_86 ( .A(_697_), .B(_699_), .C(_698_), .Y(_700_) );
NOR2X1 NOR2X1_95 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_694_) );
AND2X2 AND2X2_75 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_695_) );
OAI21X1 OAI21X1_67 ( .A(_694_), .B(_695_), .C(w_C_46_), .Y(_696_) );
NAND2X1 NAND2X1_105 ( .A(_696_), .B(_700_), .Y(_399__46_) );
INVX1 INVX1_179 ( .A(w_C_47_), .Y(_704_) );
OR2X2 OR2X2_49 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_705_) );
NAND2X1 NAND2X1_106 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_706_) );
NAND3X1 NAND3X1_87 ( .A(_704_), .B(_706_), .C(_705_), .Y(_707_) );
NOR2X1 NOR2X1_96 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_701_) );
AND2X2 AND2X2_76 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_702_) );
OAI21X1 OAI21X1_68 ( .A(_701_), .B(_702_), .C(w_C_47_), .Y(_703_) );
NAND2X1 NAND2X1_107 ( .A(_703_), .B(_707_), .Y(_399__47_) );
INVX1 INVX1_180 ( .A(w_C_48_), .Y(_711_) );
OR2X2 OR2X2_50 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_712_) );
NAND2X1 NAND2X1_108 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_713_) );
NAND3X1 NAND3X1_88 ( .A(_711_), .B(_713_), .C(_712_), .Y(_714_) );
NOR2X1 NOR2X1_97 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_708_) );
AND2X2 AND2X2_77 ( .A(i_add2[48]), .B(i_add1[48]), .Y(_709_) );
OAI21X1 OAI21X1_69 ( .A(_708_), .B(_709_), .C(w_C_48_), .Y(_710_) );
NAND2X1 NAND2X1_109 ( .A(_710_), .B(_714_), .Y(_399__48_) );
INVX1 INVX1_181 ( .A(w_C_49_), .Y(_718_) );
OR2X2 OR2X2_51 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_719_) );
NAND2X1 NAND2X1_110 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_720_) );
NAND3X1 NAND3X1_89 ( .A(_718_), .B(_720_), .C(_719_), .Y(_721_) );
NOR2X1 NOR2X1_98 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_715_) );
AND2X2 AND2X2_78 ( .A(i_add2[49]), .B(i_add1[49]), .Y(_716_) );
OAI21X1 OAI21X1_70 ( .A(_715_), .B(_716_), .C(w_C_49_), .Y(_717_) );
NAND2X1 NAND2X1_111 ( .A(_717_), .B(_721_), .Y(_399__49_) );
INVX1 INVX1_182 ( .A(w_C_50_), .Y(_725_) );
OR2X2 OR2X2_52 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_726_) );
NAND2X1 NAND2X1_112 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_727_) );
NAND3X1 NAND3X1_90 ( .A(_725_), .B(_727_), .C(_726_), .Y(_728_) );
NOR2X1 NOR2X1_99 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_722_) );
AND2X2 AND2X2_79 ( .A(i_add2[50]), .B(i_add1[50]), .Y(_723_) );
OAI21X1 OAI21X1_71 ( .A(_722_), .B(_723_), .C(w_C_50_), .Y(_724_) );
NAND2X1 NAND2X1_113 ( .A(_724_), .B(_728_), .Y(_399__50_) );
INVX1 INVX1_183 ( .A(w_C_51_), .Y(_732_) );
OR2X2 OR2X2_53 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_733_) );
NAND2X1 NAND2X1_114 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_734_) );
NAND3X1 NAND3X1_91 ( .A(_732_), .B(_734_), .C(_733_), .Y(_735_) );
NOR2X1 NOR2X1_100 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_729_) );
AND2X2 AND2X2_80 ( .A(i_add2[51]), .B(i_add1[51]), .Y(_730_) );
OAI21X1 OAI21X1_72 ( .A(_729_), .B(_730_), .C(w_C_51_), .Y(_731_) );
NAND2X1 NAND2X1_115 ( .A(_731_), .B(_735_), .Y(_399__51_) );
INVX1 INVX1_184 ( .A(w_C_52_), .Y(_739_) );
OR2X2 OR2X2_54 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_740_) );
NAND2X1 NAND2X1_116 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_741_) );
NAND3X1 NAND3X1_92 ( .A(_739_), .B(_741_), .C(_740_), .Y(_742_) );
NOR2X1 NOR2X1_101 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_736_) );
AND2X2 AND2X2_81 ( .A(i_add2[52]), .B(i_add1[52]), .Y(_737_) );
OAI21X1 OAI21X1_73 ( .A(_736_), .B(_737_), .C(w_C_52_), .Y(_738_) );
NAND2X1 NAND2X1_117 ( .A(_738_), .B(_742_), .Y(_399__52_) );
INVX1 INVX1_185 ( .A(w_C_53_), .Y(_746_) );
OR2X2 OR2X2_55 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_747_) );
NAND2X1 NAND2X1_118 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_748_) );
NAND3X1 NAND3X1_93 ( .A(_746_), .B(_748_), .C(_747_), .Y(_749_) );
NOR2X1 NOR2X1_102 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_743_) );
AND2X2 AND2X2_82 ( .A(i_add2[53]), .B(i_add1[53]), .Y(_744_) );
OAI21X1 OAI21X1_74 ( .A(_743_), .B(_744_), .C(w_C_53_), .Y(_745_) );
NAND2X1 NAND2X1_119 ( .A(_745_), .B(_749_), .Y(_399__53_) );
INVX1 INVX1_186 ( .A(w_C_54_), .Y(_753_) );
OR2X2 OR2X2_56 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_754_) );
NAND2X1 NAND2X1_120 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_755_) );
NAND3X1 NAND3X1_94 ( .A(_753_), .B(_755_), .C(_754_), .Y(_756_) );
NOR2X1 NOR2X1_103 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_750_) );
AND2X2 AND2X2_83 ( .A(i_add2[54]), .B(i_add1[54]), .Y(_751_) );
OAI21X1 OAI21X1_75 ( .A(_750_), .B(_751_), .C(w_C_54_), .Y(_752_) );
NAND2X1 NAND2X1_121 ( .A(_752_), .B(_756_), .Y(_399__54_) );
INVX1 INVX1_187 ( .A(w_C_55_), .Y(_760_) );
OR2X2 OR2X2_57 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_761_) );
NAND2X1 NAND2X1_122 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_762_) );
NAND3X1 NAND3X1_95 ( .A(_760_), .B(_762_), .C(_761_), .Y(_763_) );
NOR2X1 NOR2X1_104 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_757_) );
AND2X2 AND2X2_84 ( .A(i_add2[55]), .B(i_add1[55]), .Y(_758_) );
OAI21X1 OAI21X1_76 ( .A(_757_), .B(_758_), .C(w_C_55_), .Y(_759_) );
NAND2X1 NAND2X1_123 ( .A(_759_), .B(_763_), .Y(_399__55_) );
INVX1 INVX1_188 ( .A(w_C_56_), .Y(_767_) );
OR2X2 OR2X2_58 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_768_) );
NAND2X1 NAND2X1_124 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_769_) );
NAND3X1 NAND3X1_96 ( .A(_767_), .B(_769_), .C(_768_), .Y(_770_) );
NOR2X1 NOR2X1_105 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_764_) );
AND2X2 AND2X2_85 ( .A(i_add2[56]), .B(i_add1[56]), .Y(_765_) );
OAI21X1 OAI21X1_77 ( .A(_764_), .B(_765_), .C(w_C_56_), .Y(_766_) );
NAND2X1 NAND2X1_125 ( .A(_766_), .B(_770_), .Y(_399__56_) );
INVX1 INVX1_189 ( .A(w_C_57_), .Y(_774_) );
OR2X2 OR2X2_59 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_775_) );
NAND2X1 NAND2X1_126 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_776_) );
NAND3X1 NAND3X1_97 ( .A(_774_), .B(_776_), .C(_775_), .Y(_777_) );
NOR2X1 NOR2X1_106 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_771_) );
AND2X2 AND2X2_86 ( .A(i_add2[57]), .B(i_add1[57]), .Y(_772_) );
OAI21X1 OAI21X1_78 ( .A(_771_), .B(_772_), .C(w_C_57_), .Y(_773_) );
NAND2X1 NAND2X1_127 ( .A(_773_), .B(_777_), .Y(_399__57_) );
INVX1 INVX1_190 ( .A(w_C_58_), .Y(_781_) );
OR2X2 OR2X2_60 ( .A(i_add2[58]), .B(i_add1[58]), .Y(_782_) );
NAND2X1 NAND2X1_128 ( .A(i_add2[58]), .B(i_add1[58]), .Y(_783_) );
NAND3X1 NAND3X1_98 ( .A(_781_), .B(_783_), .C(_782_), .Y(_784_) );
NOR2X1 NOR2X1_107 ( .A(i_add2[58]), .B(i_add1[58]), .Y(_778_) );
AND2X2 AND2X2_87 ( .A(i_add2[58]), .B(i_add1[58]), .Y(_779_) );
OAI21X1 OAI21X1_79 ( .A(_778_), .B(_779_), .C(w_C_58_), .Y(_780_) );
NAND2X1 NAND2X1_129 ( .A(_780_), .B(_784_), .Y(_399__58_) );
INVX1 INVX1_191 ( .A(w_C_59_), .Y(_788_) );
OR2X2 OR2X2_61 ( .A(i_add2[59]), .B(i_add1[59]), .Y(_789_) );
NAND2X1 NAND2X1_130 ( .A(i_add2[59]), .B(i_add1[59]), .Y(_790_) );
NAND3X1 NAND3X1_99 ( .A(_788_), .B(_790_), .C(_789_), .Y(_791_) );
NOR2X1 NOR2X1_108 ( .A(i_add2[59]), .B(i_add1[59]), .Y(_785_) );
AND2X2 AND2X2_88 ( .A(i_add2[59]), .B(i_add1[59]), .Y(_786_) );
OAI21X1 OAI21X1_80 ( .A(_785_), .B(_786_), .C(w_C_59_), .Y(_787_) );
NAND2X1 NAND2X1_131 ( .A(_787_), .B(_791_), .Y(_399__59_) );
INVX1 INVX1_192 ( .A(w_C_60_), .Y(_795_) );
OR2X2 OR2X2_62 ( .A(i_add2[60]), .B(i_add1[60]), .Y(_796_) );
NAND2X1 NAND2X1_132 ( .A(i_add2[60]), .B(i_add1[60]), .Y(_797_) );
NAND3X1 NAND3X1_100 ( .A(_795_), .B(_797_), .C(_796_), .Y(_798_) );
NOR2X1 NOR2X1_109 ( .A(i_add2[60]), .B(i_add1[60]), .Y(_792_) );
AND2X2 AND2X2_89 ( .A(i_add2[60]), .B(i_add1[60]), .Y(_793_) );
OAI21X1 OAI21X1_81 ( .A(_792_), .B(_793_), .C(w_C_60_), .Y(_794_) );
NAND2X1 NAND2X1_133 ( .A(_794_), .B(_798_), .Y(_399__60_) );
INVX1 INVX1_193 ( .A(w_C_61_), .Y(_802_) );
OR2X2 OR2X2_63 ( .A(i_add2[61]), .B(i_add1[61]), .Y(_803_) );
NAND2X1 NAND2X1_134 ( .A(i_add2[61]), .B(i_add1[61]), .Y(_804_) );
NAND3X1 NAND3X1_101 ( .A(_802_), .B(_804_), .C(_803_), .Y(_805_) );
NOR2X1 NOR2X1_110 ( .A(i_add2[61]), .B(i_add1[61]), .Y(_799_) );
AND2X2 AND2X2_90 ( .A(i_add2[61]), .B(i_add1[61]), .Y(_800_) );
OAI21X1 OAI21X1_82 ( .A(_799_), .B(_800_), .C(w_C_61_), .Y(_801_) );
NAND2X1 NAND2X1_135 ( .A(_801_), .B(_805_), .Y(_399__61_) );
INVX1 INVX1_194 ( .A(w_C_62_), .Y(_809_) );
OR2X2 OR2X2_64 ( .A(i_add2[62]), .B(i_add1[62]), .Y(_810_) );
NAND2X1 NAND2X1_136 ( .A(i_add2[62]), .B(i_add1[62]), .Y(_811_) );
NAND3X1 NAND3X1_102 ( .A(_809_), .B(_811_), .C(_810_), .Y(_812_) );
NOR2X1 NOR2X1_111 ( .A(i_add2[62]), .B(i_add1[62]), .Y(_806_) );
AND2X2 AND2X2_91 ( .A(i_add2[62]), .B(i_add1[62]), .Y(_807_) );
OAI21X1 OAI21X1_83 ( .A(_806_), .B(_807_), .C(w_C_62_), .Y(_808_) );
NAND2X1 NAND2X1_137 ( .A(_808_), .B(_812_), .Y(_399__62_) );
INVX1 INVX1_195 ( .A(w_C_63_), .Y(_816_) );
OR2X2 OR2X2_65 ( .A(i_add2[63]), .B(i_add1[63]), .Y(_817_) );
NAND2X1 NAND2X1_138 ( .A(i_add2[63]), .B(i_add1[63]), .Y(_818_) );
NAND3X1 NAND3X1_103 ( .A(_816_), .B(_818_), .C(_817_), .Y(_819_) );
NOR2X1 NOR2X1_112 ( .A(i_add2[63]), .B(i_add1[63]), .Y(_813_) );
AND2X2 AND2X2_92 ( .A(i_add2[63]), .B(i_add1[63]), .Y(_814_) );
OAI21X1 OAI21X1_84 ( .A(_813_), .B(_814_), .C(w_C_63_), .Y(_815_) );
NAND2X1 NAND2X1_139 ( .A(_815_), .B(_819_), .Y(_399__63_) );
INVX1 INVX1_196 ( .A(gnd), .Y(_823_) );
OR2X2 OR2X2_66 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_824_) );
NAND2X1 NAND2X1_140 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_825_) );
NAND3X1 NAND3X1_104 ( .A(_823_), .B(_825_), .C(_824_), .Y(_826_) );
NOR2X1 NOR2X1_113 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_820_) );
AND2X2 AND2X2_93 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_821_) );
OAI21X1 OAI21X1_85 ( .A(_820_), .B(_821_), .C(gnd), .Y(_822_) );
NAND2X1 NAND2X1_141 ( .A(_822_), .B(_826_), .Y(_399__0_) );
INVX1 INVX1_197 ( .A(w_C_1_), .Y(_830_) );
OR2X2 OR2X2_67 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_831_) );
NAND2X1 NAND2X1_142 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_832_) );
NAND3X1 NAND3X1_105 ( .A(_830_), .B(_832_), .C(_831_), .Y(_833_) );
NOR2X1 NOR2X1_114 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_827_) );
AND2X2 AND2X2_94 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_828_) );
OAI21X1 OAI21X1_86 ( .A(_827_), .B(_828_), .C(w_C_1_), .Y(_829_) );
NAND2X1 NAND2X1_143 ( .A(_829_), .B(_833_), .Y(_399__1_) );
INVX1 INVX1_198 ( .A(w_C_2_), .Y(_837_) );
OR2X2 OR2X2_68 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_838_) );
NAND2X1 NAND2X1_144 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_839_) );
NAND3X1 NAND3X1_106 ( .A(_837_), .B(_839_), .C(_838_), .Y(_840_) );
NOR2X1 NOR2X1_115 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_834_) );
AND2X2 AND2X2_95 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_835_) );
OAI21X1 OAI21X1_87 ( .A(_834_), .B(_835_), .C(w_C_2_), .Y(_836_) );
NAND2X1 NAND2X1_145 ( .A(_836_), .B(_840_), .Y(_399__2_) );
INVX1 INVX1_199 ( .A(w_C_3_), .Y(_844_) );
OR2X2 OR2X2_69 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_845_) );
NAND2X1 NAND2X1_146 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_846_) );
NAND3X1 NAND3X1_107 ( .A(_844_), .B(_846_), .C(_845_), .Y(_847_) );
NOR2X1 NOR2X1_116 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_841_) );
AND2X2 AND2X2_96 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_842_) );
OAI21X1 OAI21X1_88 ( .A(_841_), .B(_842_), .C(w_C_3_), .Y(_843_) );
NAND2X1 NAND2X1_147 ( .A(_843_), .B(_847_), .Y(_399__3_) );
INVX1 INVX1_200 ( .A(i_add1[5]), .Y(_15_) );
NOR2X1 NOR2X1_117 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_16_) );
INVX1 INVX1_201 ( .A(_16_), .Y(_17_) );
NOR2X1 NOR2X1_118 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_18_) );
INVX1 INVX1_202 ( .A(_18_), .Y(_19_) );
NAND3X1 NAND3X1_108 ( .A(_17_), .B(_19_), .C(_12_), .Y(_20_) );
OAI21X1 OAI21X1_89 ( .A(_14_), .B(_15_), .C(_20_), .Y(w_C_6_) );
NOR2X1 NOR2X1_119 ( .A(_14_), .B(_15_), .Y(_21_) );
INVX1 INVX1_203 ( .A(_21_), .Y(_22_) );
AND2X2 AND2X2_97 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_23_) );
INVX1 INVX1_204 ( .A(_23_), .Y(_24_) );
NAND3X1 NAND3X1_109 ( .A(_22_), .B(_24_), .C(_20_), .Y(_25_) );
OAI21X1 OAI21X1_90 ( .A(i_add2[6]), .B(i_add1[6]), .C(_25_), .Y(_26_) );
INVX1 INVX1_205 ( .A(_26_), .Y(w_C_7_) );
INVX1 INVX1_206 ( .A(i_add2[7]), .Y(_27_) );
INVX1 INVX1_207 ( .A(i_add1[7]), .Y(_28_) );
NOR2X1 NOR2X1_120 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_29_) );
INVX1 INVX1_208 ( .A(_29_), .Y(_30_) );
NOR2X1 NOR2X1_121 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_31_) );
INVX1 INVX1_209 ( .A(_31_), .Y(_32_) );
NAND3X1 NAND3X1_110 ( .A(_30_), .B(_32_), .C(_25_), .Y(_33_) );
OAI21X1 OAI21X1_91 ( .A(_27_), .B(_28_), .C(_33_), .Y(w_C_8_) );
NOR2X1 NOR2X1_122 ( .A(_27_), .B(_28_), .Y(_34_) );
INVX1 INVX1_210 ( .A(_34_), .Y(_35_) );
AND2X2 AND2X2_98 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_36_) );
INVX1 INVX1_211 ( .A(_36_), .Y(_37_) );
NAND3X1 NAND3X1_111 ( .A(_35_), .B(_37_), .C(_33_), .Y(_38_) );
OAI21X1 OAI21X1_92 ( .A(i_add2[8]), .B(i_add1[8]), .C(_38_), .Y(_39_) );
INVX1 INVX1_212 ( .A(_39_), .Y(w_C_9_) );
INVX1 INVX1_213 ( .A(i_add2[9]), .Y(_40_) );
INVX1 INVX1_214 ( .A(i_add1[9]), .Y(_41_) );
NOR2X1 NOR2X1_123 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_42_) );
INVX1 INVX1_215 ( .A(_42_), .Y(_43_) );
NOR2X1 NOR2X1_124 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_44_) );
INVX1 INVX1_216 ( .A(_44_), .Y(_45_) );
NAND3X1 NAND3X1_112 ( .A(_43_), .B(_45_), .C(_38_), .Y(_46_) );
OAI21X1 OAI21X1_93 ( .A(_40_), .B(_41_), .C(_46_), .Y(w_C_10_) );
NOR2X1 NOR2X1_125 ( .A(_40_), .B(_41_), .Y(_47_) );
INVX1 INVX1_217 ( .A(_47_), .Y(_48_) );
AND2X2 AND2X2_99 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_49_) );
INVX1 INVX1_218 ( .A(_49_), .Y(_50_) );
NAND3X1 NAND3X1_113 ( .A(_48_), .B(_50_), .C(_46_), .Y(_51_) );
OAI21X1 OAI21X1_94 ( .A(i_add2[10]), .B(i_add1[10]), .C(_51_), .Y(_52_) );
INVX1 INVX1_219 ( .A(_52_), .Y(w_C_11_) );
INVX1 INVX1_220 ( .A(i_add2[11]), .Y(_53_) );
INVX1 INVX1_221 ( .A(i_add1[11]), .Y(_54_) );
NOR2X1 NOR2X1_126 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_55_) );
INVX1 INVX1_222 ( .A(_55_), .Y(_56_) );
NOR2X1 NOR2X1_127 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_57_) );
INVX1 INVX1_223 ( .A(_57_), .Y(_58_) );
NAND3X1 NAND3X1_114 ( .A(_56_), .B(_58_), .C(_51_), .Y(_59_) );
OAI21X1 OAI21X1_95 ( .A(_53_), .B(_54_), .C(_59_), .Y(w_C_12_) );
NOR2X1 NOR2X1_128 ( .A(_53_), .B(_54_), .Y(_60_) );
INVX1 INVX1_224 ( .A(_60_), .Y(_61_) );
AND2X2 AND2X2_100 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_62_) );
INVX1 INVX1_225 ( .A(_62_), .Y(_63_) );
NAND3X1 NAND3X1_115 ( .A(_61_), .B(_63_), .C(_59_), .Y(_64_) );
OAI21X1 OAI21X1_96 ( .A(i_add2[12]), .B(i_add1[12]), .C(_64_), .Y(_65_) );
INVX1 INVX1_226 ( .A(_65_), .Y(w_C_13_) );
INVX1 INVX1_227 ( .A(i_add2[13]), .Y(_66_) );
INVX1 INVX1_228 ( .A(i_add1[13]), .Y(_67_) );
NOR2X1 NOR2X1_129 ( .A(_66_), .B(_67_), .Y(_68_) );
INVX1 INVX1_229 ( .A(_68_), .Y(_69_) );
NOR2X1 NOR2X1_130 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_70_) );
INVX1 INVX1_230 ( .A(_70_), .Y(_71_) );
NOR2X1 NOR2X1_131 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_72_) );
INVX1 INVX1_231 ( .A(_72_), .Y(_73_) );
NAND3X1 NAND3X1_116 ( .A(_71_), .B(_73_), .C(_64_), .Y(_74_) );
AND2X2 AND2X2_101 ( .A(_74_), .B(_69_), .Y(_75_) );
INVX1 INVX1_232 ( .A(_75_), .Y(w_C_14_) );
AND2X2 AND2X2_102 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_76_) );
INVX1 INVX1_233 ( .A(_76_), .Y(_77_) );
NAND3X1 NAND3X1_117 ( .A(_69_), .B(_77_), .C(_74_), .Y(_78_) );
OAI21X1 OAI21X1_97 ( .A(i_add2[14]), .B(i_add1[14]), .C(_78_), .Y(_79_) );
INVX1 INVX1_234 ( .A(_79_), .Y(w_C_15_) );
INVX1 INVX1_235 ( .A(i_add2[15]), .Y(_80_) );
INVX1 INVX1_236 ( .A(i_add1[15]), .Y(_81_) );
NOR2X1 NOR2X1_132 ( .A(_80_), .B(_81_), .Y(_82_) );
INVX1 INVX1_237 ( .A(_82_), .Y(_83_) );
NOR2X1 NOR2X1_133 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_84_) );
INVX1 INVX1_238 ( .A(_84_), .Y(_85_) );
NOR2X1 NOR2X1_134 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_86_) );
INVX1 INVX1_239 ( .A(_86_), .Y(_87_) );
NAND3X1 NAND3X1_118 ( .A(_85_), .B(_87_), .C(_78_), .Y(_88_) );
AND2X2 AND2X2_103 ( .A(_88_), .B(_83_), .Y(_89_) );
INVX1 INVX1_240 ( .A(_89_), .Y(w_C_16_) );
AND2X2 AND2X2_104 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_90_) );
INVX1 INVX1_241 ( .A(_90_), .Y(_91_) );
NAND3X1 NAND3X1_119 ( .A(_83_), .B(_91_), .C(_88_), .Y(_92_) );
OAI21X1 OAI21X1_98 ( .A(i_add2[16]), .B(i_add1[16]), .C(_92_), .Y(_93_) );
INVX1 INVX1_242 ( .A(_93_), .Y(w_C_17_) );
INVX1 INVX1_243 ( .A(i_add2[17]), .Y(_94_) );
INVX1 INVX1_244 ( .A(i_add1[17]), .Y(_95_) );
NOR2X1 NOR2X1_135 ( .A(_94_), .B(_95_), .Y(_96_) );
INVX1 INVX1_245 ( .A(_96_), .Y(_97_) );
NOR2X1 NOR2X1_136 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_98_) );
INVX1 INVX1_246 ( .A(_98_), .Y(_99_) );
NOR2X1 NOR2X1_137 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_100_) );
INVX1 INVX1_247 ( .A(_100_), .Y(_101_) );
NAND3X1 NAND3X1_120 ( .A(_99_), .B(_101_), .C(_92_), .Y(_102_) );
AND2X2 AND2X2_105 ( .A(_102_), .B(_97_), .Y(_103_) );
INVX1 INVX1_248 ( .A(_103_), .Y(w_C_18_) );
AND2X2 AND2X2_106 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_104_) );
INVX1 INVX1_249 ( .A(_104_), .Y(_105_) );
NAND3X1 NAND3X1_121 ( .A(_97_), .B(_105_), .C(_102_), .Y(_106_) );
OAI21X1 OAI21X1_99 ( .A(i_add2[18]), .B(i_add1[18]), .C(_106_), .Y(_107_) );
INVX1 INVX1_250 ( .A(_107_), .Y(w_C_19_) );
INVX1 INVX1_251 ( .A(i_add2[19]), .Y(_108_) );
INVX1 INVX1_252 ( .A(i_add1[19]), .Y(_109_) );
NOR2X1 NOR2X1_138 ( .A(_108_), .B(_109_), .Y(_110_) );
INVX1 INVX1_253 ( .A(_110_), .Y(_111_) );
NOR2X1 NOR2X1_139 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_112_) );
INVX1 INVX1_254 ( .A(_112_), .Y(_113_) );
NOR2X1 NOR2X1_140 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_114_) );
INVX1 INVX1_255 ( .A(_114_), .Y(_115_) );
NAND3X1 NAND3X1_122 ( .A(_113_), .B(_115_), .C(_106_), .Y(_116_) );
AND2X2 AND2X2_107 ( .A(_116_), .B(_111_), .Y(_117_) );
INVX1 INVX1_256 ( .A(_117_), .Y(w_C_20_) );
AND2X2 AND2X2_108 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_118_) );
INVX1 INVX1_257 ( .A(_118_), .Y(_119_) );
NAND3X1 NAND3X1_123 ( .A(_111_), .B(_119_), .C(_116_), .Y(_120_) );
OAI21X1 OAI21X1_100 ( .A(i_add2[20]), .B(i_add1[20]), .C(_120_), .Y(_121_) );
INVX1 INVX1_258 ( .A(_121_), .Y(w_C_21_) );
INVX1 INVX1_259 ( .A(i_add2[21]), .Y(_122_) );
INVX1 INVX1_260 ( .A(i_add1[21]), .Y(_123_) );
NOR2X1 NOR2X1_141 ( .A(_122_), .B(_123_), .Y(_124_) );
INVX1 INVX1_261 ( .A(_124_), .Y(_125_) );
NOR2X1 NOR2X1_142 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_126_) );
INVX1 INVX1_262 ( .A(_126_), .Y(_127_) );
NOR2X1 NOR2X1_143 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_128_) );
INVX1 INVX1_263 ( .A(_128_), .Y(_129_) );
NAND3X1 NAND3X1_124 ( .A(_127_), .B(_129_), .C(_120_), .Y(_130_) );
AND2X2 AND2X2_109 ( .A(_130_), .B(_125_), .Y(_131_) );
INVX1 INVX1_264 ( .A(_131_), .Y(w_C_22_) );
AND2X2 AND2X2_110 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_132_) );
INVX1 INVX1_265 ( .A(_132_), .Y(_133_) );
NAND3X1 NAND3X1_125 ( .A(_125_), .B(_133_), .C(_130_), .Y(_134_) );
OAI21X1 OAI21X1_101 ( .A(i_add2[22]), .B(i_add1[22]), .C(_134_), .Y(_135_) );
INVX1 INVX1_266 ( .A(_135_), .Y(w_C_23_) );
INVX1 INVX1_267 ( .A(i_add2[23]), .Y(_136_) );
INVX1 INVX1_268 ( .A(i_add1[23]), .Y(_137_) );
NOR2X1 NOR2X1_144 ( .A(_136_), .B(_137_), .Y(_138_) );
INVX1 INVX1_269 ( .A(_138_), .Y(_139_) );
NOR2X1 NOR2X1_145 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_140_) );
INVX1 INVX1_270 ( .A(_140_), .Y(_141_) );
NOR2X1 NOR2X1_146 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_142_) );
INVX1 INVX1_271 ( .A(_142_), .Y(_143_) );
NAND3X1 NAND3X1_126 ( .A(_141_), .B(_143_), .C(_134_), .Y(_144_) );
AND2X2 AND2X2_111 ( .A(_144_), .B(_139_), .Y(_145_) );
INVX1 INVX1_272 ( .A(_145_), .Y(w_C_24_) );
AND2X2 AND2X2_112 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_146_) );
INVX1 INVX1_273 ( .A(_146_), .Y(_147_) );
BUFX2 BUFX2_66 ( .A(w_C_64_), .Y(_399__64_) );
BUFX2 BUFX2_67 ( .A(gnd), .Y(w_C_0_) );
endmodule
