module cla_34bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add1[19], i_add1[20], i_add1[21], i_add1[22], i_add1[23], i_add1[24], i_add1[25], i_add1[26], i_add1[27], i_add1[28], i_add1[29], i_add1[30], i_add1[31], i_add1[32], i_add1[33], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], i_add2[19], i_add2[20], i_add2[21], i_add2[22], i_add2[23], i_add2[24], i_add2[25], i_add2[26], i_add2[27], i_add2[28], i_add2[29], i_add2[30], i_add2[31], i_add2[32], i_add2[33], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21], o_result[22], o_result[23], o_result[24], o_result[25], o_result[26], o_result[27], o_result[28], o_result[29], o_result[30], o_result[31], o_result[32], o_result[33], o_result[34]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add1[19];
input i_add1[20];
input i_add1[21];
input i_add1[22];
input i_add1[23];
input i_add1[24];
input i_add1[25];
input i_add1[26];
input i_add1[27];
input i_add1[28];
input i_add1[29];
input i_add1[30];
input i_add1[31];
input i_add1[32];
input i_add1[33];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
input i_add2[19];
input i_add2[20];
input i_add2[21];
input i_add2[22];
input i_add2[23];
input i_add2[24];
input i_add2[25];
input i_add2[26];
input i_add2[27];
input i_add2[28];
input i_add2[29];
input i_add2[30];
input i_add2[31];
input i_add2[32];
input i_add2[33];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];
output o_result[22];
output o_result[23];
output o_result[24];
output o_result[25];
output o_result[26];
output o_result[27];
output o_result[28];
output o_result[29];
output o_result[30];
output o_result[31];
output o_result[32];
output o_result[33];
output o_result[34];

NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_1 ( .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_2 ( .A(_1_), .B(_2_), .Y(w_C_2_) );
INVX1 INVX1_2 ( .A(i_add2[2]), .Y(_3_) );
INVX1 INVX1_3 ( .A(i_add1[2]), .Y(_4_) );
NAND2X1 NAND2X1_2 ( .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
OAI21X1 OAI21X1_1 ( .A(_1_), .B(_2_), .C(_6_), .Y(_7_) );
AND2X2 AND2X2_1 ( .A(_7_), .B(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
OR2X2 OR2X2_1 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_1 ( .A(_5_), .B(_9_), .C(_7_), .Y(_10_) );
AND2X2 AND2X2_2 ( .A(_10_), .B(_8_), .Y(_11_) );
INVX1 INVX1_4 ( .A(_11_), .Y(w_C_4_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_12_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
OAI21X1 OAI21X1_2 ( .A(_13_), .B(_11_), .C(_12_), .Y(w_C_5_) );
AND2X2 AND2X2_3 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_14_) );
INVX1 INVX1_5 ( .A(_14_), .Y(_15_) );
INVX1 INVX1_6 ( .A(_13_), .Y(_16_) );
NAND3X1 NAND3X1_2 ( .A(_8_), .B(_12_), .C(_10_), .Y(_17_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_18_) );
INVX1 INVX1_7 ( .A(_18_), .Y(_19_) );
NAND3X1 NAND3X1_3 ( .A(_16_), .B(_19_), .C(_17_), .Y(_20_) );
AND2X2 AND2X2_4 ( .A(_20_), .B(_15_), .Y(_21_) );
INVX1 INVX1_8 ( .A(_21_), .Y(w_C_6_) );
AND2X2 AND2X2_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_9 ( .A(_22_), .Y(_23_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_24_) );
OAI21X1 OAI21X1_3 ( .A(_24_), .B(_21_), .C(_23_), .Y(w_C_7_) );
INVX1 INVX1_10 ( .A(i_add2[7]), .Y(_25_) );
INVX1 INVX1_11 ( .A(i_add1[7]), .Y(_26_) );
INVX1 INVX1_12 ( .A(_24_), .Y(_27_) );
NAND3X1 NAND3X1_4 ( .A(_15_), .B(_23_), .C(_20_), .Y(_28_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_29_) );
INVX1 INVX1_13 ( .A(_29_), .Y(_30_) );
NAND3X1 NAND3X1_5 ( .A(_27_), .B(_30_), .C(_28_), .Y(_31_) );
OAI21X1 OAI21X1_4 ( .A(_25_), .B(_26_), .C(_31_), .Y(w_C_8_) );
NOR2X1 NOR2X1_7 ( .A(_25_), .B(_26_), .Y(_32_) );
INVX1 INVX1_14 ( .A(_32_), .Y(_33_) );
AND2X2 AND2X2_6 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_34_) );
INVX1 INVX1_15 ( .A(_34_), .Y(_35_) );
NAND3X1 NAND3X1_6 ( .A(_33_), .B(_35_), .C(_31_), .Y(_36_) );
OAI21X1 OAI21X1_5 ( .A(i_add2[8]), .B(i_add1[8]), .C(_36_), .Y(_37_) );
INVX1 INVX1_16 ( .A(_37_), .Y(w_C_9_) );
INVX1 INVX1_17 ( .A(i_add2[9]), .Y(_38_) );
INVX1 INVX1_18 ( .A(i_add1[9]), .Y(_39_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_40_) );
INVX1 INVX1_19 ( .A(_40_), .Y(_41_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_42_) );
INVX1 INVX1_20 ( .A(_42_), .Y(_43_) );
NAND3X1 NAND3X1_7 ( .A(_41_), .B(_43_), .C(_36_), .Y(_44_) );
OAI21X1 OAI21X1_6 ( .A(_38_), .B(_39_), .C(_44_), .Y(w_C_10_) );
NOR2X1 NOR2X1_10 ( .A(_38_), .B(_39_), .Y(_45_) );
INVX1 INVX1_21 ( .A(_45_), .Y(_46_) );
AND2X2 AND2X2_7 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_47_) );
INVX1 INVX1_22 ( .A(_47_), .Y(_48_) );
NAND3X1 NAND3X1_8 ( .A(_46_), .B(_48_), .C(_44_), .Y(_49_) );
OAI21X1 OAI21X1_7 ( .A(i_add2[10]), .B(i_add1[10]), .C(_49_), .Y(_50_) );
INVX1 INVX1_23 ( .A(_50_), .Y(w_C_11_) );
INVX1 INVX1_24 ( .A(i_add2[11]), .Y(_51_) );
INVX1 INVX1_25 ( .A(i_add1[11]), .Y(_52_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_53_) );
INVX1 INVX1_26 ( .A(_53_), .Y(_54_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_55_) );
INVX1 INVX1_27 ( .A(_55_), .Y(_56_) );
NAND3X1 NAND3X1_9 ( .A(_54_), .B(_56_), .C(_49_), .Y(_57_) );
OAI21X1 OAI21X1_8 ( .A(_51_), .B(_52_), .C(_57_), .Y(w_C_12_) );
NOR2X1 NOR2X1_13 ( .A(_51_), .B(_52_), .Y(_58_) );
INVX1 INVX1_28 ( .A(_58_), .Y(_59_) );
AND2X2 AND2X2_8 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_60_) );
INVX1 INVX1_29 ( .A(_60_), .Y(_61_) );
NAND3X1 NAND3X1_10 ( .A(_59_), .B(_61_), .C(_57_), .Y(_62_) );
OAI21X1 OAI21X1_9 ( .A(i_add2[12]), .B(i_add1[12]), .C(_62_), .Y(_63_) );
INVX1 INVX1_30 ( .A(_63_), .Y(w_C_13_) );
INVX1 INVX1_31 ( .A(i_add2[13]), .Y(_64_) );
INVX1 INVX1_32 ( .A(i_add1[13]), .Y(_65_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_66_) );
INVX1 INVX1_33 ( .A(_66_), .Y(_67_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_68_) );
INVX1 INVX1_34 ( .A(_68_), .Y(_69_) );
NAND3X1 NAND3X1_11 ( .A(_67_), .B(_69_), .C(_62_), .Y(_70_) );
OAI21X1 OAI21X1_10 ( .A(_64_), .B(_65_), .C(_70_), .Y(w_C_14_) );
NOR2X1 NOR2X1_16 ( .A(_64_), .B(_65_), .Y(_71_) );
INVX1 INVX1_35 ( .A(_71_), .Y(_72_) );
AND2X2 AND2X2_9 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_73_) );
INVX1 INVX1_36 ( .A(_73_), .Y(_74_) );
NAND3X1 NAND3X1_12 ( .A(_72_), .B(_74_), .C(_70_), .Y(_75_) );
OAI21X1 OAI21X1_11 ( .A(i_add2[14]), .B(i_add1[14]), .C(_75_), .Y(_76_) );
INVX1 INVX1_37 ( .A(_76_), .Y(w_C_15_) );
INVX1 INVX1_38 ( .A(i_add2[15]), .Y(_77_) );
INVX1 INVX1_39 ( .A(i_add1[15]), .Y(_78_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_79_) );
INVX1 INVX1_40 ( .A(_79_), .Y(_80_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_81_) );
INVX1 INVX1_41 ( .A(_81_), .Y(_82_) );
NAND3X1 NAND3X1_13 ( .A(_80_), .B(_82_), .C(_75_), .Y(_83_) );
OAI21X1 OAI21X1_12 ( .A(_77_), .B(_78_), .C(_83_), .Y(w_C_16_) );
NOR2X1 NOR2X1_19 ( .A(_77_), .B(_78_), .Y(_84_) );
INVX1 INVX1_42 ( .A(_84_), .Y(_85_) );
AND2X2 AND2X2_10 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_86_) );
INVX1 INVX1_43 ( .A(_86_), .Y(_87_) );
NAND3X1 NAND3X1_14 ( .A(_85_), .B(_87_), .C(_83_), .Y(_88_) );
OAI21X1 OAI21X1_13 ( .A(i_add2[16]), .B(i_add1[16]), .C(_88_), .Y(_89_) );
INVX1 INVX1_44 ( .A(_89_), .Y(w_C_17_) );
INVX1 INVX1_45 ( .A(i_add2[17]), .Y(_90_) );
INVX1 INVX1_46 ( .A(i_add1[17]), .Y(_91_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_92_) );
INVX1 INVX1_47 ( .A(_92_), .Y(_93_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_94_) );
INVX1 INVX1_48 ( .A(_94_), .Y(_95_) );
NAND3X1 NAND3X1_15 ( .A(_93_), .B(_95_), .C(_88_), .Y(_96_) );
OAI21X1 OAI21X1_14 ( .A(_90_), .B(_91_), .C(_96_), .Y(w_C_18_) );
NOR2X1 NOR2X1_22 ( .A(_90_), .B(_91_), .Y(_97_) );
INVX1 INVX1_49 ( .A(_97_), .Y(_98_) );
AND2X2 AND2X2_11 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_99_) );
INVX1 INVX1_50 ( .A(_99_), .Y(_100_) );
NAND3X1 NAND3X1_16 ( .A(_98_), .B(_100_), .C(_96_), .Y(_101_) );
OAI21X1 OAI21X1_15 ( .A(i_add2[18]), .B(i_add1[18]), .C(_101_), .Y(_102_) );
INVX1 INVX1_51 ( .A(_102_), .Y(w_C_19_) );
INVX1 INVX1_52 ( .A(i_add2[19]), .Y(_103_) );
INVX1 INVX1_53 ( .A(i_add1[19]), .Y(_104_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_105_) );
INVX1 INVX1_54 ( .A(_105_), .Y(_106_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_107_) );
INVX1 INVX1_55 ( .A(_107_), .Y(_108_) );
NAND3X1 NAND3X1_17 ( .A(_106_), .B(_108_), .C(_101_), .Y(_109_) );
OAI21X1 OAI21X1_16 ( .A(_103_), .B(_104_), .C(_109_), .Y(w_C_20_) );
NOR2X1 NOR2X1_25 ( .A(_103_), .B(_104_), .Y(_110_) );
INVX1 INVX1_56 ( .A(_110_), .Y(_111_) );
AND2X2 AND2X2_12 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_112_) );
INVX1 INVX1_57 ( .A(_112_), .Y(_113_) );
NAND3X1 NAND3X1_18 ( .A(_111_), .B(_113_), .C(_109_), .Y(_114_) );
OAI21X1 OAI21X1_17 ( .A(i_add2[20]), .B(i_add1[20]), .C(_114_), .Y(_115_) );
INVX1 INVX1_58 ( .A(_115_), .Y(w_C_21_) );
INVX1 INVX1_59 ( .A(i_add2[21]), .Y(_116_) );
INVX1 INVX1_60 ( .A(i_add1[21]), .Y(_117_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_118_) );
INVX1 INVX1_61 ( .A(_118_), .Y(_119_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_120_) );
INVX1 INVX1_62 ( .A(_120_), .Y(_121_) );
NAND3X1 NAND3X1_19 ( .A(_119_), .B(_121_), .C(_114_), .Y(_122_) );
OAI21X1 OAI21X1_18 ( .A(_116_), .B(_117_), .C(_122_), .Y(w_C_22_) );
NOR2X1 NOR2X1_28 ( .A(_116_), .B(_117_), .Y(_123_) );
INVX1 INVX1_63 ( .A(_123_), .Y(_124_) );
AND2X2 AND2X2_13 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_125_) );
INVX1 INVX1_64 ( .A(_125_), .Y(_126_) );
NAND3X1 NAND3X1_20 ( .A(_124_), .B(_126_), .C(_122_), .Y(_127_) );
OAI21X1 OAI21X1_19 ( .A(i_add2[22]), .B(i_add1[22]), .C(_127_), .Y(_128_) );
INVX1 INVX1_65 ( .A(_128_), .Y(w_C_23_) );
INVX1 INVX1_66 ( .A(i_add2[23]), .Y(_129_) );
INVX1 INVX1_67 ( .A(i_add1[23]), .Y(_130_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_131_) );
INVX1 INVX1_68 ( .A(_131_), .Y(_132_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_133_) );
INVX1 INVX1_69 ( .A(_133_), .Y(_134_) );
NAND3X1 NAND3X1_21 ( .A(_132_), .B(_134_), .C(_127_), .Y(_135_) );
OAI21X1 OAI21X1_20 ( .A(_129_), .B(_130_), .C(_135_), .Y(w_C_24_) );
NOR2X1 NOR2X1_31 ( .A(_129_), .B(_130_), .Y(_136_) );
INVX1 INVX1_70 ( .A(_136_), .Y(_137_) );
AND2X2 AND2X2_14 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_138_) );
INVX1 INVX1_71 ( .A(_138_), .Y(_139_) );
NAND3X1 NAND3X1_22 ( .A(_137_), .B(_139_), .C(_135_), .Y(_140_) );
OAI21X1 OAI21X1_21 ( .A(i_add2[24]), .B(i_add1[24]), .C(_140_), .Y(_141_) );
INVX1 INVX1_72 ( .A(_141_), .Y(w_C_25_) );
INVX1 INVX1_73 ( .A(i_add2[25]), .Y(_142_) );
INVX1 INVX1_74 ( .A(i_add1[25]), .Y(_143_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_144_) );
INVX1 INVX1_75 ( .A(_144_), .Y(_145_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_146_) );
INVX1 INVX1_76 ( .A(_146_), .Y(_147_) );
NAND3X1 NAND3X1_23 ( .A(_145_), .B(_147_), .C(_140_), .Y(_148_) );
OAI21X1 OAI21X1_22 ( .A(_142_), .B(_143_), .C(_148_), .Y(w_C_26_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_149_) );
INVX1 INVX1_77 ( .A(_149_), .Y(_150_) );
NOR2X1 NOR2X1_35 ( .A(_142_), .B(_143_), .Y(_151_) );
INVX1 INVX1_78 ( .A(_151_), .Y(_152_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_153_) );
NAND3X1 NAND3X1_24 ( .A(_152_), .B(_153_), .C(_148_), .Y(_154_) );
AND2X2 AND2X2_15 ( .A(_154_), .B(_150_), .Y(w_C_27_) );
INVX1 INVX1_79 ( .A(i_add2[27]), .Y(_155_) );
INVX1 INVX1_80 ( .A(i_add1[27]), .Y(_156_) );
NAND2X1 NAND2X1_7 ( .A(_155_), .B(_156_), .Y(_157_) );
NAND3X1 NAND3X1_25 ( .A(_150_), .B(_157_), .C(_154_), .Y(_158_) );
OAI21X1 OAI21X1_23 ( .A(_155_), .B(_156_), .C(_158_), .Y(w_C_28_) );
INVX1 INVX1_81 ( .A(i_add2[28]), .Y(_159_) );
INVX1 INVX1_82 ( .A(i_add1[28]), .Y(_160_) );
NAND2X1 NAND2X1_8 ( .A(_159_), .B(_160_), .Y(_161_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_162_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_163_) );
NAND3X1 NAND3X1_26 ( .A(_162_), .B(_163_), .C(_158_), .Y(_164_) );
AND2X2 AND2X2_16 ( .A(_164_), .B(_161_), .Y(w_C_29_) );
INVX1 INVX1_83 ( .A(i_add2[29]), .Y(_165_) );
INVX1 INVX1_84 ( .A(i_add1[29]), .Y(_166_) );
NAND2X1 NAND2X1_11 ( .A(_165_), .B(_166_), .Y(_167_) );
NAND3X1 NAND3X1_27 ( .A(_161_), .B(_167_), .C(_164_), .Y(_168_) );
OAI21X1 OAI21X1_24 ( .A(_165_), .B(_166_), .C(_168_), .Y(w_C_30_) );
NOR2X1 NOR2X1_36 ( .A(_165_), .B(_166_), .Y(_169_) );
INVX1 INVX1_85 ( .A(_169_), .Y(_170_) );
AND2X2 AND2X2_17 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_171_) );
INVX1 INVX1_86 ( .A(_171_), .Y(_172_) );
NAND3X1 NAND3X1_28 ( .A(_170_), .B(_172_), .C(_168_), .Y(_173_) );
OAI21X1 OAI21X1_25 ( .A(i_add2[30]), .B(i_add1[30]), .C(_173_), .Y(_174_) );
INVX1 INVX1_87 ( .A(_174_), .Y(w_C_31_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_175_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_176_) );
OAI21X1 OAI21X1_26 ( .A(_176_), .B(_174_), .C(_175_), .Y(w_C_32_) );
OR2X2 OR2X2_2 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_177_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_178_) );
INVX1 INVX1_88 ( .A(_178_), .Y(_179_) );
INVX1 INVX1_89 ( .A(_176_), .Y(_180_) );
NAND3X1 NAND3X1_29 ( .A(_179_), .B(_180_), .C(_173_), .Y(_181_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_182_) );
NAND3X1 NAND3X1_30 ( .A(_175_), .B(_182_), .C(_181_), .Y(_183_) );
AND2X2 AND2X2_18 ( .A(_183_), .B(_177_), .Y(w_C_33_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_184_) );
OR2X2 OR2X2_3 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_185_) );
NAND3X1 NAND3X1_31 ( .A(_177_), .B(_185_), .C(_183_), .Y(_186_) );
NAND2X1 NAND2X1_15 ( .A(_184_), .B(_186_), .Y(w_C_34_) );
BUFX2 BUFX2_1 ( .A(_187__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_187__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_187__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_187__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_187__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_187__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_187__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_187__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_187__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_187__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_187__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_187__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_187__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_187__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_187__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_187__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_187__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_187__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_187__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_187__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_187__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_187__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_187__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_187__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_187__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_187__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_187__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_187__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_187__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_187__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_187__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_187__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_187__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_187__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(w_C_34_), .Y(o_result[34]) );
INVX1 INVX1_90 ( .A(w_C_4_), .Y(_191_) );
OR2X2 OR2X2_4 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_192_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_193_) );
NAND3X1 NAND3X1_32 ( .A(_191_), .B(_193_), .C(_192_), .Y(_194_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_188_) );
AND2X2 AND2X2_19 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_189_) );
OAI21X1 OAI21X1_27 ( .A(_188_), .B(_189_), .C(w_C_4_), .Y(_190_) );
NAND2X1 NAND2X1_17 ( .A(_190_), .B(_194_), .Y(_187__4_) );
INVX1 INVX1_91 ( .A(w_C_5_), .Y(_198_) );
OR2X2 OR2X2_5 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_199_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_200_) );
NAND3X1 NAND3X1_33 ( .A(_198_), .B(_200_), .C(_199_), .Y(_201_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_195_) );
AND2X2 AND2X2_20 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_196_) );
OAI21X1 OAI21X1_28 ( .A(_195_), .B(_196_), .C(w_C_5_), .Y(_197_) );
NAND2X1 NAND2X1_19 ( .A(_197_), .B(_201_), .Y(_187__5_) );
INVX1 INVX1_92 ( .A(w_C_6_), .Y(_205_) );
OR2X2 OR2X2_6 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_206_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_207_) );
NAND3X1 NAND3X1_34 ( .A(_205_), .B(_207_), .C(_206_), .Y(_208_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_202_) );
AND2X2 AND2X2_21 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_203_) );
OAI21X1 OAI21X1_29 ( .A(_202_), .B(_203_), .C(w_C_6_), .Y(_204_) );
NAND2X1 NAND2X1_21 ( .A(_204_), .B(_208_), .Y(_187__6_) );
INVX1 INVX1_93 ( .A(w_C_7_), .Y(_212_) );
OR2X2 OR2X2_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_213_) );
NAND2X1 NAND2X1_22 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_214_) );
NAND3X1 NAND3X1_35 ( .A(_212_), .B(_214_), .C(_213_), .Y(_215_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_209_) );
AND2X2 AND2X2_22 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_210_) );
OAI21X1 OAI21X1_30 ( .A(_209_), .B(_210_), .C(w_C_7_), .Y(_211_) );
NAND2X1 NAND2X1_23 ( .A(_211_), .B(_215_), .Y(_187__7_) );
INVX1 INVX1_94 ( .A(w_C_8_), .Y(_219_) );
OR2X2 OR2X2_8 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_220_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_221_) );
NAND3X1 NAND3X1_36 ( .A(_219_), .B(_221_), .C(_220_), .Y(_222_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_216_) );
AND2X2 AND2X2_23 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_217_) );
OAI21X1 OAI21X1_31 ( .A(_216_), .B(_217_), .C(w_C_8_), .Y(_218_) );
NAND2X1 NAND2X1_25 ( .A(_218_), .B(_222_), .Y(_187__8_) );
INVX1 INVX1_95 ( .A(w_C_9_), .Y(_226_) );
OR2X2 OR2X2_9 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_227_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_228_) );
NAND3X1 NAND3X1_37 ( .A(_226_), .B(_228_), .C(_227_), .Y(_229_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_223_) );
AND2X2 AND2X2_24 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_224_) );
OAI21X1 OAI21X1_32 ( .A(_223_), .B(_224_), .C(w_C_9_), .Y(_225_) );
NAND2X1 NAND2X1_27 ( .A(_225_), .B(_229_), .Y(_187__9_) );
INVX1 INVX1_96 ( .A(w_C_10_), .Y(_233_) );
OR2X2 OR2X2_10 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_234_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_235_) );
NAND3X1 NAND3X1_38 ( .A(_233_), .B(_235_), .C(_234_), .Y(_236_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_230_) );
AND2X2 AND2X2_25 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_231_) );
OAI21X1 OAI21X1_33 ( .A(_230_), .B(_231_), .C(w_C_10_), .Y(_232_) );
NAND2X1 NAND2X1_29 ( .A(_232_), .B(_236_), .Y(_187__10_) );
INVX1 INVX1_97 ( .A(w_C_11_), .Y(_240_) );
OR2X2 OR2X2_11 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_241_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_242_) );
NAND3X1 NAND3X1_39 ( .A(_240_), .B(_242_), .C(_241_), .Y(_243_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_237_) );
AND2X2 AND2X2_26 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_238_) );
OAI21X1 OAI21X1_34 ( .A(_237_), .B(_238_), .C(w_C_11_), .Y(_239_) );
NAND2X1 NAND2X1_31 ( .A(_239_), .B(_243_), .Y(_187__11_) );
INVX1 INVX1_98 ( .A(w_C_12_), .Y(_247_) );
OR2X2 OR2X2_12 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_248_) );
NAND2X1 NAND2X1_32 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_249_) );
NAND3X1 NAND3X1_40 ( .A(_247_), .B(_249_), .C(_248_), .Y(_250_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_244_) );
AND2X2 AND2X2_27 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_245_) );
OAI21X1 OAI21X1_35 ( .A(_244_), .B(_245_), .C(w_C_12_), .Y(_246_) );
NAND2X1 NAND2X1_33 ( .A(_246_), .B(_250_), .Y(_187__12_) );
INVX1 INVX1_99 ( .A(w_C_13_), .Y(_254_) );
OR2X2 OR2X2_13 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_255_) );
NAND2X1 NAND2X1_34 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_256_) );
NAND3X1 NAND3X1_41 ( .A(_254_), .B(_256_), .C(_255_), .Y(_257_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_251_) );
AND2X2 AND2X2_28 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_252_) );
OAI21X1 OAI21X1_36 ( .A(_251_), .B(_252_), .C(w_C_13_), .Y(_253_) );
NAND2X1 NAND2X1_35 ( .A(_253_), .B(_257_), .Y(_187__13_) );
INVX1 INVX1_100 ( .A(w_C_14_), .Y(_261_) );
OR2X2 OR2X2_14 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_262_) );
NAND2X1 NAND2X1_36 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_263_) );
NAND3X1 NAND3X1_42 ( .A(_261_), .B(_263_), .C(_262_), .Y(_264_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_258_) );
AND2X2 AND2X2_29 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_259_) );
OAI21X1 OAI21X1_37 ( .A(_258_), .B(_259_), .C(w_C_14_), .Y(_260_) );
NAND2X1 NAND2X1_37 ( .A(_260_), .B(_264_), .Y(_187__14_) );
INVX1 INVX1_101 ( .A(w_C_15_), .Y(_268_) );
OR2X2 OR2X2_15 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_269_) );
NAND2X1 NAND2X1_38 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_270_) );
NAND3X1 NAND3X1_43 ( .A(_268_), .B(_270_), .C(_269_), .Y(_271_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_265_) );
AND2X2 AND2X2_30 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_266_) );
OAI21X1 OAI21X1_38 ( .A(_265_), .B(_266_), .C(w_C_15_), .Y(_267_) );
NAND2X1 NAND2X1_39 ( .A(_267_), .B(_271_), .Y(_187__15_) );
INVX1 INVX1_102 ( .A(w_C_16_), .Y(_275_) );
OR2X2 OR2X2_16 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_276_) );
NAND2X1 NAND2X1_40 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_277_) );
NAND3X1 NAND3X1_44 ( .A(_275_), .B(_277_), .C(_276_), .Y(_278_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_272_) );
AND2X2 AND2X2_31 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_273_) );
OAI21X1 OAI21X1_39 ( .A(_272_), .B(_273_), .C(w_C_16_), .Y(_274_) );
NAND2X1 NAND2X1_41 ( .A(_274_), .B(_278_), .Y(_187__16_) );
INVX1 INVX1_103 ( .A(w_C_17_), .Y(_282_) );
OR2X2 OR2X2_17 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_283_) );
NAND2X1 NAND2X1_42 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_284_) );
NAND3X1 NAND3X1_45 ( .A(_282_), .B(_284_), .C(_283_), .Y(_285_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_279_) );
AND2X2 AND2X2_32 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_280_) );
OAI21X1 OAI21X1_40 ( .A(_279_), .B(_280_), .C(w_C_17_), .Y(_281_) );
NAND2X1 NAND2X1_43 ( .A(_281_), .B(_285_), .Y(_187__17_) );
INVX1 INVX1_104 ( .A(w_C_18_), .Y(_289_) );
OR2X2 OR2X2_18 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_290_) );
NAND2X1 NAND2X1_44 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_291_) );
NAND3X1 NAND3X1_46 ( .A(_289_), .B(_291_), .C(_290_), .Y(_292_) );
NOR2X1 NOR2X1_53 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_286_) );
AND2X2 AND2X2_33 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_287_) );
OAI21X1 OAI21X1_41 ( .A(_286_), .B(_287_), .C(w_C_18_), .Y(_288_) );
NAND2X1 NAND2X1_45 ( .A(_288_), .B(_292_), .Y(_187__18_) );
INVX1 INVX1_105 ( .A(w_C_19_), .Y(_296_) );
OR2X2 OR2X2_19 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_297_) );
NAND2X1 NAND2X1_46 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_298_) );
NAND3X1 NAND3X1_47 ( .A(_296_), .B(_298_), .C(_297_), .Y(_299_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_293_) );
AND2X2 AND2X2_34 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_294_) );
OAI21X1 OAI21X1_42 ( .A(_293_), .B(_294_), .C(w_C_19_), .Y(_295_) );
NAND2X1 NAND2X1_47 ( .A(_295_), .B(_299_), .Y(_187__19_) );
INVX1 INVX1_106 ( .A(w_C_20_), .Y(_303_) );
OR2X2 OR2X2_20 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_304_) );
NAND2X1 NAND2X1_48 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_305_) );
NAND3X1 NAND3X1_48 ( .A(_303_), .B(_305_), .C(_304_), .Y(_306_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_300_) );
AND2X2 AND2X2_35 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_301_) );
OAI21X1 OAI21X1_43 ( .A(_300_), .B(_301_), .C(w_C_20_), .Y(_302_) );
NAND2X1 NAND2X1_49 ( .A(_302_), .B(_306_), .Y(_187__20_) );
INVX1 INVX1_107 ( .A(w_C_21_), .Y(_310_) );
OR2X2 OR2X2_21 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_311_) );
NAND2X1 NAND2X1_50 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_312_) );
NAND3X1 NAND3X1_49 ( .A(_310_), .B(_312_), .C(_311_), .Y(_313_) );
NOR2X1 NOR2X1_56 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_307_) );
AND2X2 AND2X2_36 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_308_) );
OAI21X1 OAI21X1_44 ( .A(_307_), .B(_308_), .C(w_C_21_), .Y(_309_) );
NAND2X1 NAND2X1_51 ( .A(_309_), .B(_313_), .Y(_187__21_) );
INVX1 INVX1_108 ( .A(w_C_22_), .Y(_317_) );
OR2X2 OR2X2_22 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_318_) );
NAND2X1 NAND2X1_52 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_319_) );
NAND3X1 NAND3X1_50 ( .A(_317_), .B(_319_), .C(_318_), .Y(_320_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_314_) );
AND2X2 AND2X2_37 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_315_) );
OAI21X1 OAI21X1_45 ( .A(_314_), .B(_315_), .C(w_C_22_), .Y(_316_) );
NAND2X1 NAND2X1_53 ( .A(_316_), .B(_320_), .Y(_187__22_) );
INVX1 INVX1_109 ( .A(w_C_23_), .Y(_324_) );
OR2X2 OR2X2_23 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_325_) );
NAND2X1 NAND2X1_54 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_326_) );
NAND3X1 NAND3X1_51 ( .A(_324_), .B(_326_), .C(_325_), .Y(_327_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_321_) );
AND2X2 AND2X2_38 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_322_) );
OAI21X1 OAI21X1_46 ( .A(_321_), .B(_322_), .C(w_C_23_), .Y(_323_) );
NAND2X1 NAND2X1_55 ( .A(_323_), .B(_327_), .Y(_187__23_) );
INVX1 INVX1_110 ( .A(w_C_24_), .Y(_331_) );
OR2X2 OR2X2_24 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_332_) );
NAND2X1 NAND2X1_56 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_333_) );
NAND3X1 NAND3X1_52 ( .A(_331_), .B(_333_), .C(_332_), .Y(_334_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_328_) );
AND2X2 AND2X2_39 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_329_) );
OAI21X1 OAI21X1_47 ( .A(_328_), .B(_329_), .C(w_C_24_), .Y(_330_) );
NAND2X1 NAND2X1_57 ( .A(_330_), .B(_334_), .Y(_187__24_) );
INVX1 INVX1_111 ( .A(w_C_25_), .Y(_338_) );
OR2X2 OR2X2_25 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_339_) );
NAND2X1 NAND2X1_58 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_340_) );
NAND3X1 NAND3X1_53 ( .A(_338_), .B(_340_), .C(_339_), .Y(_341_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_335_) );
AND2X2 AND2X2_40 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_336_) );
OAI21X1 OAI21X1_48 ( .A(_335_), .B(_336_), .C(w_C_25_), .Y(_337_) );
NAND2X1 NAND2X1_59 ( .A(_337_), .B(_341_), .Y(_187__25_) );
INVX1 INVX1_112 ( .A(w_C_26_), .Y(_345_) );
OR2X2 OR2X2_26 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_346_) );
NAND2X1 NAND2X1_60 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_347_) );
NAND3X1 NAND3X1_54 ( .A(_345_), .B(_347_), .C(_346_), .Y(_348_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_342_) );
AND2X2 AND2X2_41 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_343_) );
OAI21X1 OAI21X1_49 ( .A(_342_), .B(_343_), .C(w_C_26_), .Y(_344_) );
NAND2X1 NAND2X1_61 ( .A(_344_), .B(_348_), .Y(_187__26_) );
INVX1 INVX1_113 ( .A(w_C_27_), .Y(_352_) );
OR2X2 OR2X2_27 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_353_) );
NAND2X1 NAND2X1_62 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_354_) );
NAND3X1 NAND3X1_55 ( .A(_352_), .B(_354_), .C(_353_), .Y(_355_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_349_) );
AND2X2 AND2X2_42 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_350_) );
OAI21X1 OAI21X1_50 ( .A(_349_), .B(_350_), .C(w_C_27_), .Y(_351_) );
NAND2X1 NAND2X1_63 ( .A(_351_), .B(_355_), .Y(_187__27_) );
INVX1 INVX1_114 ( .A(w_C_28_), .Y(_359_) );
OR2X2 OR2X2_28 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_360_) );
NAND2X1 NAND2X1_64 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_361_) );
NAND3X1 NAND3X1_56 ( .A(_359_), .B(_361_), .C(_360_), .Y(_362_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_356_) );
AND2X2 AND2X2_43 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_357_) );
OAI21X1 OAI21X1_51 ( .A(_356_), .B(_357_), .C(w_C_28_), .Y(_358_) );
NAND2X1 NAND2X1_65 ( .A(_358_), .B(_362_), .Y(_187__28_) );
INVX1 INVX1_115 ( .A(w_C_29_), .Y(_366_) );
OR2X2 OR2X2_29 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_367_) );
NAND2X1 NAND2X1_66 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_368_) );
NAND3X1 NAND3X1_57 ( .A(_366_), .B(_368_), .C(_367_), .Y(_369_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_363_) );
AND2X2 AND2X2_44 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_364_) );
OAI21X1 OAI21X1_52 ( .A(_363_), .B(_364_), .C(w_C_29_), .Y(_365_) );
NAND2X1 NAND2X1_67 ( .A(_365_), .B(_369_), .Y(_187__29_) );
INVX1 INVX1_116 ( .A(w_C_30_), .Y(_373_) );
OR2X2 OR2X2_30 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_374_) );
NAND2X1 NAND2X1_68 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_375_) );
NAND3X1 NAND3X1_58 ( .A(_373_), .B(_375_), .C(_374_), .Y(_376_) );
NOR2X1 NOR2X1_65 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_370_) );
AND2X2 AND2X2_45 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_371_) );
OAI21X1 OAI21X1_53 ( .A(_370_), .B(_371_), .C(w_C_30_), .Y(_372_) );
NAND2X1 NAND2X1_69 ( .A(_372_), .B(_376_), .Y(_187__30_) );
INVX1 INVX1_117 ( .A(w_C_31_), .Y(_380_) );
OR2X2 OR2X2_31 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_381_) );
NAND2X1 NAND2X1_70 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_382_) );
NAND3X1 NAND3X1_59 ( .A(_380_), .B(_382_), .C(_381_), .Y(_383_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_377_) );
AND2X2 AND2X2_46 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_378_) );
OAI21X1 OAI21X1_54 ( .A(_377_), .B(_378_), .C(w_C_31_), .Y(_379_) );
NAND2X1 NAND2X1_71 ( .A(_379_), .B(_383_), .Y(_187__31_) );
INVX1 INVX1_118 ( .A(w_C_32_), .Y(_387_) );
OR2X2 OR2X2_32 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_388_) );
NAND2X1 NAND2X1_72 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_389_) );
NAND3X1 NAND3X1_60 ( .A(_387_), .B(_389_), .C(_388_), .Y(_390_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_384_) );
AND2X2 AND2X2_47 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_385_) );
OAI21X1 OAI21X1_55 ( .A(_384_), .B(_385_), .C(w_C_32_), .Y(_386_) );
NAND2X1 NAND2X1_73 ( .A(_386_), .B(_390_), .Y(_187__32_) );
INVX1 INVX1_119 ( .A(w_C_33_), .Y(_394_) );
OR2X2 OR2X2_33 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_395_) );
NAND2X1 NAND2X1_74 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_396_) );
NAND3X1 NAND3X1_61 ( .A(_394_), .B(_396_), .C(_395_), .Y(_397_) );
NOR2X1 NOR2X1_68 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_391_) );
AND2X2 AND2X2_48 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_392_) );
OAI21X1 OAI21X1_56 ( .A(_391_), .B(_392_), .C(w_C_33_), .Y(_393_) );
NAND2X1 NAND2X1_75 ( .A(_393_), .B(_397_), .Y(_187__33_) );
INVX1 INVX1_120 ( .A(1'b0), .Y(_401_) );
OR2X2 OR2X2_34 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_402_) );
NAND2X1 NAND2X1_76 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_403_) );
NAND3X1 NAND3X1_62 ( .A(_401_), .B(_403_), .C(_402_), .Y(_404_) );
NOR2X1 NOR2X1_69 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_398_) );
AND2X2 AND2X2_49 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_399_) );
OAI21X1 OAI21X1_57 ( .A(_398_), .B(_399_), .C(1'b0), .Y(_400_) );
NAND2X1 NAND2X1_77 ( .A(_400_), .B(_404_), .Y(_187__0_) );
INVX1 INVX1_121 ( .A(w_C_1_), .Y(_408_) );
OR2X2 OR2X2_35 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_409_) );
NAND2X1 NAND2X1_78 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_410_) );
NAND3X1 NAND3X1_63 ( .A(_408_), .B(_410_), .C(_409_), .Y(_411_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_405_) );
AND2X2 AND2X2_50 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_406_) );
OAI21X1 OAI21X1_58 ( .A(_405_), .B(_406_), .C(w_C_1_), .Y(_407_) );
NAND2X1 NAND2X1_79 ( .A(_407_), .B(_411_), .Y(_187__1_) );
INVX1 INVX1_122 ( .A(w_C_2_), .Y(_415_) );
OR2X2 OR2X2_36 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_416_) );
NAND2X1 NAND2X1_80 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_417_) );
NAND3X1 NAND3X1_64 ( .A(_415_), .B(_417_), .C(_416_), .Y(_418_) );
NOR2X1 NOR2X1_71 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_412_) );
AND2X2 AND2X2_51 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_413_) );
OAI21X1 OAI21X1_59 ( .A(_412_), .B(_413_), .C(w_C_2_), .Y(_414_) );
NAND2X1 NAND2X1_81 ( .A(_414_), .B(_418_), .Y(_187__2_) );
INVX1 INVX1_123 ( .A(w_C_3_), .Y(_422_) );
OR2X2 OR2X2_37 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_423_) );
NAND2X1 NAND2X1_82 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_424_) );
NAND3X1 NAND3X1_65 ( .A(_422_), .B(_424_), .C(_423_), .Y(_425_) );
NOR2X1 NOR2X1_72 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_419_) );
AND2X2 AND2X2_52 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_420_) );
OAI21X1 OAI21X1_60 ( .A(_419_), .B(_420_), .C(w_C_3_), .Y(_421_) );
NAND2X1 NAND2X1_83 ( .A(_421_), .B(_425_), .Y(_187__3_) );
BUFX2 BUFX2_36 ( .A(w_C_34_), .Y(_187__34_) );
BUFX2 BUFX2_37 ( .A(1'b0), .Y(w_C_0_) );
endmodule
