module CSkipA_35bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_8_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_17_) );
OAI21X1 OAI21X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .C(1'b0), .Y(_18_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_19_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_20_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_21_) );
NAND3X1 NAND3X1_1 ( .A(_19_), .B(_20_), .C(_21_), .Y(_22_) );
OAI21X1 OAI21X1_2 ( .A(_18_), .B(_22_), .C(_17_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3_), .Y(_23_) );
OAI21X1 OAI21X1_3 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .C(1'b0), .Y(_24_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_25_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_26_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_27_) );
NAND3X1 NAND3X1_2 ( .A(_25_), .B(_26_), .C(_27_), .Y(_28_) );
OAI21X1 OAI21X1_4 ( .A(_24_), .B(_28_), .C(_23_), .Y(w_cout_2_) );
INVX1 INVX1_3 ( .A(_5_), .Y(_29_) );
OAI21X1 OAI21X1_5 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .C(1'b0), .Y(_30_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_31_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_32_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_33_) );
NAND3X1 NAND3X1_3 ( .A(_31_), .B(_32_), .C(_33_), .Y(_34_) );
OAI21X1 OAI21X1_6 ( .A(_30_), .B(_34_), .C(_29_), .Y(w_cout_3_) );
INVX1 INVX1_4 ( .A(_7_), .Y(_35_) );
OAI21X1 OAI21X1_7 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .C(1'b0), .Y(_36_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_37_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_38_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_39_) );
NAND3X1 NAND3X1_4 ( .A(_37_), .B(_38_), .C(_39_), .Y(_40_) );
OAI21X1 OAI21X1_8 ( .A(_36_), .B(_40_), .C(_35_), .Y(w_cout_4_) );
INVX1 INVX1_5 ( .A(_9_), .Y(_41_) );
OAI21X1 OAI21X1_9 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .C(1'b0), .Y(_42_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_43_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_44_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_45_) );
NAND3X1 NAND3X1_5 ( .A(_43_), .B(_44_), .C(_45_), .Y(_46_) );
OAI21X1 OAI21X1_10 ( .A(_42_), .B(_46_), .C(_41_), .Y(w_cout_5_) );
INVX1 INVX1_6 ( .A(_11_), .Y(_47_) );
OAI21X1 OAI21X1_11 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .C(1'b0), .Y(_48_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_49_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_50_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_51_) );
NAND3X1 NAND3X1_6 ( .A(_49_), .B(_50_), .C(_51_), .Y(_52_) );
OAI21X1 OAI21X1_12 ( .A(_48_), .B(_52_), .C(_47_), .Y(w_cout_6_) );
INVX1 INVX1_7 ( .A(_13_), .Y(_53_) );
OAI21X1 OAI21X1_13 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .C(1'b0), .Y(_54_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_55_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_56_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_57_) );
NAND3X1 NAND3X1_7 ( .A(_55_), .B(_56_), .C(_57_), .Y(_58_) );
OAI21X1 OAI21X1_14 ( .A(_54_), .B(_58_), .C(_53_), .Y(w_cout_7_) );
INVX1 INVX1_8 ( .A(_15_), .Y(_59_) );
OAI21X1 OAI21X1_15 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .C(1'b0), .Y(_60_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_61_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_62_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_63_) );
NAND3X1 NAND3X1_8 ( .A(_61_), .B(_62_), .C(_63_), .Y(_64_) );
OAI21X1 OAI21X1_16 ( .A(_60_), .B(_64_), .C(_59_), .Y(w_cout_8_) );
INVX1 INVX1_9 ( .A(skip0_cin_next), .Y(_68_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_69_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_70_) );
NAND3X1 NAND3X1_9 ( .A(_68_), .B(_70_), .C(_69_), .Y(_71_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_65_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_66_) );
OAI21X1 OAI21X1_17 ( .A(_65_), .B(_66_), .C(skip0_cin_next), .Y(_67_) );
NAND2X1 NAND2X1_2 ( .A(_67_), .B(_71_), .Y(_0__4_) );
OAI21X1 OAI21X1_18 ( .A(_68_), .B(_65_), .C(_70_), .Y(_2__1_) );
INVX1 INVX1_10 ( .A(_2__1_), .Y(_75_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_76_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_77_) );
NAND3X1 NAND3X1_10 ( .A(_75_), .B(_77_), .C(_76_), .Y(_78_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_72_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_73_) );
OAI21X1 OAI21X1_19 ( .A(_72_), .B(_73_), .C(_2__1_), .Y(_74_) );
NAND2X1 NAND2X1_4 ( .A(_74_), .B(_78_), .Y(_0__5_) );
OAI21X1 OAI21X1_20 ( .A(_75_), .B(_72_), .C(_77_), .Y(_2__2_) );
INVX1 INVX1_11 ( .A(_2__2_), .Y(_82_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_83_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_84_) );
NAND3X1 NAND3X1_11 ( .A(_82_), .B(_84_), .C(_83_), .Y(_85_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_79_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_80_) );
OAI21X1 OAI21X1_21 ( .A(_79_), .B(_80_), .C(_2__2_), .Y(_81_) );
NAND2X1 NAND2X1_6 ( .A(_81_), .B(_85_), .Y(_0__6_) );
OAI21X1 OAI21X1_22 ( .A(_82_), .B(_79_), .C(_84_), .Y(_2__3_) );
INVX1 INVX1_12 ( .A(_2__3_), .Y(_89_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_90_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_91_) );
NAND3X1 NAND3X1_12 ( .A(_89_), .B(_91_), .C(_90_), .Y(_92_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_86_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_87_) );
OAI21X1 OAI21X1_23 ( .A(_86_), .B(_87_), .C(_2__3_), .Y(_88_) );
NAND2X1 NAND2X1_8 ( .A(_88_), .B(_92_), .Y(_0__7_) );
OAI21X1 OAI21X1_24 ( .A(_89_), .B(_86_), .C(_91_), .Y(_1_) );
INVX1 INVX1_13 ( .A(w_cout_1_), .Y(_96_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_97_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_98_) );
NAND3X1 NAND3X1_13 ( .A(_96_), .B(_98_), .C(_97_), .Y(_99_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_93_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_94_) );
OAI21X1 OAI21X1_25 ( .A(_93_), .B(_94_), .C(w_cout_1_), .Y(_95_) );
NAND2X1 NAND2X1_10 ( .A(_95_), .B(_99_), .Y(_0__8_) );
OAI21X1 OAI21X1_26 ( .A(_96_), .B(_93_), .C(_98_), .Y(_4__1_) );
INVX1 INVX1_14 ( .A(_4__1_), .Y(_103_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_104_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_105_) );
NAND3X1 NAND3X1_14 ( .A(_103_), .B(_105_), .C(_104_), .Y(_106_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_100_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_101_) );
OAI21X1 OAI21X1_27 ( .A(_100_), .B(_101_), .C(_4__1_), .Y(_102_) );
NAND2X1 NAND2X1_12 ( .A(_102_), .B(_106_), .Y(_0__9_) );
OAI21X1 OAI21X1_28 ( .A(_103_), .B(_100_), .C(_105_), .Y(_4__2_) );
INVX1 INVX1_15 ( .A(_4__2_), .Y(_110_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_111_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_112_) );
NAND3X1 NAND3X1_15 ( .A(_110_), .B(_112_), .C(_111_), .Y(_113_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_107_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_108_) );
OAI21X1 OAI21X1_29 ( .A(_107_), .B(_108_), .C(_4__2_), .Y(_109_) );
NAND2X1 NAND2X1_14 ( .A(_109_), .B(_113_), .Y(_0__10_) );
OAI21X1 OAI21X1_30 ( .A(_110_), .B(_107_), .C(_112_), .Y(_4__3_) );
INVX1 INVX1_16 ( .A(_4__3_), .Y(_117_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_118_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_119_) );
NAND3X1 NAND3X1_16 ( .A(_117_), .B(_119_), .C(_118_), .Y(_120_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_114_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_115_) );
OAI21X1 OAI21X1_31 ( .A(_114_), .B(_115_), .C(_4__3_), .Y(_116_) );
NAND2X1 NAND2X1_16 ( .A(_116_), .B(_120_), .Y(_0__11_) );
OAI21X1 OAI21X1_32 ( .A(_117_), .B(_114_), .C(_119_), .Y(_3_) );
INVX1 INVX1_17 ( .A(w_cout_2_), .Y(_124_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_125_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_126_) );
NAND3X1 NAND3X1_17 ( .A(_124_), .B(_126_), .C(_125_), .Y(_127_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_121_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_122_) );
OAI21X1 OAI21X1_33 ( .A(_121_), .B(_122_), .C(w_cout_2_), .Y(_123_) );
NAND2X1 NAND2X1_18 ( .A(_123_), .B(_127_), .Y(_0__12_) );
OAI21X1 OAI21X1_34 ( .A(_124_), .B(_121_), .C(_126_), .Y(_6__1_) );
INVX1 INVX1_18 ( .A(_6__1_), .Y(_131_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_132_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_133_) );
NAND3X1 NAND3X1_18 ( .A(_131_), .B(_133_), .C(_132_), .Y(_134_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_128_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_129_) );
OAI21X1 OAI21X1_35 ( .A(_128_), .B(_129_), .C(_6__1_), .Y(_130_) );
NAND2X1 NAND2X1_20 ( .A(_130_), .B(_134_), .Y(_0__13_) );
OAI21X1 OAI21X1_36 ( .A(_131_), .B(_128_), .C(_133_), .Y(_6__2_) );
INVX1 INVX1_19 ( .A(_6__2_), .Y(_138_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_139_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_140_) );
NAND3X1 NAND3X1_19 ( .A(_138_), .B(_140_), .C(_139_), .Y(_141_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_135_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_136_) );
OAI21X1 OAI21X1_37 ( .A(_135_), .B(_136_), .C(_6__2_), .Y(_137_) );
NAND2X1 NAND2X1_22 ( .A(_137_), .B(_141_), .Y(_0__14_) );
OAI21X1 OAI21X1_38 ( .A(_138_), .B(_135_), .C(_140_), .Y(_6__3_) );
INVX1 INVX1_20 ( .A(_6__3_), .Y(_145_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_146_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_147_) );
NAND3X1 NAND3X1_20 ( .A(_145_), .B(_147_), .C(_146_), .Y(_148_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_142_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_143_) );
OAI21X1 OAI21X1_39 ( .A(_142_), .B(_143_), .C(_6__3_), .Y(_144_) );
NAND2X1 NAND2X1_24 ( .A(_144_), .B(_148_), .Y(_0__15_) );
OAI21X1 OAI21X1_40 ( .A(_145_), .B(_142_), .C(_147_), .Y(_5_) );
INVX1 INVX1_21 ( .A(w_cout_3_), .Y(_152_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_153_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_154_) );
NAND3X1 NAND3X1_21 ( .A(_152_), .B(_154_), .C(_153_), .Y(_155_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_149_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_150_) );
OAI21X1 OAI21X1_41 ( .A(_149_), .B(_150_), .C(w_cout_3_), .Y(_151_) );
NAND2X1 NAND2X1_26 ( .A(_151_), .B(_155_), .Y(_0__16_) );
OAI21X1 OAI21X1_42 ( .A(_152_), .B(_149_), .C(_154_), .Y(_8__1_) );
INVX1 INVX1_22 ( .A(_8__1_), .Y(_159_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_160_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_161_) );
NAND3X1 NAND3X1_22 ( .A(_159_), .B(_161_), .C(_160_), .Y(_162_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_156_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_157_) );
OAI21X1 OAI21X1_43 ( .A(_156_), .B(_157_), .C(_8__1_), .Y(_158_) );
NAND2X1 NAND2X1_28 ( .A(_158_), .B(_162_), .Y(_0__17_) );
OAI21X1 OAI21X1_44 ( .A(_159_), .B(_156_), .C(_161_), .Y(_8__2_) );
INVX1 INVX1_23 ( .A(_8__2_), .Y(_166_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_167_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_168_) );
NAND3X1 NAND3X1_23 ( .A(_166_), .B(_168_), .C(_167_), .Y(_169_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_163_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_164_) );
OAI21X1 OAI21X1_45 ( .A(_163_), .B(_164_), .C(_8__2_), .Y(_165_) );
NAND2X1 NAND2X1_30 ( .A(_165_), .B(_169_), .Y(_0__18_) );
OAI21X1 OAI21X1_46 ( .A(_166_), .B(_163_), .C(_168_), .Y(_8__3_) );
INVX1 INVX1_24 ( .A(_8__3_), .Y(_173_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_174_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_175_) );
NAND3X1 NAND3X1_24 ( .A(_173_), .B(_175_), .C(_174_), .Y(_176_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_170_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_171_) );
OAI21X1 OAI21X1_47 ( .A(_170_), .B(_171_), .C(_8__3_), .Y(_172_) );
NAND2X1 NAND2X1_32 ( .A(_172_), .B(_176_), .Y(_0__19_) );
OAI21X1 OAI21X1_48 ( .A(_173_), .B(_170_), .C(_175_), .Y(_7_) );
INVX1 INVX1_25 ( .A(w_cout_4_), .Y(_180_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_181_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_182_) );
NAND3X1 NAND3X1_25 ( .A(_180_), .B(_182_), .C(_181_), .Y(_183_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_177_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_178_) );
OAI21X1 OAI21X1_49 ( .A(_177_), .B(_178_), .C(w_cout_4_), .Y(_179_) );
NAND2X1 NAND2X1_34 ( .A(_179_), .B(_183_), .Y(_0__20_) );
OAI21X1 OAI21X1_50 ( .A(_180_), .B(_177_), .C(_182_), .Y(_10__1_) );
INVX1 INVX1_26 ( .A(_10__1_), .Y(_187_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_188_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_189_) );
NAND3X1 NAND3X1_26 ( .A(_187_), .B(_189_), .C(_188_), .Y(_190_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_184_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_185_) );
OAI21X1 OAI21X1_51 ( .A(_184_), .B(_185_), .C(_10__1_), .Y(_186_) );
NAND2X1 NAND2X1_36 ( .A(_186_), .B(_190_), .Y(_0__21_) );
OAI21X1 OAI21X1_52 ( .A(_187_), .B(_184_), .C(_189_), .Y(_10__2_) );
INVX1 INVX1_27 ( .A(_10__2_), .Y(_194_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_195_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_196_) );
NAND3X1 NAND3X1_27 ( .A(_194_), .B(_196_), .C(_195_), .Y(_197_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_191_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_192_) );
OAI21X1 OAI21X1_53 ( .A(_191_), .B(_192_), .C(_10__2_), .Y(_193_) );
NAND2X1 NAND2X1_38 ( .A(_193_), .B(_197_), .Y(_0__22_) );
OAI21X1 OAI21X1_54 ( .A(_194_), .B(_191_), .C(_196_), .Y(_10__3_) );
INVX1 INVX1_28 ( .A(_10__3_), .Y(_201_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_202_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_203_) );
NAND3X1 NAND3X1_28 ( .A(_201_), .B(_203_), .C(_202_), .Y(_204_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_198_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_199_) );
OAI21X1 OAI21X1_55 ( .A(_198_), .B(_199_), .C(_10__3_), .Y(_200_) );
NAND2X1 NAND2X1_40 ( .A(_200_), .B(_204_), .Y(_0__23_) );
OAI21X1 OAI21X1_56 ( .A(_201_), .B(_198_), .C(_203_), .Y(_9_) );
INVX1 INVX1_29 ( .A(w_cout_5_), .Y(_208_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_209_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_210_) );
NAND3X1 NAND3X1_29 ( .A(_208_), .B(_210_), .C(_209_), .Y(_211_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_205_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_206_) );
OAI21X1 OAI21X1_57 ( .A(_205_), .B(_206_), .C(w_cout_5_), .Y(_207_) );
NAND2X1 NAND2X1_42 ( .A(_207_), .B(_211_), .Y(_0__24_) );
OAI21X1 OAI21X1_58 ( .A(_208_), .B(_205_), .C(_210_), .Y(_12__1_) );
INVX1 INVX1_30 ( .A(_12__1_), .Y(_215_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_216_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_217_) );
NAND3X1 NAND3X1_30 ( .A(_215_), .B(_217_), .C(_216_), .Y(_218_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_212_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_213_) );
OAI21X1 OAI21X1_59 ( .A(_212_), .B(_213_), .C(_12__1_), .Y(_214_) );
NAND2X1 NAND2X1_44 ( .A(_214_), .B(_218_), .Y(_0__25_) );
OAI21X1 OAI21X1_60 ( .A(_215_), .B(_212_), .C(_217_), .Y(_12__2_) );
INVX1 INVX1_31 ( .A(_12__2_), .Y(_222_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_223_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_224_) );
NAND3X1 NAND3X1_31 ( .A(_222_), .B(_224_), .C(_223_), .Y(_225_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_219_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_220_) );
OAI21X1 OAI21X1_61 ( .A(_219_), .B(_220_), .C(_12__2_), .Y(_221_) );
NAND2X1 NAND2X1_46 ( .A(_221_), .B(_225_), .Y(_0__26_) );
OAI21X1 OAI21X1_62 ( .A(_222_), .B(_219_), .C(_224_), .Y(_12__3_) );
INVX1 INVX1_32 ( .A(_12__3_), .Y(_229_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_230_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_231_) );
NAND3X1 NAND3X1_32 ( .A(_229_), .B(_231_), .C(_230_), .Y(_232_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_226_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_227_) );
OAI21X1 OAI21X1_63 ( .A(_226_), .B(_227_), .C(_12__3_), .Y(_228_) );
NAND2X1 NAND2X1_48 ( .A(_228_), .B(_232_), .Y(_0__27_) );
OAI21X1 OAI21X1_64 ( .A(_229_), .B(_226_), .C(_231_), .Y(_11_) );
INVX1 INVX1_33 ( .A(w_cout_6_), .Y(_236_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_237_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_238_) );
NAND3X1 NAND3X1_33 ( .A(_236_), .B(_238_), .C(_237_), .Y(_239_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_233_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_234_) );
OAI21X1 OAI21X1_65 ( .A(_233_), .B(_234_), .C(w_cout_6_), .Y(_235_) );
NAND2X1 NAND2X1_50 ( .A(_235_), .B(_239_), .Y(_0__28_) );
OAI21X1 OAI21X1_66 ( .A(_236_), .B(_233_), .C(_238_), .Y(_14__1_) );
INVX1 INVX1_34 ( .A(_14__1_), .Y(_243_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_244_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_245_) );
NAND3X1 NAND3X1_34 ( .A(_243_), .B(_245_), .C(_244_), .Y(_246_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_240_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_241_) );
OAI21X1 OAI21X1_67 ( .A(_240_), .B(_241_), .C(_14__1_), .Y(_242_) );
NAND2X1 NAND2X1_52 ( .A(_242_), .B(_246_), .Y(_0__29_) );
OAI21X1 OAI21X1_68 ( .A(_243_), .B(_240_), .C(_245_), .Y(_14__2_) );
INVX1 INVX1_35 ( .A(_14__2_), .Y(_250_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_251_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_252_) );
NAND3X1 NAND3X1_35 ( .A(_250_), .B(_252_), .C(_251_), .Y(_253_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_247_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_248_) );
OAI21X1 OAI21X1_69 ( .A(_247_), .B(_248_), .C(_14__2_), .Y(_249_) );
NAND2X1 NAND2X1_54 ( .A(_249_), .B(_253_), .Y(_0__30_) );
OAI21X1 OAI21X1_70 ( .A(_250_), .B(_247_), .C(_252_), .Y(_14__3_) );
INVX1 INVX1_36 ( .A(_14__3_), .Y(_257_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_258_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_259_) );
NAND3X1 NAND3X1_36 ( .A(_257_), .B(_259_), .C(_258_), .Y(_260_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_254_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_255_) );
OAI21X1 OAI21X1_71 ( .A(_254_), .B(_255_), .C(_14__3_), .Y(_256_) );
NAND2X1 NAND2X1_56 ( .A(_256_), .B(_260_), .Y(_0__31_) );
OAI21X1 OAI21X1_72 ( .A(_257_), .B(_254_), .C(_259_), .Y(_13_) );
INVX1 INVX1_37 ( .A(w_cout_7_), .Y(_264_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_265_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_266_) );
NAND3X1 NAND3X1_37 ( .A(_264_), .B(_266_), .C(_265_), .Y(_267_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_261_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_262_) );
OAI21X1 OAI21X1_73 ( .A(_261_), .B(_262_), .C(w_cout_7_), .Y(_263_) );
NAND2X1 NAND2X1_58 ( .A(_263_), .B(_267_), .Y(_0__32_) );
OAI21X1 OAI21X1_74 ( .A(_264_), .B(_261_), .C(_266_), .Y(_16__1_) );
INVX1 INVX1_38 ( .A(_16__1_), .Y(_271_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_272_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_273_) );
NAND3X1 NAND3X1_38 ( .A(_271_), .B(_273_), .C(_272_), .Y(_274_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_268_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_269_) );
OAI21X1 OAI21X1_75 ( .A(_268_), .B(_269_), .C(_16__1_), .Y(_270_) );
NAND2X1 NAND2X1_60 ( .A(_270_), .B(_274_), .Y(_0__33_) );
OAI21X1 OAI21X1_76 ( .A(_271_), .B(_268_), .C(_273_), .Y(_16__2_) );
INVX1 INVX1_39 ( .A(_16__2_), .Y(_278_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_279_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_280_) );
NAND3X1 NAND3X1_39 ( .A(_278_), .B(_280_), .C(_279_), .Y(_281_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_275_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_276_) );
OAI21X1 OAI21X1_77 ( .A(_275_), .B(_276_), .C(_16__2_), .Y(_277_) );
NAND2X1 NAND2X1_62 ( .A(_277_), .B(_281_), .Y(_0__34_) );
OAI21X1 OAI21X1_78 ( .A(_278_), .B(_275_), .C(_280_), .Y(_16__3_) );
INVX1 INVX1_40 ( .A(_16__3_), .Y(_285_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_286_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_287_) );
NAND3X1 NAND3X1_40 ( .A(_285_), .B(_287_), .C(_286_), .Y(_288_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_282_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_283_) );
OAI21X1 OAI21X1_79 ( .A(_282_), .B(_283_), .C(_16__3_), .Y(_284_) );
NAND2X1 NAND2X1_64 ( .A(_284_), .B(_288_), .Y(_0__35_) );
OAI21X1 OAI21X1_80 ( .A(_285_), .B(_282_), .C(_287_), .Y(_15_) );
INVX1 INVX1_41 ( .A(1'b0), .Y(_292_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_293_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_294_) );
NAND3X1 NAND3X1_41 ( .A(_292_), .B(_294_), .C(_293_), .Y(_295_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_289_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_290_) );
OAI21X1 OAI21X1_81 ( .A(_289_), .B(_290_), .C(1'b0), .Y(_291_) );
NAND2X1 NAND2X1_66 ( .A(_291_), .B(_295_), .Y(_0__0_) );
OAI21X1 OAI21X1_82 ( .A(_292_), .B(_289_), .C(_294_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_42 ( .A(rca_inst_w_CARRY_1_), .Y(_299_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_300_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_301_) );
NAND3X1 NAND3X1_42 ( .A(_299_), .B(_301_), .C(_300_), .Y(_302_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_296_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_297_) );
OAI21X1 OAI21X1_83 ( .A(_296_), .B(_297_), .C(rca_inst_w_CARRY_1_), .Y(_298_) );
NAND2X1 NAND2X1_68 ( .A(_298_), .B(_302_), .Y(_0__1_) );
OAI21X1 OAI21X1_84 ( .A(_299_), .B(_296_), .C(_301_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_43 ( .A(rca_inst_w_CARRY_2_), .Y(_306_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_307_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_308_) );
NAND3X1 NAND3X1_43 ( .A(_306_), .B(_308_), .C(_307_), .Y(_309_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_303_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_304_) );
OAI21X1 OAI21X1_85 ( .A(_303_), .B(_304_), .C(rca_inst_w_CARRY_2_), .Y(_305_) );
NAND2X1 NAND2X1_70 ( .A(_305_), .B(_309_), .Y(_0__2_) );
OAI21X1 OAI21X1_86 ( .A(_306_), .B(_303_), .C(_308_), .Y(rca_inst_w_CARRY_3_) );
INVX1 INVX1_44 ( .A(rca_inst_w_CARRY_3_), .Y(_313_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_314_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_315_) );
NAND3X1 NAND3X1_44 ( .A(_313_), .B(_315_), .C(_314_), .Y(_316_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_310_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_311_) );
OAI21X1 OAI21X1_87 ( .A(_310_), .B(_311_), .C(rca_inst_w_CARRY_3_), .Y(_312_) );
NAND2X1 NAND2X1_72 ( .A(_312_), .B(_316_), .Y(_0__3_) );
OAI21X1 OAI21X1_88 ( .A(_313_), .B(_310_), .C(_315_), .Y(cout0) );
INVX1 INVX1_45 ( .A(cout0), .Y(_317_) );
OAI21X1 OAI21X1_89 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .C(1'b0), .Y(_318_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_319_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_320_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_321_) );
NAND3X1 NAND3X1_45 ( .A(_319_), .B(_320_), .C(_321_), .Y(_322_) );
OAI21X1 OAI21X1_90 ( .A(_318_), .B(_322_), .C(_317_), .Y(skip0_cin_next) );
BUFX2 BUFX2_38 ( .A(skip0_cin_next), .Y(_2__0_) );
BUFX2 BUFX2_39 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_40 ( .A(w_cout_1_), .Y(_4__0_) );
BUFX2 BUFX2_41 ( .A(_3_), .Y(_4__4_) );
BUFX2 BUFX2_42 ( .A(w_cout_2_), .Y(_6__0_) );
BUFX2 BUFX2_43 ( .A(_5_), .Y(_6__4_) );
BUFX2 BUFX2_44 ( .A(w_cout_3_), .Y(_8__0_) );
BUFX2 BUFX2_45 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_46 ( .A(w_cout_4_), .Y(_10__0_) );
BUFX2 BUFX2_47 ( .A(_9_), .Y(_10__4_) );
BUFX2 BUFX2_48 ( .A(w_cout_5_), .Y(_12__0_) );
BUFX2 BUFX2_49 ( .A(_11_), .Y(_12__4_) );
BUFX2 BUFX2_50 ( .A(w_cout_6_), .Y(_14__0_) );
BUFX2 BUFX2_51 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_52 ( .A(w_cout_7_), .Y(_16__0_) );
BUFX2 BUFX2_53 ( .A(_15_), .Y(_16__4_) );
BUFX2 BUFX2_54 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_55 ( .A(cout0), .Y(rca_inst_w_CARRY_4_) );
BUFX2 BUFX2_56 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
