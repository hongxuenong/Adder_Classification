module cla_48bit (i_add1, i_add2, o_result);

input [47:0] i_add1;
input [47:0] i_add2;
output [48:0] o_result;

wire vdd = 1'b1;
wire gnd = 1'b0;

NAND2X1 NAND2X1_1 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_294_) );
NAND3X1 NAND3X1_1 ( .A(_292_), .B(_294_), .C(_293_), .Y(_295_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_289_) );
AND2X2 AND2X2_1 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_290_) );
OAI21X1 OAI21X1_1 ( .A(_289_), .B(_290_), .C(w_C_6_), .Y(_291_) );
NAND2X1 NAND2X1_2 ( .A(_291_), .B(_295_), .Y(_274__6_) );
INVX1 INVX1_1 ( .A(w_C_7_), .Y(_299_) );
OR2X2 OR2X2_1 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_300_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_301_) );
NAND3X1 NAND3X1_2 ( .A(_299_), .B(_301_), .C(_300_), .Y(_302_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_296_) );
AND2X2 AND2X2_2 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_297_) );
OAI21X1 OAI21X1_2 ( .A(_296_), .B(_297_), .C(w_C_7_), .Y(_298_) );
NAND2X1 NAND2X1_4 ( .A(_298_), .B(_302_), .Y(_274__7_) );
INVX1 INVX1_2 ( .A(w_C_8_), .Y(_306_) );
OR2X2 OR2X2_2 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_307_) );
NAND2X1 NAND2X1_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_308_) );
NAND3X1 NAND3X1_3 ( .A(_306_), .B(_308_), .C(_307_), .Y(_309_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_303_) );
AND2X2 AND2X2_3 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_304_) );
OAI21X1 OAI21X1_3 ( .A(_303_), .B(_304_), .C(w_C_8_), .Y(_305_) );
NAND2X1 NAND2X1_6 ( .A(_305_), .B(_309_), .Y(_274__8_) );
INVX1 INVX1_3 ( .A(w_C_9_), .Y(_313_) );
OR2X2 OR2X2_3 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_314_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_315_) );
NAND3X1 NAND3X1_4 ( .A(_313_), .B(_315_), .C(_314_), .Y(_316_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_310_) );
AND2X2 AND2X2_4 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_311_) );
OAI21X1 OAI21X1_4 ( .A(_310_), .B(_311_), .C(w_C_9_), .Y(_312_) );
NAND2X1 NAND2X1_8 ( .A(_312_), .B(_316_), .Y(_274__9_) );
INVX1 INVX1_4 ( .A(w_C_10_), .Y(_320_) );
OR2X2 OR2X2_4 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_321_) );
NAND2X1 NAND2X1_9 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_322_) );
NAND3X1 NAND3X1_5 ( .A(_320_), .B(_322_), .C(_321_), .Y(_323_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_317_) );
AND2X2 AND2X2_5 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_318_) );
OAI21X1 OAI21X1_5 ( .A(_317_), .B(_318_), .C(w_C_10_), .Y(_319_) );
NAND2X1 NAND2X1_10 ( .A(_319_), .B(_323_), .Y(_274__10_) );
INVX1 INVX1_5 ( .A(w_C_11_), .Y(_327_) );
OR2X2 OR2X2_5 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_328_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_329_) );
NAND3X1 NAND3X1_6 ( .A(_327_), .B(_329_), .C(_328_), .Y(_330_) );
NOR2X1 NOR2X1_6 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_324_) );
AND2X2 AND2X2_6 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_325_) );
OAI21X1 OAI21X1_6 ( .A(_324_), .B(_325_), .C(w_C_11_), .Y(_326_) );
NAND2X1 NAND2X1_12 ( .A(_326_), .B(_330_), .Y(_274__11_) );
INVX1 INVX1_6 ( .A(w_C_12_), .Y(_334_) );
OR2X2 OR2X2_6 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_335_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_336_) );
NAND3X1 NAND3X1_7 ( .A(_334_), .B(_336_), .C(_335_), .Y(_337_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_331_) );
AND2X2 AND2X2_7 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_332_) );
OAI21X1 OAI21X1_7 ( .A(_331_), .B(_332_), .C(w_C_12_), .Y(_333_) );
NAND2X1 NAND2X1_14 ( .A(_333_), .B(_337_), .Y(_274__12_) );
INVX1 INVX1_7 ( .A(w_C_13_), .Y(_341_) );
OR2X2 OR2X2_7 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_342_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_343_) );
NAND3X1 NAND3X1_8 ( .A(_341_), .B(_343_), .C(_342_), .Y(_344_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_338_) );
AND2X2 AND2X2_8 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_339_) );
OAI21X1 OAI21X1_8 ( .A(_338_), .B(_339_), .C(w_C_13_), .Y(_340_) );
NAND2X1 NAND2X1_16 ( .A(_340_), .B(_344_), .Y(_274__13_) );
INVX1 INVX1_8 ( .A(w_C_14_), .Y(_348_) );
OR2X2 OR2X2_8 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_349_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_350_) );
NAND3X1 NAND3X1_9 ( .A(_348_), .B(_350_), .C(_349_), .Y(_351_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_345_) );
AND2X2 AND2X2_9 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_346_) );
OAI21X1 OAI21X1_9 ( .A(_345_), .B(_346_), .C(w_C_14_), .Y(_347_) );
NAND2X1 NAND2X1_18 ( .A(_347_), .B(_351_), .Y(_274__14_) );
INVX1 INVX1_9 ( .A(w_C_15_), .Y(_355_) );
OR2X2 OR2X2_9 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_356_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_357_) );
NAND3X1 NAND3X1_10 ( .A(_355_), .B(_357_), .C(_356_), .Y(_358_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_352_) );
AND2X2 AND2X2_10 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_353_) );
OAI21X1 OAI21X1_10 ( .A(_352_), .B(_353_), .C(w_C_15_), .Y(_354_) );
NAND2X1 NAND2X1_20 ( .A(_354_), .B(_358_), .Y(_274__15_) );
INVX1 INVX1_10 ( .A(w_C_16_), .Y(_362_) );
OR2X2 OR2X2_10 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_363_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_364_) );
NAND3X1 NAND3X1_11 ( .A(_362_), .B(_364_), .C(_363_), .Y(_365_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_359_) );
AND2X2 AND2X2_11 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_360_) );
OAI21X1 OAI21X1_11 ( .A(_359_), .B(_360_), .C(w_C_16_), .Y(_361_) );
NAND2X1 NAND2X1_22 ( .A(_361_), .B(_365_), .Y(_274__16_) );
INVX1 INVX1_11 ( .A(w_C_17_), .Y(_369_) );
OR2X2 OR2X2_11 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_370_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_371_) );
NAND3X1 NAND3X1_12 ( .A(_369_), .B(_371_), .C(_370_), .Y(_372_) );
NOR2X1 NOR2X1_12 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_366_) );
AND2X2 AND2X2_12 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_367_) );
OAI21X1 OAI21X1_12 ( .A(_366_), .B(_367_), .C(w_C_17_), .Y(_368_) );
NAND2X1 NAND2X1_24 ( .A(_368_), .B(_372_), .Y(_274__17_) );
INVX1 INVX1_12 ( .A(w_C_18_), .Y(_376_) );
OR2X2 OR2X2_12 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_377_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_378_) );
NAND3X1 NAND3X1_13 ( .A(_376_), .B(_378_), .C(_377_), .Y(_379_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_373_) );
AND2X2 AND2X2_13 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_374_) );
OAI21X1 OAI21X1_13 ( .A(_373_), .B(_374_), .C(w_C_18_), .Y(_375_) );
NAND2X1 NAND2X1_26 ( .A(_375_), .B(_379_), .Y(_274__18_) );
INVX1 INVX1_13 ( .A(w_C_19_), .Y(_383_) );
OR2X2 OR2X2_13 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_384_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_385_) );
NAND3X1 NAND3X1_14 ( .A(_383_), .B(_385_), .C(_384_), .Y(_386_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_380_) );
AND2X2 AND2X2_14 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_381_) );
OAI21X1 OAI21X1_14 ( .A(_380_), .B(_381_), .C(w_C_19_), .Y(_382_) );
NAND2X1 NAND2X1_28 ( .A(_382_), .B(_386_), .Y(_274__19_) );
INVX1 INVX1_14 ( .A(w_C_20_), .Y(_390_) );
OR2X2 OR2X2_14 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_391_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_392_) );
NAND3X1 NAND3X1_15 ( .A(_390_), .B(_392_), .C(_391_), .Y(_393_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_387_) );
AND2X2 AND2X2_15 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_388_) );
OAI21X1 OAI21X1_15 ( .A(_387_), .B(_388_), .C(w_C_20_), .Y(_389_) );
NAND2X1 NAND2X1_30 ( .A(_389_), .B(_393_), .Y(_274__20_) );
INVX1 INVX1_15 ( .A(w_C_21_), .Y(_397_) );
OR2X2 OR2X2_15 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_398_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_399_) );
NAND3X1 NAND3X1_16 ( .A(_397_), .B(_399_), .C(_398_), .Y(_400_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_394_) );
AND2X2 AND2X2_16 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_395_) );
OAI21X1 OAI21X1_16 ( .A(_394_), .B(_395_), .C(w_C_21_), .Y(_396_) );
NAND2X1 NAND2X1_32 ( .A(_396_), .B(_400_), .Y(_274__21_) );
INVX1 INVX1_16 ( .A(w_C_22_), .Y(_404_) );
OR2X2 OR2X2_16 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_405_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_406_) );
NAND3X1 NAND3X1_17 ( .A(_404_), .B(_406_), .C(_405_), .Y(_407_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_401_) );
AND2X2 AND2X2_17 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_402_) );
OAI21X1 OAI21X1_17 ( .A(_401_), .B(_402_), .C(w_C_22_), .Y(_403_) );
NAND2X1 NAND2X1_34 ( .A(_403_), .B(_407_), .Y(_274__22_) );
INVX1 INVX1_17 ( .A(w_C_23_), .Y(_411_) );
OR2X2 OR2X2_17 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_412_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_413_) );
NAND3X1 NAND3X1_18 ( .A(_411_), .B(_413_), .C(_412_), .Y(_414_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_408_) );
AND2X2 AND2X2_18 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_409_) );
OAI21X1 OAI21X1_18 ( .A(_408_), .B(_409_), .C(w_C_23_), .Y(_410_) );
NAND2X1 NAND2X1_36 ( .A(_410_), .B(_414_), .Y(_274__23_) );
INVX1 INVX1_18 ( .A(w_C_24_), .Y(_418_) );
OR2X2 OR2X2_18 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_419_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_420_) );
NAND3X1 NAND3X1_19 ( .A(_418_), .B(_420_), .C(_419_), .Y(_421_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_415_) );
AND2X2 AND2X2_19 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_416_) );
OAI21X1 OAI21X1_19 ( .A(_415_), .B(_416_), .C(w_C_24_), .Y(_417_) );
NAND2X1 NAND2X1_38 ( .A(_417_), .B(_421_), .Y(_274__24_) );
INVX1 INVX1_19 ( .A(w_C_25_), .Y(_425_) );
OR2X2 OR2X2_19 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_426_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_427_) );
NAND3X1 NAND3X1_20 ( .A(_425_), .B(_427_), .C(_426_), .Y(_428_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_422_) );
AND2X2 AND2X2_20 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_423_) );
OAI21X1 OAI21X1_20 ( .A(_422_), .B(_423_), .C(w_C_25_), .Y(_424_) );
NAND2X1 NAND2X1_40 ( .A(_424_), .B(_428_), .Y(_274__25_) );
INVX1 INVX1_20 ( .A(w_C_26_), .Y(_432_) );
OR2X2 OR2X2_20 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_433_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_434_) );
NAND3X1 NAND3X1_21 ( .A(_432_), .B(_434_), .C(_433_), .Y(_435_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_429_) );
AND2X2 AND2X2_21 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_430_) );
OAI21X1 OAI21X1_21 ( .A(_429_), .B(_430_), .C(w_C_26_), .Y(_431_) );
NAND2X1 NAND2X1_42 ( .A(_431_), .B(_435_), .Y(_274__26_) );
INVX1 INVX1_21 ( .A(w_C_27_), .Y(_439_) );
OR2X2 OR2X2_21 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_440_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_441_) );
NAND3X1 NAND3X1_22 ( .A(_439_), .B(_441_), .C(_440_), .Y(_442_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_436_) );
AND2X2 AND2X2_22 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_437_) );
OAI21X1 OAI21X1_22 ( .A(_436_), .B(_437_), .C(w_C_27_), .Y(_438_) );
NAND2X1 NAND2X1_44 ( .A(_438_), .B(_442_), .Y(_274__27_) );
INVX1 INVX1_22 ( .A(w_C_28_), .Y(_446_) );
OR2X2 OR2X2_22 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_447_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_448_) );
NAND3X1 NAND3X1_23 ( .A(_446_), .B(_448_), .C(_447_), .Y(_449_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_443_) );
AND2X2 AND2X2_23 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_444_) );
OAI21X1 OAI21X1_23 ( .A(_443_), .B(_444_), .C(w_C_28_), .Y(_445_) );
NAND2X1 NAND2X1_46 ( .A(_445_), .B(_449_), .Y(_274__28_) );
INVX1 INVX1_23 ( .A(w_C_29_), .Y(_453_) );
OR2X2 OR2X2_23 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_454_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_455_) );
NAND3X1 NAND3X1_24 ( .A(_453_), .B(_455_), .C(_454_), .Y(_456_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_450_) );
AND2X2 AND2X2_24 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_451_) );
OAI21X1 OAI21X1_24 ( .A(_450_), .B(_451_), .C(w_C_29_), .Y(_452_) );
NAND2X1 NAND2X1_48 ( .A(_452_), .B(_456_), .Y(_274__29_) );
INVX1 INVX1_24 ( .A(w_C_30_), .Y(_460_) );
OR2X2 OR2X2_24 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_461_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_462_) );
NAND3X1 NAND3X1_25 ( .A(_460_), .B(_462_), .C(_461_), .Y(_463_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_457_) );
AND2X2 AND2X2_25 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_458_) );
OAI21X1 OAI21X1_25 ( .A(_457_), .B(_458_), .C(w_C_30_), .Y(_459_) );
NAND2X1 NAND2X1_50 ( .A(_459_), .B(_463_), .Y(_274__30_) );
INVX1 INVX1_25 ( .A(w_C_31_), .Y(_467_) );
OR2X2 OR2X2_25 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_468_) );
NAND2X1 NAND2X1_51 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_469_) );
NAND3X1 NAND3X1_26 ( .A(_467_), .B(_469_), .C(_468_), .Y(_470_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_464_) );
AND2X2 AND2X2_26 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_465_) );
OAI21X1 OAI21X1_26 ( .A(_464_), .B(_465_), .C(w_C_31_), .Y(_466_) );
NAND2X1 NAND2X1_52 ( .A(_466_), .B(_470_), .Y(_274__31_) );
INVX1 INVX1_26 ( .A(w_C_32_), .Y(_474_) );
OR2X2 OR2X2_26 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_475_) );
NAND2X1 NAND2X1_53 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_476_) );
NAND3X1 NAND3X1_27 ( .A(_474_), .B(_476_), .C(_475_), .Y(_477_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_471_) );
AND2X2 AND2X2_27 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_472_) );
OAI21X1 OAI21X1_27 ( .A(_471_), .B(_472_), .C(w_C_32_), .Y(_473_) );
NAND2X1 NAND2X1_54 ( .A(_473_), .B(_477_), .Y(_274__32_) );
INVX1 INVX1_27 ( .A(w_C_33_), .Y(_481_) );
OR2X2 OR2X2_27 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_482_) );
NAND2X1 NAND2X1_55 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_483_) );
NAND3X1 NAND3X1_28 ( .A(_481_), .B(_483_), .C(_482_), .Y(_484_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_478_) );
AND2X2 AND2X2_28 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_479_) );
OAI21X1 OAI21X1_28 ( .A(_478_), .B(_479_), .C(w_C_33_), .Y(_480_) );
NAND2X1 NAND2X1_56 ( .A(_480_), .B(_484_), .Y(_274__33_) );
INVX1 INVX1_28 ( .A(w_C_34_), .Y(_488_) );
OR2X2 OR2X2_28 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_489_) );
NAND2X1 NAND2X1_57 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_490_) );
NAND3X1 NAND3X1_29 ( .A(_488_), .B(_490_), .C(_489_), .Y(_491_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_485_) );
AND2X2 AND2X2_29 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_486_) );
OAI21X1 OAI21X1_29 ( .A(_485_), .B(_486_), .C(w_C_34_), .Y(_487_) );
NAND2X1 NAND2X1_58 ( .A(_487_), .B(_491_), .Y(_274__34_) );
INVX1 INVX1_29 ( .A(w_C_35_), .Y(_495_) );
OR2X2 OR2X2_29 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_496_) );
NAND2X1 NAND2X1_59 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_497_) );
NAND3X1 NAND3X1_30 ( .A(_495_), .B(_497_), .C(_496_), .Y(_498_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_492_) );
AND2X2 AND2X2_30 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_493_) );
OAI21X1 OAI21X1_30 ( .A(_492_), .B(_493_), .C(w_C_35_), .Y(_494_) );
NAND2X1 NAND2X1_60 ( .A(_494_), .B(_498_), .Y(_274__35_) );
INVX1 INVX1_30 ( .A(w_C_36_), .Y(_502_) );
OR2X2 OR2X2_30 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_503_) );
NAND2X1 NAND2X1_61 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_504_) );
NAND3X1 NAND3X1_31 ( .A(_502_), .B(_504_), .C(_503_), .Y(_505_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_499_) );
AND2X2 AND2X2_31 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_500_) );
OAI21X1 OAI21X1_31 ( .A(_499_), .B(_500_), .C(w_C_36_), .Y(_501_) );
NAND2X1 NAND2X1_62 ( .A(_501_), .B(_505_), .Y(_274__36_) );
INVX1 INVX1_31 ( .A(w_C_37_), .Y(_509_) );
OR2X2 OR2X2_31 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_510_) );
NAND2X1 NAND2X1_63 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_511_) );
NAND3X1 NAND3X1_32 ( .A(_509_), .B(_511_), .C(_510_), .Y(_512_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_506_) );
AND2X2 AND2X2_32 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_507_) );
OAI21X1 OAI21X1_32 ( .A(_506_), .B(_507_), .C(w_C_37_), .Y(_508_) );
NAND2X1 NAND2X1_64 ( .A(_508_), .B(_512_), .Y(_274__37_) );
INVX1 INVX1_32 ( .A(w_C_38_), .Y(_516_) );
OR2X2 OR2X2_32 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_517_) );
NAND2X1 NAND2X1_65 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_518_) );
NAND3X1 NAND3X1_33 ( .A(_516_), .B(_518_), .C(_517_), .Y(_519_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_513_) );
AND2X2 AND2X2_33 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_514_) );
OAI21X1 OAI21X1_33 ( .A(_513_), .B(_514_), .C(w_C_38_), .Y(_515_) );
NAND2X1 NAND2X1_66 ( .A(_515_), .B(_519_), .Y(_274__38_) );
INVX1 INVX1_33 ( .A(w_C_39_), .Y(_523_) );
OR2X2 OR2X2_33 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_524_) );
NAND2X1 NAND2X1_67 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_525_) );
NAND3X1 NAND3X1_34 ( .A(_523_), .B(_525_), .C(_524_), .Y(_526_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_520_) );
AND2X2 AND2X2_34 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_521_) );
OAI21X1 OAI21X1_34 ( .A(_520_), .B(_521_), .C(w_C_39_), .Y(_522_) );
NAND2X1 NAND2X1_68 ( .A(_522_), .B(_526_), .Y(_274__39_) );
INVX1 INVX1_34 ( .A(w_C_40_), .Y(_530_) );
OR2X2 OR2X2_34 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_531_) );
NAND2X1 NAND2X1_69 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_532_) );
NAND3X1 NAND3X1_35 ( .A(_530_), .B(_532_), .C(_531_), .Y(_533_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_527_) );
AND2X2 AND2X2_35 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_528_) );
OAI21X1 OAI21X1_35 ( .A(_527_), .B(_528_), .C(w_C_40_), .Y(_529_) );
NAND2X1 NAND2X1_70 ( .A(_529_), .B(_533_), .Y(_274__40_) );
INVX1 INVX1_35 ( .A(w_C_41_), .Y(_537_) );
OR2X2 OR2X2_35 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_538_) );
NAND2X1 NAND2X1_71 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_539_) );
NAND3X1 NAND3X1_36 ( .A(_537_), .B(_539_), .C(_538_), .Y(_540_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_534_) );
AND2X2 AND2X2_36 ( .A(i_add2[41]), .B(i_add1[41]), .Y(_535_) );
OAI21X1 OAI21X1_36 ( .A(_534_), .B(_535_), .C(w_C_41_), .Y(_536_) );
NAND2X1 NAND2X1_72 ( .A(_536_), .B(_540_), .Y(_274__41_) );
INVX1 INVX1_36 ( .A(w_C_42_), .Y(_544_) );
OR2X2 OR2X2_36 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_545_) );
NAND2X1 NAND2X1_73 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_546_) );
NAND3X1 NAND3X1_37 ( .A(_544_), .B(_546_), .C(_545_), .Y(_547_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_541_) );
AND2X2 AND2X2_37 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_542_) );
OAI21X1 OAI21X1_37 ( .A(_541_), .B(_542_), .C(w_C_42_), .Y(_543_) );
NAND2X1 NAND2X1_74 ( .A(_543_), .B(_547_), .Y(_274__42_) );
INVX1 INVX1_37 ( .A(w_C_43_), .Y(_551_) );
OR2X2 OR2X2_37 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_552_) );
NAND2X1 NAND2X1_75 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_553_) );
NAND3X1 NAND3X1_38 ( .A(_551_), .B(_553_), .C(_552_), .Y(_554_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_548_) );
AND2X2 AND2X2_38 ( .A(i_add2[43]), .B(i_add1[43]), .Y(_549_) );
OAI21X1 OAI21X1_38 ( .A(_548_), .B(_549_), .C(w_C_43_), .Y(_550_) );
NAND2X1 NAND2X1_76 ( .A(_550_), .B(_554_), .Y(_274__43_) );
INVX1 INVX1_38 ( .A(w_C_44_), .Y(_558_) );
OR2X2 OR2X2_38 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_559_) );
NAND2X1 NAND2X1_77 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_560_) );
NAND3X1 NAND3X1_39 ( .A(_558_), .B(_560_), .C(_559_), .Y(_561_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_555_) );
AND2X2 AND2X2_39 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_556_) );
OAI21X1 OAI21X1_39 ( .A(_555_), .B(_556_), .C(w_C_44_), .Y(_557_) );
NAND2X1 NAND2X1_78 ( .A(_557_), .B(_561_), .Y(_274__44_) );
INVX1 INVX1_39 ( .A(w_C_45_), .Y(_565_) );
OR2X2 OR2X2_39 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_566_) );
NAND2X1 NAND2X1_79 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_567_) );
NAND3X1 NAND3X1_40 ( .A(_565_), .B(_567_), .C(_566_), .Y(_568_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_562_) );
AND2X2 AND2X2_40 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_563_) );
OAI21X1 OAI21X1_40 ( .A(_562_), .B(_563_), .C(w_C_45_), .Y(_564_) );
NAND2X1 NAND2X1_80 ( .A(_564_), .B(_568_), .Y(_274__45_) );
INVX1 INVX1_40 ( .A(w_C_46_), .Y(_572_) );
OR2X2 OR2X2_40 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_573_) );
NAND2X1 NAND2X1_81 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_574_) );
NAND3X1 NAND3X1_41 ( .A(_572_), .B(_574_), .C(_573_), .Y(_575_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_569_) );
AND2X2 AND2X2_41 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_570_) );
OAI21X1 OAI21X1_41 ( .A(_569_), .B(_570_), .C(w_C_46_), .Y(_571_) );
NAND2X1 NAND2X1_82 ( .A(_571_), .B(_575_), .Y(_274__46_) );
INVX1 INVX1_41 ( .A(w_C_47_), .Y(_579_) );
OR2X2 OR2X2_41 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_580_) );
NAND2X1 NAND2X1_83 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_581_) );
NAND3X1 NAND3X1_42 ( .A(_579_), .B(_581_), .C(_580_), .Y(_582_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_576_) );
AND2X2 AND2X2_42 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_577_) );
OAI21X1 OAI21X1_42 ( .A(_576_), .B(_577_), .C(w_C_47_), .Y(_578_) );
NAND2X1 NAND2X1_84 ( .A(_578_), .B(_582_), .Y(_274__47_) );
INVX1 INVX1_42 ( .A(gnd), .Y(_586_) );
OR2X2 OR2X2_42 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_587_) );
NAND2X1 NAND2X1_85 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_588_) );
NAND3X1 NAND3X1_43 ( .A(_586_), .B(_588_), .C(_587_), .Y(_589_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_583_) );
AND2X2 AND2X2_43 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_584_) );
OAI21X1 OAI21X1_43 ( .A(_583_), .B(_584_), .C(gnd), .Y(_585_) );
NAND2X1 NAND2X1_86 ( .A(_585_), .B(_589_), .Y(_274__0_) );
INVX1 INVX1_43 ( .A(w_C_1_), .Y(_593_) );
OR2X2 OR2X2_43 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_594_) );
NAND2X1 NAND2X1_87 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_595_) );
NAND3X1 NAND3X1_44 ( .A(_593_), .B(_595_), .C(_594_), .Y(_596_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_590_) );
AND2X2 AND2X2_44 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_591_) );
OAI21X1 OAI21X1_44 ( .A(_590_), .B(_591_), .C(w_C_1_), .Y(_592_) );
NAND2X1 NAND2X1_88 ( .A(_592_), .B(_596_), .Y(_274__1_) );
INVX1 INVX1_44 ( .A(w_C_2_), .Y(_600_) );
OR2X2 OR2X2_44 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_601_) );
NAND2X1 NAND2X1_89 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_602_) );
NAND3X1 NAND3X1_45 ( .A(_600_), .B(_602_), .C(_601_), .Y(_603_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_597_) );
AND2X2 AND2X2_45 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_598_) );
OAI21X1 OAI21X1_45 ( .A(_597_), .B(_598_), .C(w_C_2_), .Y(_599_) );
NAND2X1 NAND2X1_90 ( .A(_599_), .B(_603_), .Y(_274__2_) );
INVX1 INVX1_45 ( .A(w_C_3_), .Y(_607_) );
OR2X2 OR2X2_45 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_608_) );
NAND2X1 NAND2X1_91 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_609_) );
NAND3X1 NAND3X1_46 ( .A(_607_), .B(_609_), .C(_608_), .Y(_610_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_604_) );
AND2X2 AND2X2_46 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_605_) );
OAI21X1 OAI21X1_46 ( .A(_604_), .B(_605_), .C(w_C_3_), .Y(_606_) );
NAND2X1 NAND2X1_92 ( .A(_606_), .B(_610_), .Y(_274__3_) );
INVX1 INVX1_46 ( .A(_215_), .Y(w_C_37_) );
INVX1 INVX1_47 ( .A(i_add2[37]), .Y(_216_) );
INVX1 INVX1_48 ( .A(i_add1[37]), .Y(_217_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_218_) );
INVX1 INVX1_49 ( .A(_218_), .Y(_219_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[37]), .B(i_add1[37]), .Y(_220_) );
INVX1 INVX1_50 ( .A(_220_), .Y(_221_) );
NAND3X1 NAND3X1_47 ( .A(_219_), .B(_221_), .C(_214_), .Y(_222_) );
OAI21X1 OAI21X1_47 ( .A(_216_), .B(_217_), .C(_222_), .Y(w_C_38_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_223_) );
INVX1 INVX1_51 ( .A(_223_), .Y(_224_) );
NOR2X1 NOR2X1_50 ( .A(_216_), .B(_217_), .Y(_225_) );
INVX1 INVX1_52 ( .A(_225_), .Y(_226_) );
NAND2X1 NAND2X1_93 ( .A(i_add2[38]), .B(i_add1[38]), .Y(_227_) );
NAND3X1 NAND3X1_48 ( .A(_226_), .B(_227_), .C(_222_), .Y(_228_) );
AND2X2 AND2X2_47 ( .A(_228_), .B(_224_), .Y(w_C_39_) );
INVX1 INVX1_53 ( .A(i_add2[39]), .Y(_229_) );
INVX1 INVX1_54 ( .A(i_add1[39]), .Y(_230_) );
NAND2X1 NAND2X1_94 ( .A(_229_), .B(_230_), .Y(_231_) );
NAND3X1 NAND3X1_49 ( .A(_224_), .B(_231_), .C(_228_), .Y(_232_) );
OAI21X1 OAI21X1_48 ( .A(_229_), .B(_230_), .C(_232_), .Y(w_C_40_) );
INVX1 INVX1_55 ( .A(i_add2[40]), .Y(_233_) );
INVX1 INVX1_56 ( .A(i_add1[40]), .Y(_234_) );
OAI21X1 OAI21X1_49 ( .A(i_add2[40]), .B(i_add1[40]), .C(w_C_40_), .Y(_235_) );
OAI21X1 OAI21X1_50 ( .A(_233_), .B(_234_), .C(_235_), .Y(w_C_41_) );
INVX1 INVX1_57 ( .A(i_add2[41]), .Y(_236_) );
INVX1 INVX1_58 ( .A(i_add1[41]), .Y(_237_) );
NOR2X1 NOR2X1_51 ( .A(_236_), .B(_237_), .Y(_238_) );
OR2X2 OR2X2_46 ( .A(w_C_41_), .B(_238_), .Y(_239_) );
OAI21X1 OAI21X1_51 ( .A(i_add2[41]), .B(i_add1[41]), .C(_239_), .Y(_240_) );
INVX1 INVX1_59 ( .A(_240_), .Y(w_C_42_) );
INVX1 INVX1_60 ( .A(_238_), .Y(_241_) );
NAND2X1 NAND2X1_95 ( .A(_233_), .B(_234_), .Y(_242_) );
NAND2X1 NAND2X1_96 ( .A(i_add2[39]), .B(i_add1[39]), .Y(_243_) );
NAND2X1 NAND2X1_97 ( .A(i_add2[40]), .B(i_add1[40]), .Y(_244_) );
NAND3X1 NAND3X1_50 ( .A(_243_), .B(_244_), .C(_232_), .Y(_245_) );
NAND2X1 NAND2X1_98 ( .A(_236_), .B(_237_), .Y(_246_) );
NAND3X1 NAND3X1_51 ( .A(_242_), .B(_246_), .C(_245_), .Y(_247_) );
NAND2X1 NAND2X1_99 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_248_) );
NAND3X1 NAND3X1_52 ( .A(_241_), .B(_248_), .C(_247_), .Y(_249_) );
OAI21X1 OAI21X1_52 ( .A(i_add2[42]), .B(i_add1[42]), .C(_249_), .Y(_250_) );
INVX1 INVX1_61 ( .A(_250_), .Y(w_C_43_) );
INVX1 INVX1_62 ( .A(i_add2[43]), .Y(_251_) );
INVX1 INVX1_63 ( .A(i_add1[43]), .Y(_252_) );
OAI21X1 OAI21X1_53 ( .A(_251_), .B(_252_), .C(_250_), .Y(_253_) );
OAI21X1 OAI21X1_54 ( .A(i_add2[43]), .B(i_add1[43]), .C(_253_), .Y(_254_) );
INVX1 INVX1_64 ( .A(_254_), .Y(w_C_44_) );
NAND2X1 NAND2X1_100 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_255_) );
NOR2X1 NOR2X1_52 ( .A(i_add2[44]), .B(i_add1[44]), .Y(_256_) );
OAI21X1 OAI21X1_55 ( .A(_256_), .B(_254_), .C(_255_), .Y(w_C_45_) );
NAND2X1 NAND2X1_101 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_257_) );
INVX1 INVX1_65 ( .A(_256_), .Y(_258_) );
NOR2X1 NOR2X1_53 ( .A(_251_), .B(_252_), .Y(_259_) );
INVX1 INVX1_66 ( .A(_259_), .Y(_260_) );
NOR2X1 NOR2X1_54 ( .A(i_add2[42]), .B(i_add1[42]), .Y(_261_) );
INVX1 INVX1_67 ( .A(_261_), .Y(_262_) );
NAND2X1 NAND2X1_102 ( .A(_251_), .B(_252_), .Y(_263_) );
NAND3X1 NAND3X1_53 ( .A(_262_), .B(_263_), .C(_249_), .Y(_264_) );
NAND3X1 NAND3X1_54 ( .A(_260_), .B(_255_), .C(_264_), .Y(_265_) );
OR2X2 OR2X2_47 ( .A(i_add2[45]), .B(i_add1[45]), .Y(_266_) );
NAND3X1 NAND3X1_55 ( .A(_258_), .B(_266_), .C(_265_), .Y(_267_) );
NAND2X1 NAND2X1_103 ( .A(_257_), .B(_267_), .Y(w_C_46_) );
OR2X2 OR2X2_48 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_268_) );
NAND2X1 NAND2X1_104 ( .A(i_add2[46]), .B(i_add1[46]), .Y(_269_) );
NAND3X1 NAND3X1_56 ( .A(_257_), .B(_269_), .C(_267_), .Y(_270_) );
AND2X2 AND2X2_48 ( .A(_270_), .B(_268_), .Y(w_C_47_) );
NAND2X1 NAND2X1_105 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_271_) );
OR2X2 OR2X2_49 ( .A(i_add2[47]), .B(i_add1[47]), .Y(_272_) );
NAND3X1 NAND3X1_57 ( .A(_268_), .B(_272_), .C(_270_), .Y(_273_) );
NAND2X1 NAND2X1_106 ( .A(_271_), .B(_273_), .Y(w_C_48_) );
NAND2X1 NAND2X1_107 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_68 ( .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_55 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_56 ( .A(_1_), .B(_2_), .Y(w_C_2_) );
INVX1 INVX1_69 ( .A(i_add2[2]), .Y(_3_) );
INVX1 INVX1_70 ( .A(i_add1[2]), .Y(_4_) );
NAND2X1 NAND2X1_108 ( .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_109 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
OAI21X1 OAI21X1_56 ( .A(_1_), .B(_2_), .C(_6_), .Y(_7_) );
AND2X2 AND2X2_49 ( .A(_7_), .B(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_110 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
OR2X2 OR2X2_50 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_9_) );
NAND3X1 NAND3X1_58 ( .A(_5_), .B(_9_), .C(_7_), .Y(_10_) );
NAND2X1 NAND2X1_111 ( .A(_8_), .B(_10_), .Y(w_C_4_) );
NOR2X1 NOR2X1_57 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_11_) );
INVX1 INVX1_71 ( .A(_11_), .Y(_12_) );
NAND2X1 NAND2X1_112 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
NAND3X1 NAND3X1_59 ( .A(_8_), .B(_13_), .C(_10_), .Y(_14_) );
AND2X2 AND2X2_50 ( .A(_14_), .B(_12_), .Y(w_C_5_) );
AND2X2 AND2X2_51 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_15_) );
INVX1 INVX1_72 ( .A(_15_), .Y(_16_) );
NOR2X1 NOR2X1_58 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_17_) );
INVX1 INVX1_73 ( .A(_17_), .Y(_18_) );
NAND3X1 NAND3X1_60 ( .A(_12_), .B(_18_), .C(_14_), .Y(_19_) );
AND2X2 AND2X2_52 ( .A(_19_), .B(_16_), .Y(_20_) );
INVX1 INVX1_74 ( .A(_20_), .Y(w_C_6_) );
AND2X2 AND2X2_53 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_21_) );
INVX1 INVX1_75 ( .A(_21_), .Y(_22_) );
NOR2X1 NOR2X1_59 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_23_) );
OAI21X1 OAI21X1_57 ( .A(_23_), .B(_20_), .C(_22_), .Y(w_C_7_) );
AND2X2 AND2X2_54 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_24_) );
INVX1 INVX1_76 ( .A(_24_), .Y(_25_) );
INVX1 INVX1_77 ( .A(_23_), .Y(_26_) );
NAND3X1 NAND3X1_61 ( .A(_16_), .B(_22_), .C(_19_), .Y(_27_) );
NOR2X1 NOR2X1_60 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_28_) );
INVX1 INVX1_78 ( .A(_28_), .Y(_29_) );
NAND3X1 NAND3X1_62 ( .A(_26_), .B(_29_), .C(_27_), .Y(_30_) );
AND2X2 AND2X2_55 ( .A(_30_), .B(_25_), .Y(_31_) );
INVX1 INVX1_79 ( .A(_31_), .Y(w_C_8_) );
AND2X2 AND2X2_56 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_32_) );
INVX1 INVX1_80 ( .A(_32_), .Y(_33_) );
NOR2X1 NOR2X1_61 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_34_) );
OAI21X1 OAI21X1_58 ( .A(_34_), .B(_31_), .C(_33_), .Y(w_C_9_) );
AND2X2 AND2X2_57 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_35_) );
INVX1 INVX1_81 ( .A(_35_), .Y(_36_) );
INVX1 INVX1_82 ( .A(_34_), .Y(_37_) );
NAND3X1 NAND3X1_63 ( .A(_25_), .B(_33_), .C(_30_), .Y(_38_) );
NOR2X1 NOR2X1_62 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_39_) );
INVX1 INVX1_83 ( .A(_39_), .Y(_40_) );
NAND3X1 NAND3X1_64 ( .A(_37_), .B(_40_), .C(_38_), .Y(_41_) );
AND2X2 AND2X2_58 ( .A(_41_), .B(_36_), .Y(_42_) );
INVX1 INVX1_84 ( .A(_42_), .Y(w_C_10_) );
AND2X2 AND2X2_59 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_43_) );
INVX1 INVX1_85 ( .A(_43_), .Y(_44_) );
NAND3X1 NAND3X1_65 ( .A(_36_), .B(_44_), .C(_41_), .Y(_45_) );
OAI21X1 OAI21X1_59 ( .A(i_add2[10]), .B(i_add1[10]), .C(_45_), .Y(_46_) );
INVX1 INVX1_86 ( .A(_46_), .Y(w_C_11_) );
INVX1 INVX1_87 ( .A(i_add2[11]), .Y(_47_) );
INVX1 INVX1_88 ( .A(i_add1[11]), .Y(_48_) );
NOR2X1 NOR2X1_63 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_49_) );
INVX1 INVX1_89 ( .A(_49_), .Y(_50_) );
NOR2X1 NOR2X1_64 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_51_) );
INVX1 INVX1_90 ( .A(_51_), .Y(_52_) );
NAND3X1 NAND3X1_66 ( .A(_50_), .B(_52_), .C(_45_), .Y(_53_) );
OAI21X1 OAI21X1_60 ( .A(_47_), .B(_48_), .C(_53_), .Y(w_C_12_) );
NOR2X1 NOR2X1_65 ( .A(_47_), .B(_48_), .Y(_54_) );
INVX1 INVX1_91 ( .A(_54_), .Y(_55_) );
AND2X2 AND2X2_60 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_56_) );
INVX1 INVX1_92 ( .A(_56_), .Y(_57_) );
NAND3X1 NAND3X1_67 ( .A(_55_), .B(_57_), .C(_53_), .Y(_58_) );
OAI21X1 OAI21X1_61 ( .A(i_add2[12]), .B(i_add1[12]), .C(_58_), .Y(_59_) );
INVX1 INVX1_93 ( .A(_59_), .Y(w_C_13_) );
INVX1 INVX1_94 ( .A(i_add2[13]), .Y(_60_) );
INVX1 INVX1_95 ( .A(i_add1[13]), .Y(_61_) );
NOR2X1 NOR2X1_66 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_62_) );
INVX1 INVX1_96 ( .A(_62_), .Y(_63_) );
NOR2X1 NOR2X1_67 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_64_) );
INVX1 INVX1_97 ( .A(_64_), .Y(_65_) );
NAND3X1 NAND3X1_68 ( .A(_63_), .B(_65_), .C(_58_), .Y(_66_) );
OAI21X1 OAI21X1_62 ( .A(_60_), .B(_61_), .C(_66_), .Y(w_C_14_) );
NOR2X1 NOR2X1_68 ( .A(_60_), .B(_61_), .Y(_67_) );
INVX1 INVX1_98 ( .A(_67_), .Y(_68_) );
AND2X2 AND2X2_61 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_69_) );
INVX1 INVX1_99 ( .A(_69_), .Y(_70_) );
NAND3X1 NAND3X1_69 ( .A(_68_), .B(_70_), .C(_66_), .Y(_71_) );
OAI21X1 OAI21X1_63 ( .A(i_add2[14]), .B(i_add1[14]), .C(_71_), .Y(_72_) );
INVX1 INVX1_100 ( .A(_72_), .Y(w_C_15_) );
INVX1 INVX1_101 ( .A(i_add2[15]), .Y(_73_) );
INVX1 INVX1_102 ( .A(i_add1[15]), .Y(_74_) );
NOR2X1 NOR2X1_69 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_75_) );
INVX1 INVX1_103 ( .A(_75_), .Y(_76_) );
NOR2X1 NOR2X1_70 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_77_) );
INVX1 INVX1_104 ( .A(_77_), .Y(_78_) );
NAND3X1 NAND3X1_70 ( .A(_76_), .B(_78_), .C(_71_), .Y(_79_) );
OAI21X1 OAI21X1_64 ( .A(_73_), .B(_74_), .C(_79_), .Y(w_C_16_) );
NOR2X1 NOR2X1_71 ( .A(_73_), .B(_74_), .Y(_80_) );
INVX1 INVX1_105 ( .A(_80_), .Y(_81_) );
AND2X2 AND2X2_62 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_82_) );
INVX1 INVX1_106 ( .A(_82_), .Y(_83_) );
NAND3X1 NAND3X1_71 ( .A(_81_), .B(_83_), .C(_79_), .Y(_84_) );
OAI21X1 OAI21X1_65 ( .A(i_add2[16]), .B(i_add1[16]), .C(_84_), .Y(_85_) );
INVX1 INVX1_107 ( .A(_85_), .Y(w_C_17_) );
INVX1 INVX1_108 ( .A(i_add2[17]), .Y(_86_) );
INVX1 INVX1_109 ( .A(i_add1[17]), .Y(_87_) );
NOR2X1 NOR2X1_72 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_88_) );
INVX1 INVX1_110 ( .A(_88_), .Y(_89_) );
NOR2X1 NOR2X1_73 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_90_) );
INVX1 INVX1_111 ( .A(_90_), .Y(_91_) );
NAND3X1 NAND3X1_72 ( .A(_89_), .B(_91_), .C(_84_), .Y(_92_) );
OAI21X1 OAI21X1_66 ( .A(_86_), .B(_87_), .C(_92_), .Y(w_C_18_) );
NOR2X1 NOR2X1_74 ( .A(_86_), .B(_87_), .Y(_93_) );
INVX1 INVX1_112 ( .A(_93_), .Y(_94_) );
AND2X2 AND2X2_63 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_95_) );
INVX1 INVX1_113 ( .A(_95_), .Y(_96_) );
NAND3X1 NAND3X1_73 ( .A(_94_), .B(_96_), .C(_92_), .Y(_97_) );
OAI21X1 OAI21X1_67 ( .A(i_add2[18]), .B(i_add1[18]), .C(_97_), .Y(_98_) );
INVX1 INVX1_114 ( .A(_98_), .Y(w_C_19_) );
INVX1 INVX1_115 ( .A(i_add2[19]), .Y(_99_) );
INVX1 INVX1_116 ( .A(i_add1[19]), .Y(_100_) );
NOR2X1 NOR2X1_75 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_101_) );
INVX1 INVX1_117 ( .A(_101_), .Y(_102_) );
NOR2X1 NOR2X1_76 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_103_) );
INVX1 INVX1_118 ( .A(_103_), .Y(_104_) );
NAND3X1 NAND3X1_74 ( .A(_102_), .B(_104_), .C(_97_), .Y(_105_) );
OAI21X1 OAI21X1_68 ( .A(_99_), .B(_100_), .C(_105_), .Y(w_C_20_) );
NOR2X1 NOR2X1_77 ( .A(_99_), .B(_100_), .Y(_106_) );
INVX1 INVX1_119 ( .A(_106_), .Y(_107_) );
AND2X2 AND2X2_64 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_108_) );
INVX1 INVX1_120 ( .A(_108_), .Y(_109_) );
NAND3X1 NAND3X1_75 ( .A(_107_), .B(_109_), .C(_105_), .Y(_110_) );
OAI21X1 OAI21X1_69 ( .A(i_add2[20]), .B(i_add1[20]), .C(_110_), .Y(_111_) );
INVX1 INVX1_121 ( .A(_111_), .Y(w_C_21_) );
INVX1 INVX1_122 ( .A(i_add2[21]), .Y(_112_) );
INVX1 INVX1_123 ( .A(i_add1[21]), .Y(_113_) );
NOR2X1 NOR2X1_78 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_114_) );
INVX1 INVX1_124 ( .A(_114_), .Y(_115_) );
NOR2X1 NOR2X1_79 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_116_) );
INVX1 INVX1_125 ( .A(_116_), .Y(_117_) );
NAND3X1 NAND3X1_76 ( .A(_115_), .B(_117_), .C(_110_), .Y(_118_) );
OAI21X1 OAI21X1_70 ( .A(_112_), .B(_113_), .C(_118_), .Y(w_C_22_) );
NOR2X1 NOR2X1_80 ( .A(_112_), .B(_113_), .Y(_119_) );
INVX1 INVX1_126 ( .A(_119_), .Y(_120_) );
AND2X2 AND2X2_65 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_121_) );
INVX1 INVX1_127 ( .A(_121_), .Y(_122_) );
NAND3X1 NAND3X1_77 ( .A(_120_), .B(_122_), .C(_118_), .Y(_123_) );
OAI21X1 OAI21X1_71 ( .A(i_add2[22]), .B(i_add1[22]), .C(_123_), .Y(_124_) );
INVX1 INVX1_128 ( .A(_124_), .Y(w_C_23_) );
INVX1 INVX1_129 ( .A(i_add2[23]), .Y(_125_) );
INVX1 INVX1_130 ( .A(i_add1[23]), .Y(_126_) );
NOR2X1 NOR2X1_81 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_127_) );
INVX1 INVX1_131 ( .A(_127_), .Y(_128_) );
NOR2X1 NOR2X1_82 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_129_) );
INVX1 INVX1_132 ( .A(_129_), .Y(_130_) );
NAND3X1 NAND3X1_78 ( .A(_128_), .B(_130_), .C(_123_), .Y(_131_) );
OAI21X1 OAI21X1_72 ( .A(_125_), .B(_126_), .C(_131_), .Y(w_C_24_) );
NOR2X1 NOR2X1_83 ( .A(_125_), .B(_126_), .Y(_132_) );
INVX1 INVX1_133 ( .A(_132_), .Y(_133_) );
AND2X2 AND2X2_66 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_134_) );
INVX1 INVX1_134 ( .A(_134_), .Y(_135_) );
NAND3X1 NAND3X1_79 ( .A(_133_), .B(_135_), .C(_131_), .Y(_136_) );
OAI21X1 OAI21X1_73 ( .A(i_add2[24]), .B(i_add1[24]), .C(_136_), .Y(_137_) );
INVX1 INVX1_135 ( .A(_137_), .Y(w_C_25_) );
INVX1 INVX1_136 ( .A(i_add2[25]), .Y(_138_) );
INVX1 INVX1_137 ( .A(i_add1[25]), .Y(_139_) );
NOR2X1 NOR2X1_84 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_140_) );
INVX1 INVX1_138 ( .A(_140_), .Y(_141_) );
NOR2X1 NOR2X1_85 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_142_) );
INVX1 INVX1_139 ( .A(_142_), .Y(_143_) );
NAND3X1 NAND3X1_80 ( .A(_141_), .B(_143_), .C(_136_), .Y(_144_) );
OAI21X1 OAI21X1_74 ( .A(_138_), .B(_139_), .C(_144_), .Y(w_C_26_) );
NOR2X1 NOR2X1_86 ( .A(_138_), .B(_139_), .Y(_145_) );
INVX1 INVX1_140 ( .A(_145_), .Y(_146_) );
AND2X2 AND2X2_67 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_147_) );
INVX1 INVX1_141 ( .A(_147_), .Y(_148_) );
NAND3X1 NAND3X1_81 ( .A(_146_), .B(_148_), .C(_144_), .Y(_149_) );
OAI21X1 OAI21X1_75 ( .A(i_add2[26]), .B(i_add1[26]), .C(_149_), .Y(_150_) );
INVX1 INVX1_142 ( .A(_150_), .Y(w_C_27_) );
INVX1 INVX1_143 ( .A(i_add2[27]), .Y(_151_) );
INVX1 INVX1_144 ( .A(i_add1[27]), .Y(_152_) );
NOR2X1 NOR2X1_87 ( .A(i_add2[26]), .B(i_add1[26]), .Y(_153_) );
INVX1 INVX1_145 ( .A(_153_), .Y(_154_) );
NOR2X1 NOR2X1_88 ( .A(i_add2[27]), .B(i_add1[27]), .Y(_155_) );
INVX1 INVX1_146 ( .A(_155_), .Y(_156_) );
NAND3X1 NAND3X1_82 ( .A(_154_), .B(_156_), .C(_149_), .Y(_157_) );
OAI21X1 OAI21X1_76 ( .A(_151_), .B(_152_), .C(_157_), .Y(w_C_28_) );
NOR2X1 NOR2X1_89 ( .A(_151_), .B(_152_), .Y(_158_) );
INVX1 INVX1_147 ( .A(_158_), .Y(_159_) );
AND2X2 AND2X2_68 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_160_) );
INVX1 INVX1_148 ( .A(_160_), .Y(_161_) );
NAND3X1 NAND3X1_83 ( .A(_159_), .B(_161_), .C(_157_), .Y(_162_) );
OAI21X1 OAI21X1_77 ( .A(i_add2[28]), .B(i_add1[28]), .C(_162_), .Y(_163_) );
INVX1 INVX1_149 ( .A(_163_), .Y(w_C_29_) );
INVX1 INVX1_150 ( .A(i_add2[29]), .Y(_164_) );
INVX1 INVX1_151 ( .A(i_add1[29]), .Y(_165_) );
NOR2X1 NOR2X1_90 ( .A(i_add2[28]), .B(i_add1[28]), .Y(_166_) );
INVX1 INVX1_152 ( .A(_166_), .Y(_167_) );
NOR2X1 NOR2X1_91 ( .A(i_add2[29]), .B(i_add1[29]), .Y(_168_) );
INVX1 INVX1_153 ( .A(_168_), .Y(_169_) );
NAND3X1 NAND3X1_84 ( .A(_167_), .B(_169_), .C(_162_), .Y(_170_) );
OAI21X1 OAI21X1_78 ( .A(_164_), .B(_165_), .C(_170_), .Y(w_C_30_) );
NOR2X1 NOR2X1_92 ( .A(_164_), .B(_165_), .Y(_171_) );
INVX1 INVX1_154 ( .A(_171_), .Y(_172_) );
AND2X2 AND2X2_69 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_173_) );
INVX1 INVX1_155 ( .A(_173_), .Y(_174_) );
NAND3X1 NAND3X1_85 ( .A(_172_), .B(_174_), .C(_170_), .Y(_175_) );
OAI21X1 OAI21X1_79 ( .A(i_add2[30]), .B(i_add1[30]), .C(_175_), .Y(_176_) );
INVX1 INVX1_156 ( .A(_176_), .Y(w_C_31_) );
INVX1 INVX1_157 ( .A(i_add2[31]), .Y(_177_) );
INVX1 INVX1_158 ( .A(i_add1[31]), .Y(_178_) );
NOR2X1 NOR2X1_93 ( .A(i_add2[30]), .B(i_add1[30]), .Y(_179_) );
INVX1 INVX1_159 ( .A(_179_), .Y(_180_) );
NOR2X1 NOR2X1_94 ( .A(i_add2[31]), .B(i_add1[31]), .Y(_181_) );
INVX1 INVX1_160 ( .A(_181_), .Y(_182_) );
NAND3X1 NAND3X1_86 ( .A(_180_), .B(_182_), .C(_175_), .Y(_183_) );
OAI21X1 OAI21X1_80 ( .A(_177_), .B(_178_), .C(_183_), .Y(w_C_32_) );
NOR2X1 NOR2X1_95 ( .A(_177_), .B(_178_), .Y(_184_) );
INVX1 INVX1_161 ( .A(_184_), .Y(_185_) );
AND2X2 AND2X2_70 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_186_) );
INVX1 INVX1_162 ( .A(_186_), .Y(_187_) );
NAND3X1 NAND3X1_87 ( .A(_185_), .B(_187_), .C(_183_), .Y(_188_) );
OAI21X1 OAI21X1_81 ( .A(i_add2[32]), .B(i_add1[32]), .C(_188_), .Y(_189_) );
INVX1 INVX1_163 ( .A(_189_), .Y(w_C_33_) );
INVX1 INVX1_164 ( .A(i_add2[33]), .Y(_190_) );
INVX1 INVX1_165 ( .A(i_add1[33]), .Y(_191_) );
NOR2X1 NOR2X1_96 ( .A(i_add2[32]), .B(i_add1[32]), .Y(_192_) );
INVX1 INVX1_166 ( .A(_192_), .Y(_193_) );
NOR2X1 NOR2X1_97 ( .A(i_add2[33]), .B(i_add1[33]), .Y(_194_) );
INVX1 INVX1_167 ( .A(_194_), .Y(_195_) );
NAND3X1 NAND3X1_88 ( .A(_193_), .B(_195_), .C(_188_), .Y(_196_) );
OAI21X1 OAI21X1_82 ( .A(_190_), .B(_191_), .C(_196_), .Y(w_C_34_) );
NOR2X1 NOR2X1_98 ( .A(_190_), .B(_191_), .Y(_197_) );
INVX1 INVX1_168 ( .A(_197_), .Y(_198_) );
AND2X2 AND2X2_71 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_199_) );
INVX1 INVX1_169 ( .A(_199_), .Y(_200_) );
NAND3X1 NAND3X1_89 ( .A(_198_), .B(_200_), .C(_196_), .Y(_201_) );
OAI21X1 OAI21X1_83 ( .A(i_add2[34]), .B(i_add1[34]), .C(_201_), .Y(_202_) );
INVX1 INVX1_170 ( .A(_202_), .Y(w_C_35_) );
INVX1 INVX1_171 ( .A(i_add2[35]), .Y(_203_) );
INVX1 INVX1_172 ( .A(i_add1[35]), .Y(_204_) );
NOR2X1 NOR2X1_99 ( .A(i_add2[34]), .B(i_add1[34]), .Y(_205_) );
INVX1 INVX1_173 ( .A(_205_), .Y(_206_) );
NOR2X1 NOR2X1_100 ( .A(i_add2[35]), .B(i_add1[35]), .Y(_207_) );
INVX1 INVX1_174 ( .A(_207_), .Y(_208_) );
NAND3X1 NAND3X1_90 ( .A(_206_), .B(_208_), .C(_201_), .Y(_209_) );
OAI21X1 OAI21X1_84 ( .A(_203_), .B(_204_), .C(_209_), .Y(w_C_36_) );
NOR2X1 NOR2X1_101 ( .A(_203_), .B(_204_), .Y(_210_) );
INVX1 INVX1_175 ( .A(_210_), .Y(_211_) );
AND2X2 AND2X2_72 ( .A(i_add2[36]), .B(i_add1[36]), .Y(_212_) );
INVX1 INVX1_176 ( .A(_212_), .Y(_213_) );
NAND3X1 NAND3X1_91 ( .A(_211_), .B(_213_), .C(_209_), .Y(_214_) );
OAI21X1 OAI21X1_85 ( .A(i_add2[36]), .B(i_add1[36]), .C(_214_), .Y(_215_) );
BUFX2 BUFX2_1 ( .A(_274__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_274__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_274__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_274__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_274__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_274__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_274__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_274__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_274__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_274__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_274__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_274__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_274__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_274__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_274__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_274__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_274__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_274__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_274__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_274__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_274__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_274__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_274__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_274__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_274__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_274__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(_274__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .A(_274__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .A(_274__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .A(_274__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .A(_274__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .A(_274__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .A(_274__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .A(_274__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .A(_274__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .A(_274__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .A(_274__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .A(_274__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .A(_274__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .A(_274__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .A(_274__40_), .Y(o_result[40]) );
BUFX2 BUFX2_42 ( .A(_274__41_), .Y(o_result[41]) );
BUFX2 BUFX2_43 ( .A(_274__42_), .Y(o_result[42]) );
BUFX2 BUFX2_44 ( .A(_274__43_), .Y(o_result[43]) );
BUFX2 BUFX2_45 ( .A(_274__44_), .Y(o_result[44]) );
BUFX2 BUFX2_46 ( .A(_274__45_), .Y(o_result[45]) );
BUFX2 BUFX2_47 ( .A(_274__46_), .Y(o_result[46]) );
BUFX2 BUFX2_48 ( .A(_274__47_), .Y(o_result[47]) );
BUFX2 BUFX2_49 ( .A(w_C_48_), .Y(o_result[48]) );
INVX1 INVX1_177 ( .A(w_C_4_), .Y(_278_) );
OR2X2 OR2X2_51 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_279_) );
NAND2X1 NAND2X1_113 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_280_) );
NAND3X1 NAND3X1_92 ( .A(_278_), .B(_280_), .C(_279_), .Y(_281_) );
NOR2X1 NOR2X1_102 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_275_) );
AND2X2 AND2X2_73 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_276_) );
OAI21X1 OAI21X1_86 ( .A(_275_), .B(_276_), .C(w_C_4_), .Y(_277_) );
NAND2X1 NAND2X1_114 ( .A(_277_), .B(_281_), .Y(_274__4_) );
INVX1 INVX1_178 ( .A(w_C_5_), .Y(_285_) );
OR2X2 OR2X2_52 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_286_) );
NAND2X1 NAND2X1_115 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_287_) );
NAND3X1 NAND3X1_93 ( .A(_285_), .B(_287_), .C(_286_), .Y(_288_) );
NOR2X1 NOR2X1_103 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_282_) );
AND2X2 AND2X2_74 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_283_) );
OAI21X1 OAI21X1_87 ( .A(_282_), .B(_283_), .C(w_C_5_), .Y(_284_) );
NAND2X1 NAND2X1_116 ( .A(_284_), .B(_288_), .Y(_274__5_) );
INVX1 INVX1_179 ( .A(w_C_6_), .Y(_292_) );
OR2X2 OR2X2_53 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_293_) );
BUFX2 BUFX2_50 ( .A(w_C_48_), .Y(_274__48_) );
BUFX2 BUFX2_51 ( .A(gnd), .Y(w_C_0_) );
endmodule
