* NGSPICE file created from csa_16bit.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

.subckt csa_16bit vdd gnd i_add_term1[0] i_add_term1[1] i_add_term1[2] i_add_term1[3]
+ i_add_term1[4] i_add_term1[5] i_add_term1[6] i_add_term1[7] i_add_term1[8] i_add_term1[9]
+ i_add_term1[10] i_add_term1[11] i_add_term1[12] i_add_term1[13] i_add_term1[14]
+ i_add_term1[15] i_add_term2[0] i_add_term2[1] i_add_term2[2] i_add_term2[3] i_add_term2[4]
+ i_add_term2[5] i_add_term2[6] i_add_term2[7] i_add_term2[8] i_add_term2[9] i_add_term2[10]
+ i_add_term2[11] i_add_term2[12] i_add_term2[13] i_add_term2[14] i_add_term2[15]
+ sum[0] sum[1] sum[2] sum[3] sum[4] sum[5] sum[6] sum[7] sum[8] sum[9] sum[10] sum[11]
+ sum[12] sum[13] sum[14] sum[15] cout
XFILL_0_0_2 gnd vdd FILL
XNOR2X1_26 i_add_term2[3] i_add_term1[3] gnd NOR2X1_26/Y vdd NOR2X1
XFILL_1_1_0 gnd vdd FILL
XOR2X2_11 i_add_term2[9] i_add_term1[9] gnd OR2X2_11/Y vdd OR2X2
XFILL_7_0_2 gnd vdd FILL
XBUFX2_3 BUFX2_3/A gnd sum[1] vdd BUFX2
XOAI21X1_70 NOR2X1_28/Y AND2X2_28/Y INVX1_43/A gnd OAI21X1_70/Y vdd OAI21X1
XOAI21X1_34 INVX1_22/Y NOR2X1_12/Y OAI21X1_34/C gnd INVX1_20/A vdd OAI21X1
XNAND3X1_18 INVX1_33/Y NAND3X1_18/B OR2X2_18/Y gnd NAND2X1_51/B vdd NAND3X1
XNAND2X1_2 NAND2X1_2/A BUFX2_22/A gnd OAI21X1_2/C vdd NAND2X1
XNAND2X1_13 OAI21X1_12/Y NAND3X1_4/Y gnd INVX1_4/A vdd NAND2X1
XNAND2X1_49 OAI21X1_48/Y NAND2X1_49/B gnd INVX1_28/A vdd NAND2X1
XAND2X2_24 i_add_term2[14] i_add_term1[14] gnd AND2X2_24/Y vdd AND2X2
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XNOR2X1_27 i_add_term2[1] i_add_term1[1] gnd NOR2X1_27/Y vdd NOR2X1
XFILL_1_1_1 gnd vdd FILL
XOR2X2_12 i_add_term2[10] i_add_term1[10] gnd OR2X2_12/Y vdd OR2X2
XNAND2X1_14 i_add_term2[4] i_add_term1[4] gnd NAND3X1_5/B vdd NAND2X1
XNAND2X1_50 i_add_term2[15] i_add_term1[15] gnd NAND3X1_18/B vdd NAND2X1
XBUFX2_4 BUFX2_4/A gnd sum[2] vdd BUFX2
XOAI21X1_71 INVX1_43/Y NOR2X1_28/Y OAI21X1_71/C gnd INVX1_41/A vdd OAI21X1
XOAI21X1_35 NOR2X1_13/Y AND2X2_13/Y vdd gnd OAI21X1_35/Y vdd OAI21X1
XAND2X2_25 i_add_term2[0] i_add_term1[0] gnd AND2X2_25/Y vdd AND2X2
XNAND2X1_3 BUFX2_22/A NAND2X1_3/B gnd OAI21X1_3/C vdd NAND2X1
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XNAND3X1_19 INVX1_34/Y NAND2X1_52/Y OR2X2_19/Y gnd NAND3X1_19/Y vdd NAND3X1
XNOR2X1_28 i_add_term2[2] i_add_term1[2] gnd NOR2X1_28/Y vdd NOR2X1
XFILL_1_1_2 gnd vdd FILL
XOR2X2_13 i_add_term2[8] i_add_term1[8] gnd OR2X2_13/Y vdd OR2X2
XNAND2X1_51 NAND2X1_51/A NAND2X1_51/B gnd INVX1_31/A vdd NAND2X1
XNAND2X1_4 BUFX2_22/A NAND2X1_4/B gnd OAI21X1_4/C vdd NAND2X1
XNAND2X1_15 NAND2X1_15/A NAND3X1_5/Y gnd NAND2X1_2/A vdd NAND2X1
XOAI21X1_36 INVX1_23/Y NOR2X1_13/Y OAI21X1_36/C gnd INVX1_25/A vdd OAI21X1
XBUFX2_5 BUFX2_5/A gnd sum[3] vdd BUFX2
XNAND3X1_20 INVX1_35/Y OAI21X1_55/C OR2X2_20/Y gnd NAND3X1_20/Y vdd NAND3X1
XINVX1_40 gnd gnd INVX1_40/Y vdd INVX1
XAND2X2_26 i_add_term2[3] i_add_term1[3] gnd AND2X2_26/Y vdd AND2X2
XOR2X2_14 i_add_term2[11] i_add_term1[11] gnd OR2X2_14/Y vdd OR2X2
XOAI21X1_37 NOR2X1_14/Y AND2X2_14/Y INVX1_24/A gnd OAI21X1_37/Y vdd OAI21X1
XBUFX2_6 BUFX2_6/A gnd sum[4] vdd BUFX2
XFILL_4_0_0 gnd vdd FILL
XNAND2X1_16 i_add_term2[7] i_add_term1[7] gnd NAND3X1_6/B vdd NAND2X1
XNAND2X1_52 i_add_term2[13] i_add_term1[13] gnd NAND2X1_52/Y vdd NAND2X1
XNAND3X1_21 INVX1_36/Y OAI21X1_57/C OR2X2_21/Y gnd NAND3X1_21/Y vdd NAND3X1
XNAND2X1_5 BUFX2_22/A NAND2X1_5/B gnd OAI21X1_5/C vdd NAND2X1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XAND2X2_27 i_add_term2[1] i_add_term1[1] gnd AND2X2_27/Y vdd AND2X2
XOR2X2_15 i_add_term2[9] i_add_term1[9] gnd OR2X2_15/Y vdd OR2X2
XFILL_4_0_1 gnd vdd FILL
XNAND2X1_6 i_add_term2[4] i_add_term1[4] gnd OAI21X1_7/C vdd NAND2X1
XBUFX2_7 BUFX2_7/A gnd sum[5] vdd BUFX2
XOAI21X1_38 INVX1_24/Y NOR2X1_14/Y NAND2X1_37/Y gnd NAND2X1_22/A vdd OAI21X1
XNAND2X1_17 NAND2X1_17/A NAND3X1_6/Y gnd NAND2X1_5/B vdd NAND2X1
XNAND2X1_53 OAI21X1_52/Y NAND3X1_19/Y gnd INVX1_29/A vdd NAND2X1
XNAND3X1_22 INVX1_37/Y NAND2X1_58/Y OR2X2_22/Y gnd NAND3X1_22/Y vdd NAND3X1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XAND2X2_28 i_add_term2[2] i_add_term1[2] gnd AND2X2_28/Y vdd AND2X2
XFILL_4_1 gnd vdd FILL
XNOR2X1_1 i_add_term2[4] i_add_term1[4] gnd NOR2X1_1/Y vdd NOR2X1
XOR2X2_16 i_add_term2[10] i_add_term1[10] gnd OR2X2_16/Y vdd OR2X2
XBUFX2_8 BUFX2_8/A gnd sum[6] vdd BUFX2
XOAI21X1_39 NOR2X1_15/Y AND2X2_15/Y INVX1_25/A gnd NAND2X1_40/A vdd OAI21X1
XFILL_4_0_2 gnd vdd FILL
XNAND2X1_54 i_add_term2[14] i_add_term1[14] gnd OAI21X1_55/C vdd NAND2X1
XNAND2X1_18 i_add_term2[5] i_add_term1[5] gnd NAND3X1_7/B vdd NAND2X1
XNAND2X1_7 NAND2X1_7/A NAND2X1_7/B gnd INVX1_2/A vdd NAND2X1
XFILL_5_1_0 gnd vdd FILL
XNAND3X1_23 INVX1_38/Y OAI21X1_61/C OR2X2_23/Y gnd NAND3X1_23/Y vdd NAND3X1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XFILL_4_2 gnd vdd FILL
XOR2X2_17 i_add_term2[12] i_add_term1[12] gnd OR2X2_17/Y vdd OR2X2
XNAND2X1_19 NAND2X1_19/A NAND3X1_7/Y gnd NAND2X1_3/B vdd NAND2X1
XOAI21X1_40 INVX1_25/Y NOR2X1_15/Y OAI21X1_40/C gnd INVX1_26/A vdd OAI21X1
XBUFX2_9 BUFX2_9/A gnd sum[7] vdd BUFX2
XFILL_5_1_1 gnd vdd FILL
XNAND2X1_55 OAI21X1_54/Y NAND3X1_20/Y gnd INVX1_30/A vdd NAND2X1
XNOR2X1_2 i_add_term2[7] i_add_term1[7] gnd NOR2X1_2/Y vdd NOR2X1
XNAND3X1_24 INVX1_39/Y OAI21X1_63/C OR2X2_24/Y gnd NAND3X1_24/Y vdd NAND3X1
XNAND2X1_8 i_add_term2[7] i_add_term1[7] gnd NAND2X1_8/Y vdd NAND2X1
XOR2X2_1 i_add_term2[4] i_add_term1[4] gnd OR2X2_1/Y vdd OR2X2
XOR2X2_18 i_add_term2[15] i_add_term1[15] gnd OR2X2_18/Y vdd OR2X2
XOAI21X1_41 NOR2X1_16/Y AND2X2_16/Y INVX1_26/A gnd NAND2X1_42/A vdd OAI21X1
XNAND2X1_56 i_add_term2[12] i_add_term1[12] gnd OAI21X1_57/C vdd NAND2X1
XNOR2X1_3 i_add_term2[5] i_add_term1[5] gnd NOR2X1_3/Y vdd NOR2X1
XNAND3X1_25 INVX1_40/Y NAND2X1_64/Y OR2X2_25/Y gnd NAND2X1_65/B vdd NAND3X1
XNAND2X1_20 i_add_term2[6] i_add_term1[6] gnd NAND3X1_8/B vdd NAND2X1
XFILL_5_1_2 gnd vdd FILL
XNAND2X1_9 OAI21X1_8/Y NAND2X1_9/B gnd INVX1_5/A vdd NAND2X1
XOR2X2_2 i_add_term2[7] i_add_term1[7] gnd OR2X2_2/Y vdd OR2X2
XFILL_1_0_0 gnd vdd FILL
XOAI21X1_42 INVX1_26/Y NOR2X1_16/Y OAI21X1_42/C gnd INVX1_24/A vdd OAI21X1
XNAND2X1_21 OAI21X1_20/Y NAND3X1_8/Y gnd NAND2X1_4/B vdd NAND2X1
XNOR2X1_4 i_add_term2[6] i_add_term1[6] gnd NOR2X1_4/Y vdd NOR2X1
XNAND2X1_57 OAI21X1_56/Y NAND3X1_21/Y gnd NAND2X1_57/Y vdd NAND2X1
XOR2X2_19 i_add_term2[13] i_add_term1[13] gnd OR2X2_19/Y vdd OR2X2
XFILL_8_1 gnd vdd FILL
XINVX1_10 vdd gnd INVX1_10/Y vdd INVX1
XNAND3X1_26 INVX1_41/Y NAND3X1_26/B OR2X2_26/Y gnd NAND2X1_67/B vdd NAND3X1
XOR2X2_3 i_add_term2[5] i_add_term1[5] gnd OR2X2_3/Y vdd OR2X2
XFILL_1_0_1 gnd vdd FILL
XOR2X2_20 i_add_term2[14] i_add_term1[14] gnd OR2X2_20/Y vdd OR2X2
XNAND2X1_22 NAND2X1_22/A OAI21X1_1/Y gnd OAI21X1_22/C vdd NAND2X1
XOAI21X1_43 OAI21X1_47/A INVX1_27/Y OAI21X1_43/C gnd BUFX2_1/A vdd OAI21X1
XNOR2X1_5 i_add_term2[4] i_add_term1[4] gnd NOR2X1_5/Y vdd NOR2X1
XNAND2X1_58 i_add_term2[15] i_add_term1[15] gnd NAND2X1_58/Y vdd NAND2X1
XNAND3X1_27 INVX1_42/Y OAI21X1_69/C OR2X2_27/Y gnd NAND2X1_69/B vdd NAND3X1
XFILL_8_2 gnd vdd FILL
XNAND3X1_1 INVX1_6/Y OAI21X1_7/C OR2X2_1/Y gnd NAND2X1_7/B vdd NAND3X1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XOR2X2_4 i_add_term2[6] i_add_term1[6] gnd OR2X2_4/Y vdd OR2X2
XFILL_1_0_2 gnd vdd FILL
XFILL_2_1_0 gnd vdd FILL
XNAND2X1_59 NAND2X1_59/A NAND3X1_22/Y gnd NAND2X1_47/B vdd NAND2X1
XOR2X2_21 i_add_term2[12] i_add_term1[12] gnd OR2X2_21/Y vdd OR2X2
XNOR2X1_6 i_add_term2[7] i_add_term1[7] gnd NOR2X1_6/Y vdd NOR2X1
XOAI21X1_44 OAI21X1_47/A INVX1_28/Y NAND2X1_44/Y gnd BUFX2_14/A vdd OAI21X1
XNAND2X1_23 NAND2X1_36/Y OAI21X1_1/Y gnd NAND2X1_23/Y vdd NAND2X1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XNAND3X1_28 INVX1_43/Y OAI21X1_71/C OR2X2_28/Y gnd NAND3X1_28/Y vdd NAND3X1
XOR2X2_5 i_add_term2[4] i_add_term1[4] gnd OR2X2_5/Y vdd OR2X2
XNAND3X1_2 INVX1_7/Y NAND2X1_8/Y OR2X2_2/Y gnd NAND2X1_9/B vdd NAND3X1
XOR2X2_22 i_add_term2[15] i_add_term1[15] gnd OR2X2_22/Y vdd OR2X2
XNOR2X1_7 i_add_term2[5] i_add_term1[5] gnd NOR2X1_7/Y vdd NOR2X1
XFILL_2_1_1 gnd vdd FILL
XNAND2X1_24 OAI21X1_1/Y NAND2X1_40/Y gnd NAND2X1_24/Y vdd NAND2X1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XNAND2X1_60 i_add_term2[13] i_add_term1[13] gnd OAI21X1_61/C vdd NAND2X1
XOAI21X1_45 OAI21X1_47/A INVX1_29/Y NAND2X1_45/Y gnd BUFX2_15/A vdd OAI21X1
XNAND3X1_3 INVX1_8/Y NAND3X1_3/B OR2X2_3/Y gnd NAND3X1_3/Y vdd NAND3X1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XOR2X2_6 i_add_term2[7] i_add_term1[7] gnd OR2X2_6/Y vdd OR2X2
XOAI21X1_10 NOR2X1_3/Y AND2X2_3/Y INVX1_8/A gnd NAND2X1_11/A vdd OAI21X1
XNAND2X1_25 OAI21X1_1/Y NAND2X1_25/B gnd OAI21X1_25/C vdd NAND2X1
XNOR2X1_8 i_add_term2[6] i_add_term1[6] gnd NOR2X1_8/Y vdd NOR2X1
XNAND2X1_61 OAI21X1_60/Y NAND3X1_23/Y gnd NAND2X1_61/Y vdd NAND2X1
XOR2X2_23 i_add_term2[13] i_add_term1[13] gnd OR2X2_23/Y vdd OR2X2
XOAI21X1_46 OAI21X1_47/A INVX1_30/Y NAND2X1_46/Y gnd BUFX2_16/A vdd OAI21X1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XFILL_2_1_2 gnd vdd FILL
XOR2X2_7 i_add_term2[5] i_add_term1[5] gnd OR2X2_7/Y vdd OR2X2
XNAND3X1_4 INVX1_9/Y NAND3X1_4/B OR2X2_4/Y gnd NAND3X1_4/Y vdd NAND3X1
XOR2X2_24 i_add_term2[14] i_add_term1[14] gnd OR2X2_24/Y vdd OR2X2
XOAI21X1_47 OAI21X1_47/A INVX1_31/Y OAI21X1_47/C gnd BUFX2_17/A vdd OAI21X1
XOAI21X1_11 INVX1_8/Y NOR2X1_3/Y NAND3X1_3/B gnd INVX1_9/A vdd OAI21X1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XNAND2X1_26 OAI21X1_1/Y NAND2X1_38/Y gnd OAI21X1_26/C vdd NAND2X1
XFILL_3_1 gnd vdd FILL
XNAND2X1_62 i_add_term2[14] i_add_term1[14] gnd OAI21X1_63/C vdd NAND2X1
XNOR2X1_9 i_add_term2[8] i_add_term1[8] gnd NOR2X1_9/Y vdd NOR2X1
XFILL_5_0_0 gnd vdd FILL
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XNAND3X1_5 INVX1_10/Y NAND3X1_5/B OR2X2_5/Y gnd NAND3X1_5/Y vdd NAND3X1
XOR2X2_8 i_add_term2[6] i_add_term1[6] gnd OR2X2_8/Y vdd OR2X2
XOR2X2_25 i_add_term2[0] i_add_term1[0] gnd OR2X2_25/Y vdd OR2X2
XFILL_3_2 gnd vdd FILL
XOAI21X1_12 NOR2X1_4/Y AND2X2_4/Y INVX1_9/A gnd OAI21X1_12/Y vdd OAI21X1
XNAND2X1_63 OAI21X1_62/Y NAND3X1_24/Y gnd NAND2X1_63/Y vdd NAND2X1
XNAND2X1_27 i_add_term2[8] i_add_term1[8] gnd NAND3X1_9/B vdd NAND2X1
XOAI21X1_48 NOR2X1_17/Y AND2X2_17/Y gnd gnd OAI21X1_48/Y vdd OAI21X1
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XFILL_5_0_1 gnd vdd FILL
XNAND3X1_6 INVX1_11/Y NAND3X1_6/B OR2X2_6/Y gnd NAND3X1_6/Y vdd NAND3X1
XOR2X2_9 i_add_term2[8] i_add_term1[8] gnd OR2X2_9/Y vdd OR2X2
XOR2X2_26 i_add_term2[3] i_add_term1[3] gnd OR2X2_26/Y vdd OR2X2
XNAND2X1_64 i_add_term2[0] i_add_term1[0] gnd NAND2X1_64/Y vdd NAND2X1
XOAI21X1_13 INVX1_9/Y NOR2X1_4/Y NAND3X1_4/B gnd INVX1_7/A vdd OAI21X1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XOAI21X1_49 INVX1_32/Y NOR2X1_17/Y OAI21X1_49/C gnd INVX1_34/A vdd OAI21X1
XNAND2X1_28 OAI21X1_27/Y NAND3X1_9/Y gnd INVX1_15/A vdd NAND2X1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XFILL_5_0_2 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XNAND3X1_7 INVX1_12/Y NAND3X1_7/B OR2X2_7/Y gnd NAND3X1_7/Y vdd NAND3X1
XNAND2X1_65 OAI21X1_64/Y NAND2X1_65/B gnd BUFX2_2/A vdd NAND2X1
XOAI21X1_50 NOR2X1_18/Y AND2X2_18/Y INVX1_33/A gnd NAND2X1_51/A vdd OAI21X1
XOR2X2_27 i_add_term2[1] i_add_term1[1] gnd OR2X2_27/Y vdd OR2X2
XNAND2X1_29 i_add_term2[11] i_add_term1[11] gnd NAND2X1_29/Y vdd NAND2X1
XAND2X2_1 i_add_term2[4] i_add_term1[4] gnd AND2X2_1/Y vdd AND2X2
XINVX1_6 gnd gnd INVX1_6/Y vdd INVX1
XOAI21X1_14 NOR2X1_5/Y AND2X2_5/Y vdd gnd NAND2X1_15/A vdd OAI21X1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XNAND3X1_8 INVX1_13/Y NAND3X1_8/B OR2X2_8/Y gnd NAND3X1_8/Y vdd NAND3X1
XFILL_6_1_1 gnd vdd FILL
XNAND2X1_30 NAND2X1_30/A NAND3X1_10/Y gnd INVX1_18/A vdd NAND2X1
XOAI21X1_51 INVX1_33/Y NOR2X1_18/Y NAND3X1_18/B gnd INVX1_27/A vdd OAI21X1
XOAI21X1_15 INVX1_10/Y NOR2X1_5/Y NAND3X1_5/B gnd INVX1_12/A vdd OAI21X1
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XNAND2X1_66 i_add_term2[3] i_add_term1[3] gnd NAND3X1_26/B vdd NAND2X1
XOR2X2_28 i_add_term2[2] i_add_term1[2] gnd OR2X2_28/Y vdd OR2X2
XAND2X2_2 i_add_term2[7] i_add_term1[7] gnd AND2X2_2/Y vdd AND2X2
XINVX1_19 gnd gnd INVX1_19/Y vdd INVX1
XFILL_6_1_2 gnd vdd FILL
XNAND3X1_9 INVX1_19/Y NAND3X1_9/B OR2X2_9/Y gnd NAND3X1_9/Y vdd NAND3X1
XOAI21X1_52 NOR2X1_19/Y AND2X2_19/Y INVX1_34/A gnd OAI21X1_52/Y vdd OAI21X1
XNAND2X1_67 NAND2X1_67/A NAND2X1_67/B gnd BUFX2_5/A vdd NAND2X1
XAND2X2_3 i_add_term2[5] i_add_term1[5] gnd AND2X2_3/Y vdd AND2X2
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XNAND2X1_31 i_add_term2[9] i_add_term1[9] gnd NAND2X1_31/Y vdd NAND2X1
XOAI21X1_16 NOR2X1_6/Y AND2X2_6/Y INVX1_11/A gnd NAND2X1_17/A vdd OAI21X1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XFILL_2_0_0 gnd vdd FILL
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XNAND2X1_32 NAND2X1_32/A NAND2X1_32/B gnd INVX1_16/A vdd NAND2X1
XOAI21X1_17 INVX1_11/Y NOR2X1_6/Y NAND3X1_6/B gnd NAND2X1_1/A vdd OAI21X1
XOAI21X1_53 INVX1_34/Y NOR2X1_19/Y NAND2X1_52/Y gnd INVX1_35/A vdd OAI21X1
XNAND2X1_68 i_add_term2[1] i_add_term1[1] gnd OAI21X1_69/C vdd NAND2X1
XFILL_2_0_1 gnd vdd FILL
XAND2X2_4 i_add_term2[6] i_add_term1[6] gnd AND2X2_4/Y vdd AND2X2
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XNOR2X1_10 i_add_term2[11] i_add_term1[11] gnd NOR2X1_10/Y vdd NOR2X1
XOAI21X1_18 NOR2X1_7/Y AND2X2_7/Y INVX1_12/A gnd NAND2X1_19/A vdd OAI21X1
XAND2X2_5 i_add_term2[4] i_add_term1[4] gnd AND2X2_5/Y vdd AND2X2
XNAND2X1_33 i_add_term2[10] i_add_term1[10] gnd OAI21X1_34/C vdd NAND2X1
XNAND2X1_69 NAND2X1_69/A NAND2X1_69/B gnd BUFX2_3/A vdd NAND2X1
XOAI21X1_54 NOR2X1_20/Y AND2X2_20/Y INVX1_35/A gnd OAI21X1_54/Y vdd OAI21X1
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XFILL_2_0_2 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XNOR2X1_11 i_add_term2[9] i_add_term1[9] gnd NOR2X1_11/Y vdd NOR2X1
XOAI21X1_19 INVX1_12/Y NOR2X1_7/Y NAND3X1_7/B gnd INVX1_13/A vdd OAI21X1
XNAND2X1_34 NAND2X1_34/A NAND2X1_34/B gnd INVX1_17/A vdd NAND2X1
XNAND2X1_70 i_add_term2[2] i_add_term1[2] gnd OAI21X1_71/C vdd NAND2X1
XOAI21X1_55 INVX1_35/Y NOR2X1_20/Y OAI21X1_55/C gnd INVX1_33/A vdd OAI21X1
XBUFX2_10 BUFX2_10/A gnd sum[8] vdd BUFX2
XFILL_2_1 gnd vdd FILL
XINVX1_23 vdd gnd INVX1_23/Y vdd INVX1
XAND2X2_6 i_add_term2[7] i_add_term1[7] gnd AND2X2_6/Y vdd AND2X2
XNOR2X1_12 i_add_term2[10] i_add_term1[10] gnd NOR2X1_12/Y vdd NOR2X1
XFILL_3_1_1 gnd vdd FILL
XAND2X2_7 i_add_term2[5] i_add_term1[5] gnd AND2X2_7/Y vdd AND2X2
XOAI21X1_20 NOR2X1_8/Y AND2X2_8/Y INVX1_13/A gnd OAI21X1_20/Y vdd OAI21X1
XBUFX2_11 BUFX2_11/A gnd sum[9] vdd BUFX2
XOAI21X1_56 NOR2X1_21/Y AND2X2_21/Y vdd gnd OAI21X1_56/Y vdd OAI21X1
XNAND2X1_35 i_add_term2[8] i_add_term1[8] gnd OAI21X1_36/C vdd NAND2X1
XNAND2X1_71 OAI21X1_70/Y NAND3X1_28/Y gnd BUFX2_4/A vdd NAND2X1
XAND2X2_10 i_add_term2[11] i_add_term1[11] gnd AND2X2_10/Y vdd AND2X2
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XFILL_3_1_2 gnd vdd FILL
XNOR2X1_13 i_add_term2[8] i_add_term1[8] gnd NOR2X1_13/Y vdd NOR2X1
XBUFX2_12 BUFX2_12/A gnd sum[10] vdd BUFX2
XOAI21X1_21 INVX1_13/Y NOR2X1_8/Y NAND3X1_8/B gnd INVX1_11/A vdd OAI21X1
XOAI21X1_57 INVX1_36/Y NOR2X1_21/Y OAI21X1_57/C gnd INVX1_38/A vdd OAI21X1
XNAND2X1_36 OAI21X1_35/Y NAND3X1_13/Y gnd NAND2X1_36/Y vdd NAND2X1
XAND2X2_8 i_add_term2[6] i_add_term1[6] gnd AND2X2_8/Y vdd AND2X2
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XNOR2X1_14 i_add_term2[11] i_add_term1[11] gnd NOR2X1_14/Y vdd NOR2X1
XAND2X2_11 i_add_term2[9] i_add_term1[9] gnd AND2X2_11/Y vdd AND2X2
XFILL_6_0_0 gnd vdd FILL
XBUFX2_13 BUFX2_13/A gnd sum[11] vdd BUFX2
XNAND2X1_37 i_add_term2[11] i_add_term1[11] gnd NAND2X1_37/Y vdd NAND2X1
XOAI21X1_22 OAI21X1_1/Y INVX1_14/Y OAI21X1_22/C gnd OAI21X1_47/A vdd OAI21X1
XAND2X2_9 i_add_term2[8] i_add_term1[8] gnd AND2X2_9/Y vdd AND2X2
XOAI21X1_58 NOR2X1_22/Y AND2X2_22/Y INVX1_37/A gnd NAND2X1_59/A vdd OAI21X1
XAND2X2_12 i_add_term2[10] i_add_term1[10] gnd AND2X2_12/Y vdd AND2X2
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XFILL_6_1 gnd vdd FILL
XNOR2X1_15 i_add_term2[9] i_add_term1[9] gnd NOR2X1_15/Y vdd NOR2X1
XFILL_6_0_1 gnd vdd FILL
XOAI21X1_59 INVX1_37/Y NOR2X1_22/Y NAND2X1_58/Y gnd OAI21X1_59/Y vdd OAI21X1
XBUFX2_14 BUFX2_14/A gnd sum[12] vdd BUFX2
XNAND2X1_38 OAI21X1_37/Y NAND2X1_38/B gnd NAND2X1_38/Y vdd NAND2X1
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XOAI21X1_23 OAI21X1_1/Y INVX1_15/Y NAND2X1_23/Y gnd BUFX2_10/A vdd OAI21X1
XFILL_0_1_0 gnd vdd FILL
XNOR2X1_16 i_add_term2[10] i_add_term1[10] gnd NOR2X1_16/Y vdd NOR2X1
XFILL_6_2 gnd vdd FILL
XFILL_6_0_2 gnd vdd FILL
XAND2X2_13 i_add_term2[8] i_add_term1[8] gnd AND2X2_13/Y vdd AND2X2
XFILL_7_1_0 gnd vdd FILL
XOAI21X1_24 OAI21X1_1/Y INVX1_16/Y NAND2X1_24/Y gnd BUFX2_11/A vdd OAI21X1
XNAND2X1_39 i_add_term2[9] i_add_term1[9] gnd OAI21X1_40/C vdd NAND2X1
XOAI21X1_1 BUFX2_22/A INVX1_1/Y NAND2X1_1/Y gnd OAI21X1_1/Y vdd OAI21X1
XBUFX2_15 BUFX2_15/A gnd sum[13] vdd BUFX2
XOAI21X1_60 NOR2X1_23/Y AND2X2_23/Y INVX1_38/A gnd OAI21X1_60/Y vdd OAI21X1
XAND2X2_14 i_add_term2[11] i_add_term1[11] gnd AND2X2_14/Y vdd AND2X2
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XFILL_0_1_1 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XNOR2X1_17 i_add_term2[12] i_add_term1[12] gnd NOR2X1_17/Y vdd NOR2X1
XOAI21X1_2 BUFX2_22/A INVX1_2/Y OAI21X1_2/C gnd BUFX2_6/A vdd OAI21X1
XOAI21X1_61 INVX1_38/Y NOR2X1_23/Y OAI21X1_61/C gnd INVX1_39/A vdd OAI21X1
XBUFX2_16 BUFX2_16/A gnd sum[14] vdd BUFX2
XOAI21X1_25 OAI21X1_1/Y INVX1_17/Y OAI21X1_25/C gnd BUFX2_12/A vdd OAI21X1
XNAND2X1_40 NAND2X1_40/A NAND2X1_40/B gnd NAND2X1_40/Y vdd NAND2X1
XFILL_0_1_2 gnd vdd FILL
XNOR2X1_18 i_add_term2[15] i_add_term1[15] gnd NOR2X1_18/Y vdd NOR2X1
XAND2X2_15 i_add_term2[9] i_add_term1[9] gnd AND2X2_15/Y vdd AND2X2
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XFILL_7_1_2 gnd vdd FILL
XOAI21X1_26 OAI21X1_1/Y INVX1_18/Y OAI21X1_26/C gnd BUFX2_13/A vdd OAI21X1
XBUFX2_17 BUFX2_17/A gnd sum[15] vdd BUFX2
XOAI21X1_3 BUFX2_22/A INVX1_3/Y OAI21X1_3/C gnd BUFX2_7/A vdd OAI21X1
XNAND2X1_41 i_add_term2[10] i_add_term1[10] gnd OAI21X1_42/C vdd NAND2X1
XOAI21X1_62 NOR2X1_24/Y AND2X2_24/Y INVX1_39/A gnd OAI21X1_62/Y vdd OAI21X1
XNAND3X1_10 INVX1_20/Y NAND2X1_29/Y OR2X2_10/Y gnd NAND3X1_10/Y vdd NAND3X1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XAND2X2_16 i_add_term2[10] i_add_term1[10] gnd AND2X2_16/Y vdd AND2X2
XFILL_3_0_0 gnd vdd FILL
XNOR2X1_19 i_add_term2[13] i_add_term1[13] gnd NOR2X1_19/Y vdd NOR2X1
XBUFX2_18 BUFX2_2/A gnd BUFX2_18/Y vdd BUFX2
XOAI21X1_4 BUFX2_22/A INVX1_4/Y OAI21X1_4/C gnd BUFX2_8/A vdd OAI21X1
XNAND2X1_42 NAND2X1_42/A NAND2X1_42/B gnd NAND2X1_25/B vdd NAND2X1
XOAI21X1_63 INVX1_39/Y NOR2X1_24/Y OAI21X1_63/C gnd INVX1_37/A vdd OAI21X1
XOAI21X1_27 NOR2X1_9/Y AND2X2_9/Y gnd gnd OAI21X1_27/Y vdd OAI21X1
XFILL_1_1 gnd vdd FILL
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XNAND3X1_11 INVX1_21/Y NAND2X1_31/Y OR2X2_11/Y gnd NAND2X1_32/B vdd NAND3X1
XAND2X2_17 i_add_term2[12] i_add_term1[12] gnd AND2X2_17/Y vdd AND2X2
XFILL_3_0_1 gnd vdd FILL
XNOR2X1_20 i_add_term2[14] i_add_term1[14] gnd NOR2X1_20/Y vdd NOR2X1
XOAI21X1_64 NOR2X1_25/Y AND2X2_25/Y gnd gnd OAI21X1_64/Y vdd OAI21X1
XNAND2X1_43 OAI21X1_59/Y OAI21X1_47/A gnd OAI21X1_43/C vdd NAND2X1
XOAI21X1_5 BUFX2_22/A INVX1_5/Y OAI21X1_5/C gnd BUFX2_9/A vdd OAI21X1
XOAI21X1_28 INVX1_19/Y NOR2X1_9/Y NAND3X1_9/B gnd INVX1_21/A vdd OAI21X1
XBUFX2_19 BUFX2_3/A gnd BUFX2_19/Y vdd BUFX2
XNAND3X1_12 INVX1_22/Y OAI21X1_34/C OR2X2_12/Y gnd NAND2X1_34/B vdd NAND3X1
XINVX1_32 gnd gnd INVX1_32/Y vdd INVX1
XAND2X2_18 i_add_term2[15] i_add_term1[15] gnd AND2X2_18/Y vdd AND2X2
XFILL_3_0_2 gnd vdd FILL
XNOR2X1_21 i_add_term2[12] i_add_term1[12] gnd NOR2X1_21/Y vdd NOR2X1
XOAI21X1_6 NOR2X1_1/Y AND2X2_1/Y gnd gnd NAND2X1_7/A vdd OAI21X1
XFILL_4_1_0 gnd vdd FILL
XOAI21X1_29 NOR2X1_10/Y AND2X2_10/Y INVX1_20/A gnd NAND2X1_30/A vdd OAI21X1
XOAI21X1_65 INVX1_40/Y NOR2X1_25/Y NAND2X1_64/Y gnd INVX1_42/A vdd OAI21X1
XNAND2X1_44 NAND2X1_57/Y OAI21X1_47/A gnd NAND2X1_44/Y vdd NAND2X1
XBUFX2_20 BUFX2_4/A gnd BUFX2_20/Y vdd BUFX2
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XNAND3X1_13 INVX1_23/Y OAI21X1_36/C OR2X2_13/Y gnd NAND3X1_13/Y vdd NAND3X1
XAND2X2_19 i_add_term2[13] i_add_term1[13] gnd AND2X2_19/Y vdd AND2X2
XNOR2X1_22 i_add_term2[15] i_add_term1[15] gnd NOR2X1_22/Y vdd NOR2X1
XFILL_4_1_1 gnd vdd FILL
XOAI21X1_30 INVX1_20/Y NOR2X1_10/Y NAND2X1_29/Y gnd INVX1_14/A vdd OAI21X1
XOAI21X1_7 INVX1_6/Y NOR2X1_1/Y OAI21X1_7/C gnd INVX1_8/A vdd OAI21X1
XBUFX2_21 BUFX2_5/A gnd BUFX2_21/Y vdd BUFX2
XOAI21X1_66 NOR2X1_26/Y AND2X2_26/Y INVX1_41/A gnd NAND2X1_67/A vdd OAI21X1
XNAND2X1_45 OAI21X1_47/A NAND2X1_61/Y gnd NAND2X1_45/Y vdd NAND2X1
XNAND3X1_14 INVX1_24/Y NAND2X1_37/Y OR2X2_14/Y gnd NAND2X1_38/B vdd NAND3X1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XFILL_5_1 gnd vdd FILL
XAND2X2_20 i_add_term2[14] i_add_term1[14] gnd AND2X2_20/Y vdd AND2X2
XNOR2X1_23 i_add_term2[13] i_add_term1[13] gnd NOR2X1_23/Y vdd NOR2X1
XFILL_4_1_2 gnd vdd FILL
XOAI21X1_8 NOR2X1_2/Y AND2X2_2/Y INVX1_7/A gnd OAI21X1_8/Y vdd OAI21X1
XNAND2X1_10 i_add_term2[5] i_add_term1[5] gnd NAND3X1_3/B vdd NAND2X1
XBUFX2_22 BUFX2_22/A gnd BUFX2_22/Y vdd BUFX2
XOAI21X1_31 NOR2X1_11/Y AND2X2_11/Y INVX1_21/A gnd NAND2X1_32/A vdd OAI21X1
XNAND2X1_46 OAI21X1_47/A NAND2X1_63/Y gnd NAND2X1_46/Y vdd NAND2X1
XOAI21X1_67 INVX1_41/Y NOR2X1_26/Y NAND3X1_26/B gnd BUFX2_22/A vdd OAI21X1
XNAND3X1_15 INVX1_25/Y OAI21X1_40/C OR2X2_15/Y gnd NAND2X1_40/B vdd NAND3X1
XAND2X2_21 i_add_term2[12] i_add_term1[12] gnd AND2X2_21/Y vdd AND2X2
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XFILL_0_0_0 gnd vdd FILL
XNOR2X1_24 i_add_term2[14] i_add_term1[14] gnd NOR2X1_24/Y vdd NOR2X1
XBUFX2_1 BUFX2_1/A gnd cout vdd BUFX2
XNAND2X1_47 OAI21X1_47/A NAND2X1_47/B gnd OAI21X1_47/C vdd NAND2X1
XOAI21X1_32 INVX1_21/Y NOR2X1_11/Y NAND2X1_31/Y gnd INVX1_22/A vdd OAI21X1
XOAI21X1_9 INVX1_7/Y NOR2X1_2/Y NAND2X1_8/Y gnd INVX1_1/A vdd OAI21X1
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_68 NOR2X1_27/Y AND2X2_27/Y INVX1_42/A gnd NAND2X1_69/A vdd OAI21X1
XNAND2X1_11 NAND2X1_11/A NAND3X1_3/Y gnd INVX1_3/A vdd NAND2X1
XNAND3X1_16 INVX1_26/Y OAI21X1_42/C OR2X2_16/Y gnd NAND2X1_42/B vdd NAND3X1
XINVX1_36 vdd gnd INVX1_36/Y vdd INVX1
XNOR2X1_25 i_add_term2[0] i_add_term1[0] gnd NOR2X1_25/Y vdd NOR2X1
XAND2X2_22 i_add_term2[15] i_add_term1[15] gnd AND2X2_22/Y vdd AND2X2
XFILL_0_0_1 gnd vdd FILL
XOR2X2_10 i_add_term2[11] i_add_term1[11] gnd OR2X2_10/Y vdd OR2X2
XBUFX2_2 BUFX2_2/A gnd sum[0] vdd BUFX2
XOAI21X1_33 NOR2X1_12/Y AND2X2_12/Y INVX1_22/A gnd NAND2X1_34/A vdd OAI21X1
XNAND2X1_12 i_add_term2[6] i_add_term1[6] gnd NAND3X1_4/B vdd NAND2X1
XFILL_7_0_1 gnd vdd FILL
XOAI21X1_69 INVX1_42/Y NOR2X1_27/Y OAI21X1_69/C gnd INVX1_43/A vdd OAI21X1
XNAND2X1_48 i_add_term2[12] i_add_term1[12] gnd OAI21X1_49/C vdd NAND2X1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XNAND2X1_1 NAND2X1_1/A BUFX2_22/A gnd NAND2X1_1/Y vdd NAND2X1
XAND2X2_23 i_add_term2[13] i_add_term1[13] gnd AND2X2_23/Y vdd AND2X2
XNAND3X1_17 INVX1_32/Y OAI21X1_49/C OR2X2_17/Y gnd NAND2X1_49/B vdd NAND3X1
.ends

