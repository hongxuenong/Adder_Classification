module csa_25bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_6_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_w_SUM), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
INVX1 INVX1_1 ( .A(_1_), .Y(_37_) );
NAND2X1 NAND2X1_1 ( .A(_2_), .B(1'b0), .Y(_38_) );
OAI21X1 OAI21X1_1 ( .A(1'b0), .B(_37_), .C(_38_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .A(_3__2_), .Y(_39_) );
NAND2X1 NAND2X1_2 ( .A(_4__2_), .B(1'b0), .Y(_40_) );
OAI21X1 OAI21X1_2 ( .A(1'b0), .B(_39_), .C(_40_), .Y(_0__3_) );
INVX1 INVX1_3 ( .A(_3__3_), .Y(_41_) );
NAND2X1 NAND2X1_3 ( .A(1'b0), .B(_4__3_), .Y(_42_) );
OAI21X1 OAI21X1_3 ( .A(1'b0), .B(_41_), .C(_42_), .Y(_0__4_) );
INVX1 INVX1_4 ( .A(_3__0_), .Y(_43_) );
NAND2X1 NAND2X1_4 ( .A(1'b0), .B(_4__0_), .Y(_44_) );
OAI21X1 OAI21X1_4 ( .A(1'b0), .B(_43_), .C(_44_), .Y(_0__1_) );
INVX1 INVX1_5 ( .A(_3__1_), .Y(_45_) );
NAND2X1 NAND2X1_5 ( .A(1'b0), .B(_4__1_), .Y(_46_) );
OAI21X1 OAI21X1_5 ( .A(1'b0), .B(_45_), .C(_46_), .Y(_0__2_) );
INVX1 INVX1_6 ( .A(_7_), .Y(_47_) );
NAND2X1 NAND2X1_6 ( .A(_8_), .B(w_cout_1_), .Y(_48_) );
OAI21X1 OAI21X1_6 ( .A(w_cout_1_), .B(_47_), .C(_48_), .Y(w_cout_2_) );
INVX1 INVX1_7 ( .A(_9__2_), .Y(_49_) );
NAND2X1 NAND2X1_7 ( .A(_10__2_), .B(w_cout_1_), .Y(_50_) );
OAI21X1 OAI21X1_7 ( .A(w_cout_1_), .B(_49_), .C(_50_), .Y(_0__7_) );
INVX1 INVX1_8 ( .A(_9__3_), .Y(_51_) );
NAND2X1 NAND2X1_8 ( .A(w_cout_1_), .B(_10__3_), .Y(_52_) );
OAI21X1 OAI21X1_8 ( .A(w_cout_1_), .B(_51_), .C(_52_), .Y(_0__8_) );
INVX1 INVX1_9 ( .A(_9__0_), .Y(_53_) );
NAND2X1 NAND2X1_9 ( .A(w_cout_1_), .B(_10__0_), .Y(_54_) );
OAI21X1 OAI21X1_9 ( .A(w_cout_1_), .B(_53_), .C(_54_), .Y(_0__5_) );
INVX1 INVX1_10 ( .A(_9__1_), .Y(_55_) );
NAND2X1 NAND2X1_10 ( .A(w_cout_1_), .B(_10__1_), .Y(_56_) );
OAI21X1 OAI21X1_10 ( .A(w_cout_1_), .B(_55_), .C(_56_), .Y(_0__6_) );
INVX1 INVX1_11 ( .A(_13_), .Y(_57_) );
NAND2X1 NAND2X1_11 ( .A(_14_), .B(w_cout_2_), .Y(_58_) );
OAI21X1 OAI21X1_11 ( .A(w_cout_2_), .B(_57_), .C(_58_), .Y(w_cout_3_) );
INVX1 INVX1_12 ( .A(_15__2_), .Y(_59_) );
NAND2X1 NAND2X1_12 ( .A(_16__2_), .B(w_cout_2_), .Y(_60_) );
OAI21X1 OAI21X1_12 ( .A(w_cout_2_), .B(_59_), .C(_60_), .Y(_0__11_) );
INVX1 INVX1_13 ( .A(_15__3_), .Y(_61_) );
NAND2X1 NAND2X1_13 ( .A(w_cout_2_), .B(_16__3_), .Y(_62_) );
OAI21X1 OAI21X1_13 ( .A(w_cout_2_), .B(_61_), .C(_62_), .Y(_0__12_) );
INVX1 INVX1_14 ( .A(_15__0_), .Y(_63_) );
NAND2X1 NAND2X1_14 ( .A(w_cout_2_), .B(_16__0_), .Y(_64_) );
OAI21X1 OAI21X1_14 ( .A(w_cout_2_), .B(_63_), .C(_64_), .Y(_0__9_) );
INVX1 INVX1_15 ( .A(_15__1_), .Y(_65_) );
NAND2X1 NAND2X1_15 ( .A(w_cout_2_), .B(_16__1_), .Y(_66_) );
OAI21X1 OAI21X1_15 ( .A(w_cout_2_), .B(_65_), .C(_66_), .Y(_0__10_) );
INVX1 INVX1_16 ( .A(_19_), .Y(_67_) );
NAND2X1 NAND2X1_16 ( .A(_20_), .B(w_cout_3_), .Y(_68_) );
OAI21X1 OAI21X1_16 ( .A(w_cout_3_), .B(_67_), .C(_68_), .Y(w_cout_4_) );
INVX1 INVX1_17 ( .A(_21__2_), .Y(_69_) );
NAND2X1 NAND2X1_17 ( .A(_22__2_), .B(w_cout_3_), .Y(_70_) );
OAI21X1 OAI21X1_17 ( .A(w_cout_3_), .B(_69_), .C(_70_), .Y(_0__15_) );
INVX1 INVX1_18 ( .A(_21__3_), .Y(_71_) );
NAND2X1 NAND2X1_18 ( .A(w_cout_3_), .B(_22__3_), .Y(_72_) );
OAI21X1 OAI21X1_18 ( .A(w_cout_3_), .B(_71_), .C(_72_), .Y(_0__16_) );
INVX1 INVX1_19 ( .A(_21__0_), .Y(_73_) );
NAND2X1 NAND2X1_19 ( .A(w_cout_3_), .B(_22__0_), .Y(_74_) );
OAI21X1 OAI21X1_19 ( .A(w_cout_3_), .B(_73_), .C(_74_), .Y(_0__13_) );
INVX1 INVX1_20 ( .A(_21__1_), .Y(_75_) );
NAND2X1 NAND2X1_20 ( .A(w_cout_3_), .B(_22__1_), .Y(_76_) );
OAI21X1 OAI21X1_20 ( .A(w_cout_3_), .B(_75_), .C(_76_), .Y(_0__14_) );
INVX1 INVX1_21 ( .A(_25_), .Y(_77_) );
NAND2X1 NAND2X1_21 ( .A(_26_), .B(w_cout_4_), .Y(_78_) );
OAI21X1 OAI21X1_21 ( .A(w_cout_4_), .B(_77_), .C(_78_), .Y(w_cout_5_) );
INVX1 INVX1_22 ( .A(_27__2_), .Y(_79_) );
NAND2X1 NAND2X1_22 ( .A(_28__2_), .B(w_cout_4_), .Y(_80_) );
OAI21X1 OAI21X1_22 ( .A(w_cout_4_), .B(_79_), .C(_80_), .Y(_0__19_) );
INVX1 INVX1_23 ( .A(_27__3_), .Y(_81_) );
NAND2X1 NAND2X1_23 ( .A(w_cout_4_), .B(_28__3_), .Y(_82_) );
OAI21X1 OAI21X1_23 ( .A(w_cout_4_), .B(_81_), .C(_82_), .Y(_0__20_) );
INVX1 INVX1_24 ( .A(_27__0_), .Y(_83_) );
NAND2X1 NAND2X1_24 ( .A(w_cout_4_), .B(_28__0_), .Y(_84_) );
OAI21X1 OAI21X1_24 ( .A(w_cout_4_), .B(_83_), .C(_84_), .Y(_0__17_) );
INVX1 INVX1_25 ( .A(_27__1_), .Y(_85_) );
NAND2X1 NAND2X1_25 ( .A(w_cout_4_), .B(_28__1_), .Y(_86_) );
OAI21X1 OAI21X1_25 ( .A(w_cout_4_), .B(_85_), .C(_86_), .Y(_0__18_) );
INVX1 INVX1_26 ( .A(_31_), .Y(_87_) );
NAND2X1 NAND2X1_26 ( .A(_32_), .B(w_cout_5_), .Y(_88_) );
OAI21X1 OAI21X1_26 ( .A(w_cout_5_), .B(_87_), .C(_88_), .Y(w_cout_6_) );
INVX1 INVX1_27 ( .A(_33__2_), .Y(_89_) );
NAND2X1 NAND2X1_27 ( .A(_34__2_), .B(w_cout_5_), .Y(_90_) );
OAI21X1 OAI21X1_27 ( .A(w_cout_5_), .B(_89_), .C(_90_), .Y(_0__23_) );
INVX1 INVX1_28 ( .A(_33__3_), .Y(_91_) );
NAND2X1 NAND2X1_28 ( .A(w_cout_5_), .B(_34__3_), .Y(_92_) );
OAI21X1 OAI21X1_28 ( .A(w_cout_5_), .B(_91_), .C(_92_), .Y(_0__24_) );
INVX1 INVX1_29 ( .A(_33__0_), .Y(_93_) );
NAND2X1 NAND2X1_29 ( .A(w_cout_5_), .B(_34__0_), .Y(_94_) );
OAI21X1 OAI21X1_29 ( .A(w_cout_5_), .B(_93_), .C(_94_), .Y(_0__21_) );
INVX1 INVX1_30 ( .A(_33__1_), .Y(_95_) );
NAND2X1 NAND2X1_30 ( .A(w_cout_5_), .B(_34__1_), .Y(_96_) );
OAI21X1 OAI21X1_30 ( .A(w_cout_5_), .B(_95_), .C(_96_), .Y(_0__22_) );
INVX1 INVX1_31 ( .A(1'b0), .Y(_100_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_101_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_102_) );
NAND3X1 NAND3X1_1 ( .A(_100_), .B(_102_), .C(_101_), .Y(_103_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_97_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_98_) );
OAI21X1 OAI21X1_31 ( .A(_97_), .B(_98_), .C(1'b0), .Y(_99_) );
NAND2X1 NAND2X1_32 ( .A(_99_), .B(_103_), .Y(_3__0_) );
OAI21X1 OAI21X1_32 ( .A(_100_), .B(_97_), .C(_102_), .Y(_5__1_) );
INVX1 INVX1_32 ( .A(_5__1_), .Y(_107_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_108_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_109_) );
NAND3X1 NAND3X1_2 ( .A(_107_), .B(_109_), .C(_108_), .Y(_110_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_104_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_105_) );
OAI21X1 OAI21X1_33 ( .A(_104_), .B(_105_), .C(_5__1_), .Y(_106_) );
NAND2X1 NAND2X1_34 ( .A(_106_), .B(_110_), .Y(_3__1_) );
OAI21X1 OAI21X1_34 ( .A(_107_), .B(_104_), .C(_109_), .Y(_5__2_) );
INVX1 INVX1_33 ( .A(_5__2_), .Y(_114_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_115_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_116_) );
NAND3X1 NAND3X1_3 ( .A(_114_), .B(_116_), .C(_115_), .Y(_117_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_111_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_112_) );
OAI21X1 OAI21X1_35 ( .A(_111_), .B(_112_), .C(_5__2_), .Y(_113_) );
NAND2X1 NAND2X1_36 ( .A(_113_), .B(_117_), .Y(_3__2_) );
OAI21X1 OAI21X1_36 ( .A(_114_), .B(_111_), .C(_116_), .Y(_5__3_) );
INVX1 INVX1_34 ( .A(_5__3_), .Y(_121_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_122_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_123_) );
NAND3X1 NAND3X1_4 ( .A(_121_), .B(_123_), .C(_122_), .Y(_124_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_118_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_119_) );
OAI21X1 OAI21X1_37 ( .A(_118_), .B(_119_), .C(_5__3_), .Y(_120_) );
NAND2X1 NAND2X1_38 ( .A(_120_), .B(_124_), .Y(_3__3_) );
OAI21X1 OAI21X1_38 ( .A(_121_), .B(_118_), .C(_123_), .Y(_1_) );
INVX1 INVX1_35 ( .A(1'b1), .Y(_128_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_129_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_130_) );
NAND3X1 NAND3X1_5 ( .A(_128_), .B(_130_), .C(_129_), .Y(_131_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_125_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_126_) );
OAI21X1 OAI21X1_39 ( .A(_125_), .B(_126_), .C(1'b1), .Y(_127_) );
NAND2X1 NAND2X1_40 ( .A(_127_), .B(_131_), .Y(_4__0_) );
OAI21X1 OAI21X1_40 ( .A(_128_), .B(_125_), .C(_130_), .Y(_6__1_) );
INVX1 INVX1_36 ( .A(_6__1_), .Y(_135_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_136_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_137_) );
NAND3X1 NAND3X1_6 ( .A(_135_), .B(_137_), .C(_136_), .Y(_138_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_132_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_133_) );
OAI21X1 OAI21X1_41 ( .A(_132_), .B(_133_), .C(_6__1_), .Y(_134_) );
NAND2X1 NAND2X1_42 ( .A(_134_), .B(_138_), .Y(_4__1_) );
OAI21X1 OAI21X1_42 ( .A(_135_), .B(_132_), .C(_137_), .Y(_6__2_) );
INVX1 INVX1_37 ( .A(_6__2_), .Y(_142_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_143_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_144_) );
NAND3X1 NAND3X1_7 ( .A(_142_), .B(_144_), .C(_143_), .Y(_145_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_139_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_140_) );
OAI21X1 OAI21X1_43 ( .A(_139_), .B(_140_), .C(_6__2_), .Y(_141_) );
NAND2X1 NAND2X1_44 ( .A(_141_), .B(_145_), .Y(_4__2_) );
OAI21X1 OAI21X1_44 ( .A(_142_), .B(_139_), .C(_144_), .Y(_6__3_) );
INVX1 INVX1_38 ( .A(_6__3_), .Y(_149_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_150_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_151_) );
NAND3X1 NAND3X1_8 ( .A(_149_), .B(_151_), .C(_150_), .Y(_152_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_146_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_147_) );
OAI21X1 OAI21X1_45 ( .A(_146_), .B(_147_), .C(_6__3_), .Y(_148_) );
NAND2X1 NAND2X1_46 ( .A(_148_), .B(_152_), .Y(_4__3_) );
OAI21X1 OAI21X1_46 ( .A(_149_), .B(_146_), .C(_151_), .Y(_2_) );
INVX1 INVX1_39 ( .A(1'b0), .Y(_156_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_157_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_158_) );
NAND3X1 NAND3X1_9 ( .A(_156_), .B(_158_), .C(_157_), .Y(_159_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_153_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_154_) );
OAI21X1 OAI21X1_47 ( .A(_153_), .B(_154_), .C(1'b0), .Y(_155_) );
NAND2X1 NAND2X1_48 ( .A(_155_), .B(_159_), .Y(_9__0_) );
OAI21X1 OAI21X1_48 ( .A(_156_), .B(_153_), .C(_158_), .Y(_11__1_) );
INVX1 INVX1_40 ( .A(_11__1_), .Y(_163_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_164_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_165_) );
NAND3X1 NAND3X1_10 ( .A(_163_), .B(_165_), .C(_164_), .Y(_166_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_160_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_161_) );
OAI21X1 OAI21X1_49 ( .A(_160_), .B(_161_), .C(_11__1_), .Y(_162_) );
NAND2X1 NAND2X1_50 ( .A(_162_), .B(_166_), .Y(_9__1_) );
OAI21X1 OAI21X1_50 ( .A(_163_), .B(_160_), .C(_165_), .Y(_11__2_) );
INVX1 INVX1_41 ( .A(_11__2_), .Y(_170_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_171_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_172_) );
NAND3X1 NAND3X1_11 ( .A(_170_), .B(_172_), .C(_171_), .Y(_173_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_167_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_168_) );
OAI21X1 OAI21X1_51 ( .A(_167_), .B(_168_), .C(_11__2_), .Y(_169_) );
NAND2X1 NAND2X1_52 ( .A(_169_), .B(_173_), .Y(_9__2_) );
OAI21X1 OAI21X1_52 ( .A(_170_), .B(_167_), .C(_172_), .Y(_11__3_) );
INVX1 INVX1_42 ( .A(_11__3_), .Y(_177_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_178_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_179_) );
NAND3X1 NAND3X1_12 ( .A(_177_), .B(_179_), .C(_178_), .Y(_180_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_174_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_175_) );
OAI21X1 OAI21X1_53 ( .A(_174_), .B(_175_), .C(_11__3_), .Y(_176_) );
NAND2X1 NAND2X1_54 ( .A(_176_), .B(_180_), .Y(_9__3_) );
OAI21X1 OAI21X1_54 ( .A(_177_), .B(_174_), .C(_179_), .Y(_7_) );
INVX1 INVX1_43 ( .A(1'b1), .Y(_184_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_185_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_186_) );
NAND3X1 NAND3X1_13 ( .A(_184_), .B(_186_), .C(_185_), .Y(_187_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_181_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_182_) );
OAI21X1 OAI21X1_55 ( .A(_181_), .B(_182_), .C(1'b1), .Y(_183_) );
NAND2X1 NAND2X1_56 ( .A(_183_), .B(_187_), .Y(_10__0_) );
OAI21X1 OAI21X1_56 ( .A(_184_), .B(_181_), .C(_186_), .Y(_12__1_) );
INVX1 INVX1_44 ( .A(_12__1_), .Y(_191_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_192_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_193_) );
NAND3X1 NAND3X1_14 ( .A(_191_), .B(_193_), .C(_192_), .Y(_194_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_188_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_189_) );
OAI21X1 OAI21X1_57 ( .A(_188_), .B(_189_), .C(_12__1_), .Y(_190_) );
NAND2X1 NAND2X1_58 ( .A(_190_), .B(_194_), .Y(_10__1_) );
OAI21X1 OAI21X1_58 ( .A(_191_), .B(_188_), .C(_193_), .Y(_12__2_) );
INVX1 INVX1_45 ( .A(_12__2_), .Y(_198_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_199_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_200_) );
NAND3X1 NAND3X1_15 ( .A(_198_), .B(_200_), .C(_199_), .Y(_201_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_195_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_196_) );
OAI21X1 OAI21X1_59 ( .A(_195_), .B(_196_), .C(_12__2_), .Y(_197_) );
NAND2X1 NAND2X1_60 ( .A(_197_), .B(_201_), .Y(_10__2_) );
OAI21X1 OAI21X1_60 ( .A(_198_), .B(_195_), .C(_200_), .Y(_12__3_) );
INVX1 INVX1_46 ( .A(_12__3_), .Y(_205_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_206_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_207_) );
NAND3X1 NAND3X1_16 ( .A(_205_), .B(_207_), .C(_206_), .Y(_208_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_202_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_203_) );
OAI21X1 OAI21X1_61 ( .A(_202_), .B(_203_), .C(_12__3_), .Y(_204_) );
NAND2X1 NAND2X1_62 ( .A(_204_), .B(_208_), .Y(_10__3_) );
OAI21X1 OAI21X1_62 ( .A(_205_), .B(_202_), .C(_207_), .Y(_8_) );
INVX1 INVX1_47 ( .A(1'b0), .Y(_212_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_213_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_214_) );
NAND3X1 NAND3X1_17 ( .A(_212_), .B(_214_), .C(_213_), .Y(_215_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_209_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_210_) );
OAI21X1 OAI21X1_63 ( .A(_209_), .B(_210_), .C(1'b0), .Y(_211_) );
NAND2X1 NAND2X1_64 ( .A(_211_), .B(_215_), .Y(_15__0_) );
OAI21X1 OAI21X1_64 ( .A(_212_), .B(_209_), .C(_214_), .Y(_17__1_) );
INVX1 INVX1_48 ( .A(_17__1_), .Y(_219_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_220_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_221_) );
NAND3X1 NAND3X1_18 ( .A(_219_), .B(_221_), .C(_220_), .Y(_222_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_216_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_217_) );
OAI21X1 OAI21X1_65 ( .A(_216_), .B(_217_), .C(_17__1_), .Y(_218_) );
NAND2X1 NAND2X1_66 ( .A(_218_), .B(_222_), .Y(_15__1_) );
OAI21X1 OAI21X1_66 ( .A(_219_), .B(_216_), .C(_221_), .Y(_17__2_) );
INVX1 INVX1_49 ( .A(_17__2_), .Y(_226_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_227_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_228_) );
NAND3X1 NAND3X1_19 ( .A(_226_), .B(_228_), .C(_227_), .Y(_229_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_223_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_224_) );
OAI21X1 OAI21X1_67 ( .A(_223_), .B(_224_), .C(_17__2_), .Y(_225_) );
NAND2X1 NAND2X1_68 ( .A(_225_), .B(_229_), .Y(_15__2_) );
OAI21X1 OAI21X1_68 ( .A(_226_), .B(_223_), .C(_228_), .Y(_17__3_) );
INVX1 INVX1_50 ( .A(_17__3_), .Y(_233_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_234_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_235_) );
NAND3X1 NAND3X1_20 ( .A(_233_), .B(_235_), .C(_234_), .Y(_236_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_230_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_231_) );
OAI21X1 OAI21X1_69 ( .A(_230_), .B(_231_), .C(_17__3_), .Y(_232_) );
NAND2X1 NAND2X1_70 ( .A(_232_), .B(_236_), .Y(_15__3_) );
OAI21X1 OAI21X1_70 ( .A(_233_), .B(_230_), .C(_235_), .Y(_13_) );
INVX1 INVX1_51 ( .A(1'b1), .Y(_240_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_241_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_242_) );
NAND3X1 NAND3X1_21 ( .A(_240_), .B(_242_), .C(_241_), .Y(_243_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_237_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_238_) );
OAI21X1 OAI21X1_71 ( .A(_237_), .B(_238_), .C(1'b1), .Y(_239_) );
NAND2X1 NAND2X1_72 ( .A(_239_), .B(_243_), .Y(_16__0_) );
OAI21X1 OAI21X1_72 ( .A(_240_), .B(_237_), .C(_242_), .Y(_18__1_) );
INVX1 INVX1_52 ( .A(_18__1_), .Y(_247_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_248_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_249_) );
NAND3X1 NAND3X1_22 ( .A(_247_), .B(_249_), .C(_248_), .Y(_250_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_244_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_245_) );
OAI21X1 OAI21X1_73 ( .A(_244_), .B(_245_), .C(_18__1_), .Y(_246_) );
NAND2X1 NAND2X1_74 ( .A(_246_), .B(_250_), .Y(_16__1_) );
OAI21X1 OAI21X1_74 ( .A(_247_), .B(_244_), .C(_249_), .Y(_18__2_) );
INVX1 INVX1_53 ( .A(_18__2_), .Y(_254_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_255_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_256_) );
NAND3X1 NAND3X1_23 ( .A(_254_), .B(_256_), .C(_255_), .Y(_257_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_251_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_252_) );
OAI21X1 OAI21X1_75 ( .A(_251_), .B(_252_), .C(_18__2_), .Y(_253_) );
NAND2X1 NAND2X1_76 ( .A(_253_), .B(_257_), .Y(_16__2_) );
OAI21X1 OAI21X1_76 ( .A(_254_), .B(_251_), .C(_256_), .Y(_18__3_) );
INVX1 INVX1_54 ( .A(_18__3_), .Y(_261_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_262_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_263_) );
NAND3X1 NAND3X1_24 ( .A(_261_), .B(_263_), .C(_262_), .Y(_264_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_258_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_259_) );
OAI21X1 OAI21X1_77 ( .A(_258_), .B(_259_), .C(_18__3_), .Y(_260_) );
NAND2X1 NAND2X1_78 ( .A(_260_), .B(_264_), .Y(_16__3_) );
OAI21X1 OAI21X1_78 ( .A(_261_), .B(_258_), .C(_263_), .Y(_14_) );
INVX1 INVX1_55 ( .A(1'b0), .Y(_268_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_269_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_270_) );
NAND3X1 NAND3X1_25 ( .A(_268_), .B(_270_), .C(_269_), .Y(_271_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_265_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_266_) );
OAI21X1 OAI21X1_79 ( .A(_265_), .B(_266_), .C(1'b0), .Y(_267_) );
NAND2X1 NAND2X1_80 ( .A(_267_), .B(_271_), .Y(_21__0_) );
OAI21X1 OAI21X1_80 ( .A(_268_), .B(_265_), .C(_270_), .Y(_23__1_) );
INVX1 INVX1_56 ( .A(_23__1_), .Y(_275_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_276_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_277_) );
NAND3X1 NAND3X1_26 ( .A(_275_), .B(_277_), .C(_276_), .Y(_278_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_272_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_273_) );
OAI21X1 OAI21X1_81 ( .A(_272_), .B(_273_), .C(_23__1_), .Y(_274_) );
NAND2X1 NAND2X1_82 ( .A(_274_), .B(_278_), .Y(_21__1_) );
OAI21X1 OAI21X1_82 ( .A(_275_), .B(_272_), .C(_277_), .Y(_23__2_) );
INVX1 INVX1_57 ( .A(_23__2_), .Y(_282_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_283_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_284_) );
NAND3X1 NAND3X1_27 ( .A(_282_), .B(_284_), .C(_283_), .Y(_285_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_279_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_280_) );
OAI21X1 OAI21X1_83 ( .A(_279_), .B(_280_), .C(_23__2_), .Y(_281_) );
NAND2X1 NAND2X1_84 ( .A(_281_), .B(_285_), .Y(_21__2_) );
OAI21X1 OAI21X1_84 ( .A(_282_), .B(_279_), .C(_284_), .Y(_23__3_) );
INVX1 INVX1_58 ( .A(_23__3_), .Y(_289_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_290_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_291_) );
NAND3X1 NAND3X1_28 ( .A(_289_), .B(_291_), .C(_290_), .Y(_292_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_286_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_287_) );
OAI21X1 OAI21X1_85 ( .A(_286_), .B(_287_), .C(_23__3_), .Y(_288_) );
NAND2X1 NAND2X1_86 ( .A(_288_), .B(_292_), .Y(_21__3_) );
OAI21X1 OAI21X1_86 ( .A(_289_), .B(_286_), .C(_291_), .Y(_19_) );
INVX1 INVX1_59 ( .A(1'b1), .Y(_296_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_297_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_298_) );
NAND3X1 NAND3X1_29 ( .A(_296_), .B(_298_), .C(_297_), .Y(_299_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_293_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_294_) );
OAI21X1 OAI21X1_87 ( .A(_293_), .B(_294_), .C(1'b1), .Y(_295_) );
NAND2X1 NAND2X1_88 ( .A(_295_), .B(_299_), .Y(_22__0_) );
OAI21X1 OAI21X1_88 ( .A(_296_), .B(_293_), .C(_298_), .Y(_24__1_) );
INVX1 INVX1_60 ( .A(_24__1_), .Y(_303_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_304_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_305_) );
NAND3X1 NAND3X1_30 ( .A(_303_), .B(_305_), .C(_304_), .Y(_306_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_300_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_301_) );
OAI21X1 OAI21X1_89 ( .A(_300_), .B(_301_), .C(_24__1_), .Y(_302_) );
NAND2X1 NAND2X1_90 ( .A(_302_), .B(_306_), .Y(_22__1_) );
OAI21X1 OAI21X1_90 ( .A(_303_), .B(_300_), .C(_305_), .Y(_24__2_) );
INVX1 INVX1_61 ( .A(_24__2_), .Y(_310_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_311_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_312_) );
NAND3X1 NAND3X1_31 ( .A(_310_), .B(_312_), .C(_311_), .Y(_313_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_307_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_308_) );
OAI21X1 OAI21X1_91 ( .A(_307_), .B(_308_), .C(_24__2_), .Y(_309_) );
NAND2X1 NAND2X1_92 ( .A(_309_), .B(_313_), .Y(_22__2_) );
OAI21X1 OAI21X1_92 ( .A(_310_), .B(_307_), .C(_312_), .Y(_24__3_) );
INVX1 INVX1_62 ( .A(_24__3_), .Y(_317_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_318_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_319_) );
NAND3X1 NAND3X1_32 ( .A(_317_), .B(_319_), .C(_318_), .Y(_320_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_314_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_315_) );
OAI21X1 OAI21X1_93 ( .A(_314_), .B(_315_), .C(_24__3_), .Y(_316_) );
NAND2X1 NAND2X1_94 ( .A(_316_), .B(_320_), .Y(_22__3_) );
OAI21X1 OAI21X1_94 ( .A(_317_), .B(_314_), .C(_319_), .Y(_20_) );
INVX1 INVX1_63 ( .A(1'b0), .Y(_324_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_325_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_326_) );
NAND3X1 NAND3X1_33 ( .A(_324_), .B(_326_), .C(_325_), .Y(_327_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_321_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_322_) );
OAI21X1 OAI21X1_95 ( .A(_321_), .B(_322_), .C(1'b0), .Y(_323_) );
NAND2X1 NAND2X1_96 ( .A(_323_), .B(_327_), .Y(_27__0_) );
OAI21X1 OAI21X1_96 ( .A(_324_), .B(_321_), .C(_326_), .Y(_29__1_) );
INVX1 INVX1_64 ( .A(_29__1_), .Y(_331_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_332_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_333_) );
NAND3X1 NAND3X1_34 ( .A(_331_), .B(_333_), .C(_332_), .Y(_334_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_328_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_329_) );
OAI21X1 OAI21X1_97 ( .A(_328_), .B(_329_), .C(_29__1_), .Y(_330_) );
NAND2X1 NAND2X1_98 ( .A(_330_), .B(_334_), .Y(_27__1_) );
OAI21X1 OAI21X1_98 ( .A(_331_), .B(_328_), .C(_333_), .Y(_29__2_) );
INVX1 INVX1_65 ( .A(_29__2_), .Y(_338_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_339_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_340_) );
NAND3X1 NAND3X1_35 ( .A(_338_), .B(_340_), .C(_339_), .Y(_341_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_335_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_336_) );
OAI21X1 OAI21X1_99 ( .A(_335_), .B(_336_), .C(_29__2_), .Y(_337_) );
NAND2X1 NAND2X1_100 ( .A(_337_), .B(_341_), .Y(_27__2_) );
OAI21X1 OAI21X1_100 ( .A(_338_), .B(_335_), .C(_340_), .Y(_29__3_) );
INVX1 INVX1_66 ( .A(_29__3_), .Y(_345_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_346_) );
NAND2X1 NAND2X1_101 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_347_) );
NAND3X1 NAND3X1_36 ( .A(_345_), .B(_347_), .C(_346_), .Y(_348_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_342_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_343_) );
OAI21X1 OAI21X1_101 ( .A(_342_), .B(_343_), .C(_29__3_), .Y(_344_) );
NAND2X1 NAND2X1_102 ( .A(_344_), .B(_348_), .Y(_27__3_) );
OAI21X1 OAI21X1_102 ( .A(_345_), .B(_342_), .C(_347_), .Y(_25_) );
INVX1 INVX1_67 ( .A(1'b1), .Y(_352_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_353_) );
NAND2X1 NAND2X1_103 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_354_) );
NAND3X1 NAND3X1_37 ( .A(_352_), .B(_354_), .C(_353_), .Y(_355_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_349_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_350_) );
OAI21X1 OAI21X1_103 ( .A(_349_), .B(_350_), .C(1'b1), .Y(_351_) );
NAND2X1 NAND2X1_104 ( .A(_351_), .B(_355_), .Y(_28__0_) );
OAI21X1 OAI21X1_104 ( .A(_352_), .B(_349_), .C(_354_), .Y(_30__1_) );
INVX1 INVX1_68 ( .A(_30__1_), .Y(_359_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_360_) );
NAND2X1 NAND2X1_105 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_361_) );
NAND3X1 NAND3X1_38 ( .A(_359_), .B(_361_), .C(_360_), .Y(_362_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_356_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_357_) );
OAI21X1 OAI21X1_105 ( .A(_356_), .B(_357_), .C(_30__1_), .Y(_358_) );
NAND2X1 NAND2X1_106 ( .A(_358_), .B(_362_), .Y(_28__1_) );
OAI21X1 OAI21X1_106 ( .A(_359_), .B(_356_), .C(_361_), .Y(_30__2_) );
INVX1 INVX1_69 ( .A(_30__2_), .Y(_366_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_367_) );
NAND2X1 NAND2X1_107 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_368_) );
NAND3X1 NAND3X1_39 ( .A(_366_), .B(_368_), .C(_367_), .Y(_369_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_363_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_364_) );
OAI21X1 OAI21X1_107 ( .A(_363_), .B(_364_), .C(_30__2_), .Y(_365_) );
NAND2X1 NAND2X1_108 ( .A(_365_), .B(_369_), .Y(_28__2_) );
OAI21X1 OAI21X1_108 ( .A(_366_), .B(_363_), .C(_368_), .Y(_30__3_) );
INVX1 INVX1_70 ( .A(_30__3_), .Y(_373_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_374_) );
NAND2X1 NAND2X1_109 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_375_) );
NAND3X1 NAND3X1_40 ( .A(_373_), .B(_375_), .C(_374_), .Y(_376_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_370_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_371_) );
OAI21X1 OAI21X1_109 ( .A(_370_), .B(_371_), .C(_30__3_), .Y(_372_) );
NAND2X1 NAND2X1_110 ( .A(_372_), .B(_376_), .Y(_28__3_) );
OAI21X1 OAI21X1_110 ( .A(_373_), .B(_370_), .C(_375_), .Y(_26_) );
INVX1 INVX1_71 ( .A(1'b0), .Y(_380_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_381_) );
NAND2X1 NAND2X1_111 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_382_) );
NAND3X1 NAND3X1_41 ( .A(_380_), .B(_382_), .C(_381_), .Y(_383_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_377_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_378_) );
OAI21X1 OAI21X1_111 ( .A(_377_), .B(_378_), .C(1'b0), .Y(_379_) );
NAND2X1 NAND2X1_112 ( .A(_379_), .B(_383_), .Y(_33__0_) );
OAI21X1 OAI21X1_112 ( .A(_380_), .B(_377_), .C(_382_), .Y(_35__1_) );
INVX1 INVX1_72 ( .A(_35__1_), .Y(_387_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_388_) );
NAND2X1 NAND2X1_113 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_389_) );
NAND3X1 NAND3X1_42 ( .A(_387_), .B(_389_), .C(_388_), .Y(_390_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_384_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_385_) );
OAI21X1 OAI21X1_113 ( .A(_384_), .B(_385_), .C(_35__1_), .Y(_386_) );
NAND2X1 NAND2X1_114 ( .A(_386_), .B(_390_), .Y(_33__1_) );
OAI21X1 OAI21X1_114 ( .A(_387_), .B(_384_), .C(_389_), .Y(_35__2_) );
INVX1 INVX1_73 ( .A(_35__2_), .Y(_394_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_395_) );
NAND2X1 NAND2X1_115 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_396_) );
NAND3X1 NAND3X1_43 ( .A(_394_), .B(_396_), .C(_395_), .Y(_397_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_391_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_392_) );
OAI21X1 OAI21X1_115 ( .A(_391_), .B(_392_), .C(_35__2_), .Y(_393_) );
NAND2X1 NAND2X1_116 ( .A(_393_), .B(_397_), .Y(_33__2_) );
OAI21X1 OAI21X1_116 ( .A(_394_), .B(_391_), .C(_396_), .Y(_35__3_) );
INVX1 INVX1_74 ( .A(_35__3_), .Y(_401_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_402_) );
NAND2X1 NAND2X1_117 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_403_) );
NAND3X1 NAND3X1_44 ( .A(_401_), .B(_403_), .C(_402_), .Y(_404_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_398_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_399_) );
OAI21X1 OAI21X1_117 ( .A(_398_), .B(_399_), .C(_35__3_), .Y(_400_) );
NAND2X1 NAND2X1_118 ( .A(_400_), .B(_404_), .Y(_33__3_) );
OAI21X1 OAI21X1_118 ( .A(_401_), .B(_398_), .C(_403_), .Y(_31_) );
INVX1 INVX1_75 ( .A(1'b1), .Y(_408_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_409_) );
NAND2X1 NAND2X1_119 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_410_) );
NAND3X1 NAND3X1_45 ( .A(_408_), .B(_410_), .C(_409_), .Y(_411_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_405_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_406_) );
OAI21X1 OAI21X1_119 ( .A(_405_), .B(_406_), .C(1'b1), .Y(_407_) );
NAND2X1 NAND2X1_120 ( .A(_407_), .B(_411_), .Y(_34__0_) );
OAI21X1 OAI21X1_120 ( .A(_408_), .B(_405_), .C(_410_), .Y(_36__1_) );
INVX1 INVX1_76 ( .A(_36__1_), .Y(_415_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_416_) );
NAND2X1 NAND2X1_121 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_417_) );
NAND3X1 NAND3X1_46 ( .A(_415_), .B(_417_), .C(_416_), .Y(_418_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_412_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_413_) );
OAI21X1 OAI21X1_121 ( .A(_412_), .B(_413_), .C(_36__1_), .Y(_414_) );
NAND2X1 NAND2X1_122 ( .A(_414_), .B(_418_), .Y(_34__1_) );
OAI21X1 OAI21X1_122 ( .A(_415_), .B(_412_), .C(_417_), .Y(_36__2_) );
INVX1 INVX1_77 ( .A(_36__2_), .Y(_422_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_423_) );
NAND2X1 NAND2X1_123 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_424_) );
NAND3X1 NAND3X1_47 ( .A(_422_), .B(_424_), .C(_423_), .Y(_425_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_419_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_420_) );
OAI21X1 OAI21X1_123 ( .A(_419_), .B(_420_), .C(_36__2_), .Y(_421_) );
NAND2X1 NAND2X1_124 ( .A(_421_), .B(_425_), .Y(_34__2_) );
OAI21X1 OAI21X1_124 ( .A(_422_), .B(_419_), .C(_424_), .Y(_36__3_) );
INVX1 INVX1_78 ( .A(_36__3_), .Y(_429_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_430_) );
NAND2X1 NAND2X1_125 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_431_) );
NAND3X1 NAND3X1_48 ( .A(_429_), .B(_431_), .C(_430_), .Y(_432_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_426_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_427_) );
OAI21X1 OAI21X1_125 ( .A(_426_), .B(_427_), .C(_36__3_), .Y(_428_) );
NAND2X1 NAND2X1_126 ( .A(_428_), .B(_432_), .Y(_34__3_) );
OAI21X1 OAI21X1_126 ( .A(_429_), .B(_426_), .C(_431_), .Y(_32_) );
INVX1 INVX1_79 ( .A(1'b0), .Y(_436_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_437_) );
NAND2X1 NAND2X1_127 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_438_) );
NAND3X1 NAND3X1_49 ( .A(_436_), .B(_438_), .C(_437_), .Y(_439_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_433_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_434_) );
OAI21X1 OAI21X1_127 ( .A(_433_), .B(_434_), .C(1'b0), .Y(_435_) );
NAND2X1 NAND2X1_128 ( .A(_435_), .B(_439_), .Y(rca_inst_w_SUM) );
BUFX2 BUFX2_27 ( .A(rca_inst_w_SUM), .Y(_0__0_) );
BUFX2 BUFX2_28 ( .A(1'b0), .Y(_5__0_) );
BUFX2 BUFX2_29 ( .A(_1_), .Y(_5__4_) );
BUFX2 BUFX2_30 ( .A(1'b1), .Y(_6__0_) );
BUFX2 BUFX2_31 ( .A(_2_), .Y(_6__4_) );
BUFX2 BUFX2_32 ( .A(1'b0), .Y(_11__0_) );
BUFX2 BUFX2_33 ( .A(_7_), .Y(_11__4_) );
BUFX2 BUFX2_34 ( .A(1'b1), .Y(_12__0_) );
BUFX2 BUFX2_35 ( .A(_8_), .Y(_12__4_) );
BUFX2 BUFX2_36 ( .A(1'b0), .Y(_17__0_) );
BUFX2 BUFX2_37 ( .A(_13_), .Y(_17__4_) );
BUFX2 BUFX2_38 ( .A(1'b1), .Y(_18__0_) );
BUFX2 BUFX2_39 ( .A(_14_), .Y(_18__4_) );
BUFX2 BUFX2_40 ( .A(1'b0), .Y(_23__0_) );
BUFX2 BUFX2_41 ( .A(_19_), .Y(_23__4_) );
BUFX2 BUFX2_42 ( .A(1'b1), .Y(_24__0_) );
BUFX2 BUFX2_43 ( .A(_20_), .Y(_24__4_) );
BUFX2 BUFX2_44 ( .A(1'b0), .Y(_29__0_) );
BUFX2 BUFX2_45 ( .A(_25_), .Y(_29__4_) );
BUFX2 BUFX2_46 ( .A(1'b1), .Y(_30__0_) );
BUFX2 BUFX2_47 ( .A(_26_), .Y(_30__4_) );
BUFX2 BUFX2_48 ( .A(1'b0), .Y(_35__0_) );
BUFX2 BUFX2_49 ( .A(_31_), .Y(_35__4_) );
BUFX2 BUFX2_50 ( .A(1'b1), .Y(_36__0_) );
BUFX2 BUFX2_51 ( .A(_32_), .Y(_36__4_) );
BUFX2 BUFX2_52 ( .A(1'b0), .Y(w_cout_0_) );
endmodule
