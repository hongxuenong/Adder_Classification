module cla_11bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [10:0] i_add1;
input [10:0] i_add2;
output [11:0] o_result;

NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(w_C_1_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_1_), .Y(_2_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .C(_2_), .Y(_3_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_3_), .Y(w_C_2_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_4_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_5_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_6_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_6_), .C(_2_), .Y(_7_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_7_), .Y(w_C_3_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .Y(_8_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add1[3]), .Y(_9_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_9_), .Y(_10_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_11_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_11_), .C(_7_), .Y(_12_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_10_), .Y(w_C_4_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_13_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_14_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_14_), .C(_12_), .Y(_15_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_15_), .Y(w_C_5_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_16_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(_17_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_18_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_18_), .C(_15_), .Y(_19_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_17_), .Y(w_C_6_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .Y(_20_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add1[6]), .Y(_21_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_23_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_23_), .C(_19_), .Y(_24_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .C(_24_), .Y(w_C_7_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .Y(_25_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(_26_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_27_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(_28_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_28_), .C(_24_), .Y(_29_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .C(_29_), .Y(_30_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(w_C_8_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_31_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_32_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_30_), .C(_31_), .Y(w_C_9_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_33_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_34_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_34_), .Y(_35_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_32_), .Y(_36_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_36_), .C(_29_), .Y(_37_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_38_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_38_), .C(_37_), .Y(_39_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_33_), .Y(w_C_10_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_40_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_41_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_41_), .C(_39_), .Y(_42_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_42_), .Y(w_C_11_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_43__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_43__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_43__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_43__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_43__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_43__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_43__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_43__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_43__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_43__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_43__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(o_result[11]) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_47_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_48_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_49_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_49_), .C(_48_), .Y(_50_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_44_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_45_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_45_), .C(w_C_4_), .Y(_46_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_50_), .Y(_43__4_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_54_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_55_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_56_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_56_), .C(_55_), .Y(_57_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_51_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_52_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_52_), .C(w_C_5_), .Y(_53_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_57_), .Y(_43__5_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_61_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_62_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_63_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_63_), .C(_62_), .Y(_64_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_58_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_59_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_59_), .C(w_C_6_), .Y(_60_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_64_), .Y(_43__6_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_68_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_69_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_70_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_70_), .C(_69_), .Y(_71_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_65_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_66_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_66_), .C(w_C_7_), .Y(_67_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_71_), .Y(_43__7_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_75_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_76_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_77_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_77_), .C(_76_), .Y(_78_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_72_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_73_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_73_), .C(w_C_8_), .Y(_74_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_78_), .Y(_43__8_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_82_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_83_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_84_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_84_), .C(_83_), .Y(_85_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_79_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_80_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_80_), .C(w_C_9_), .Y(_81_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_85_), .Y(_43__9_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_89_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_90_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_91_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_91_), .C(_90_), .Y(_92_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_86_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_87_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_87_), .C(w_C_10_), .Y(_88_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_92_), .Y(_43__10_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_96_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_97_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_98_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_98_), .C(_97_), .Y(_99_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_93_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_94_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_94_), .C(gnd), .Y(_95_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_99_), .Y(_43__0_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_103_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_104_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_105_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_105_), .C(_104_), .Y(_106_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_100_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_101_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_101_), .C(w_C_1_), .Y(_102_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_106_), .Y(_43__1_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_110_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_111_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_112_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_112_), .C(_111_), .Y(_113_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_107_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_108_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_108_), .C(w_C_2_), .Y(_109_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_113_), .Y(_43__2_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_117_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_118_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_119_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_119_), .C(_118_), .Y(_120_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_114_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_115_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_115_), .C(w_C_3_), .Y(_116_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_120_), .Y(_43__3_) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_43__11_) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
