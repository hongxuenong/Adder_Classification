module CSkipA_4bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [3:0] i_add_term1;
input [3:0] i_add_term2;
output [3:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

NOR2X1 NOR2X1_1 ( .A(_37_), .B(_42_), .Y(skip0_P) );
INVX1 INVX1_1 ( .A(cout0), .Y(_43_) );
NAND2X1 NAND2X1_1 ( .A(gnd), .B(skip0_P), .Y(_44_) );
OAI21X1 OAI21X1_1 ( .A(skip0_P), .B(_43_), .C(_44_), .Y(_0_) );
BUFX2 BUFX2_1 ( .A(_0_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
INVX1 INVX1_2 ( .A(gnd), .Y(_4_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_5_) );
NAND2X1 NAND2X1_2 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_6_) );
NAND3X1 NAND3X1_1 ( .A(_4_), .B(_6_), .C(_5_), .Y(_7_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_1_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_2_) );
OAI21X1 OAI21X1_2 ( .A(_1_), .B(_2_), .C(gnd), .Y(_3_) );
NAND2X1 NAND2X1_3 ( .A(_3_), .B(_7_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_3 ( .A(_4_), .B(_1_), .C(_6_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_3 ( .A(rca_inst_fa3_i_carry), .Y(_11_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_12_) );
NAND2X1 NAND2X1_4 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_13_) );
NAND3X1 NAND3X1_2 ( .A(_11_), .B(_13_), .C(_12_), .Y(_14_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_8_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_9_) );
OAI21X1 OAI21X1_4 ( .A(_8_), .B(_9_), .C(rca_inst_fa3_i_carry), .Y(_10_) );
NAND2X1 NAND2X1_5 ( .A(_10_), .B(_14_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_5 ( .A(_11_), .B(_8_), .C(_13_), .Y(cout0) );
INVX1 INVX1_4 ( .A(rca_inst_fa0_o_carry), .Y(_18_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_19_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_20_) );
NAND3X1 NAND3X1_3 ( .A(_18_), .B(_20_), .C(_19_), .Y(_21_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_15_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_16_) );
OAI21X1 OAI21X1_6 ( .A(_15_), .B(_16_), .C(rca_inst_fa0_o_carry), .Y(_17_) );
NAND2X1 NAND2X1_7 ( .A(_17_), .B(_21_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_7 ( .A(_18_), .B(_15_), .C(_20_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_5 ( .A(rca_inst_fa_1__o_carry), .Y(_25_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_26_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_27_) );
NAND3X1 NAND3X1_4 ( .A(_25_), .B(_27_), .C(_26_), .Y(_28_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_22_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_23_) );
OAI21X1 OAI21X1_8 ( .A(_22_), .B(_23_), .C(rca_inst_fa_1__o_carry), .Y(_24_) );
NAND2X1 NAND2X1_9 ( .A(_24_), .B(_28_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_9 ( .A(_25_), .B(_22_), .C(_27_), .Y(rca_inst_fa3_i_carry) );
INVX1 INVX1_6 ( .A(i_add_term1[0]), .Y(_29_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[0]), .B(_29_), .Y(_30_) );
INVX1 INVX1_7 ( .A(i_add_term2[0]), .Y(_31_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term1[0]), .B(_31_), .Y(_32_) );
INVX1 INVX1_8 ( .A(i_add_term1[1]), .Y(_33_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[1]), .B(_33_), .Y(_34_) );
INVX1 INVX1_9 ( .A(i_add_term2[1]), .Y(_35_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term1[1]), .B(_35_), .Y(_36_) );
OAI22X1 OAI22X1_1 ( .A(_30_), .B(_32_), .C(_34_), .D(_36_), .Y(_37_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_38_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_39_) );
NOR2X1 NOR2X1_11 ( .A(_38_), .B(_39_), .Y(_40_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_41_) );
NAND2X1 NAND2X1_10 ( .A(_40_), .B(_41_), .Y(_42_) );
endmodule
