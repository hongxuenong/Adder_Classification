module csa_51bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term1[45], i_add_term1[46], i_add_term1[47], i_add_term1[48], i_add_term1[49], i_add_term1[50], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], i_add_term2[45], i_add_term2[46], i_add_term2[47], i_add_term2[48], i_add_term2[49], i_add_term2[50], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], sum[45], sum[46], sum[47], sum[48], sum[49], sum[50], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term1[45];
input i_add_term1[46];
input i_add_term1[47];
input i_add_term1[48];
input i_add_term1[49];
input i_add_term1[50];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
input i_add_term2[45];
input i_add_term2[46];
input i_add_term2[47];
input i_add_term2[48];
input i_add_term2[49];
input i_add_term2[50];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output sum[45];
output sum[46];
output sum[47];
output sum[48];
output sum[49];
output sum[50];
output cout;

OAI21X1 OAI21X1_1 ( .A(w_cout_4_), .B(_113_), .C(_114_), .Y(w_cout_5_) );
INVX1 INVX1_1 ( .A(_27__0_), .Y(_115_) );
NAND2X1 NAND2X1_1 ( .A(_28__0_), .B(w_cout_4_), .Y(_116_) );
OAI21X1 OAI21X1_2 ( .A(w_cout_4_), .B(_115_), .C(_116_), .Y(_0__19_) );
INVX1 INVX1_2 ( .A(_27__1_), .Y(_117_) );
NAND2X1 NAND2X1_2 ( .A(w_cout_4_), .B(_28__1_), .Y(_118_) );
OAI21X1 OAI21X1_3 ( .A(w_cout_4_), .B(_117_), .C(_118_), .Y(_0__20_) );
INVX1 INVX1_3 ( .A(_27__2_), .Y(_119_) );
NAND2X1 NAND2X1_3 ( .A(w_cout_4_), .B(_28__2_), .Y(_120_) );
OAI21X1 OAI21X1_4 ( .A(w_cout_4_), .B(_119_), .C(_120_), .Y(_0__21_) );
INVX1 INVX1_4 ( .A(_27__3_), .Y(_121_) );
NAND2X1 NAND2X1_4 ( .A(w_cout_4_), .B(_28__3_), .Y(_122_) );
OAI21X1 OAI21X1_5 ( .A(w_cout_4_), .B(_121_), .C(_122_), .Y(_0__22_) );
INVX1 INVX1_5 ( .A(_31_), .Y(_123_) );
NAND2X1 NAND2X1_5 ( .A(_32_), .B(w_cout_5_), .Y(_124_) );
OAI21X1 OAI21X1_6 ( .A(w_cout_5_), .B(_123_), .C(_124_), .Y(w_cout_6_) );
INVX1 INVX1_6 ( .A(_33__0_), .Y(_125_) );
NAND2X1 NAND2X1_6 ( .A(_34__0_), .B(w_cout_5_), .Y(_126_) );
OAI21X1 OAI21X1_7 ( .A(w_cout_5_), .B(_125_), .C(_126_), .Y(_0__23_) );
INVX1 INVX1_7 ( .A(_33__1_), .Y(_127_) );
NAND2X1 NAND2X1_7 ( .A(w_cout_5_), .B(_34__1_), .Y(_128_) );
OAI21X1 OAI21X1_8 ( .A(w_cout_5_), .B(_127_), .C(_128_), .Y(_0__24_) );
INVX1 INVX1_8 ( .A(_33__2_), .Y(_129_) );
NAND2X1 NAND2X1_8 ( .A(w_cout_5_), .B(_34__2_), .Y(_130_) );
OAI21X1 OAI21X1_9 ( .A(w_cout_5_), .B(_129_), .C(_130_), .Y(_0__25_) );
INVX1 INVX1_9 ( .A(_33__3_), .Y(_131_) );
NAND2X1 NAND2X1_9 ( .A(w_cout_5_), .B(_34__3_), .Y(_132_) );
OAI21X1 OAI21X1_10 ( .A(w_cout_5_), .B(_131_), .C(_132_), .Y(_0__26_) );
INVX1 INVX1_10 ( .A(_37_), .Y(_133_) );
NAND2X1 NAND2X1_10 ( .A(_38_), .B(w_cout_6_), .Y(_134_) );
OAI21X1 OAI21X1_11 ( .A(w_cout_6_), .B(_133_), .C(_134_), .Y(w_cout_7_) );
INVX1 INVX1_11 ( .A(_39__0_), .Y(_135_) );
NAND2X1 NAND2X1_11 ( .A(_40__0_), .B(w_cout_6_), .Y(_136_) );
OAI21X1 OAI21X1_12 ( .A(w_cout_6_), .B(_135_), .C(_136_), .Y(_0__27_) );
INVX1 INVX1_12 ( .A(_39__1_), .Y(_137_) );
NAND2X1 NAND2X1_12 ( .A(w_cout_6_), .B(_40__1_), .Y(_138_) );
OAI21X1 OAI21X1_13 ( .A(w_cout_6_), .B(_137_), .C(_138_), .Y(_0__28_) );
INVX1 INVX1_13 ( .A(_39__2_), .Y(_139_) );
NAND2X1 NAND2X1_13 ( .A(w_cout_6_), .B(_40__2_), .Y(_140_) );
OAI21X1 OAI21X1_14 ( .A(w_cout_6_), .B(_139_), .C(_140_), .Y(_0__29_) );
INVX1 INVX1_14 ( .A(_39__3_), .Y(_141_) );
NAND2X1 NAND2X1_14 ( .A(w_cout_6_), .B(_40__3_), .Y(_142_) );
OAI21X1 OAI21X1_15 ( .A(w_cout_6_), .B(_141_), .C(_142_), .Y(_0__30_) );
INVX1 INVX1_15 ( .A(_43_), .Y(_143_) );
NAND2X1 NAND2X1_15 ( .A(_44_), .B(w_cout_7_), .Y(_144_) );
OAI21X1 OAI21X1_16 ( .A(w_cout_7_), .B(_143_), .C(_144_), .Y(w_cout_8_) );
INVX1 INVX1_16 ( .A(_45__0_), .Y(_145_) );
NAND2X1 NAND2X1_16 ( .A(_46__0_), .B(w_cout_7_), .Y(_146_) );
OAI21X1 OAI21X1_17 ( .A(w_cout_7_), .B(_145_), .C(_146_), .Y(_0__31_) );
INVX1 INVX1_17 ( .A(_45__1_), .Y(_147_) );
NAND2X1 NAND2X1_17 ( .A(w_cout_7_), .B(_46__1_), .Y(_148_) );
OAI21X1 OAI21X1_18 ( .A(w_cout_7_), .B(_147_), .C(_148_), .Y(_0__32_) );
INVX1 INVX1_18 ( .A(_45__2_), .Y(_149_) );
NAND2X1 NAND2X1_18 ( .A(w_cout_7_), .B(_46__2_), .Y(_150_) );
OAI21X1 OAI21X1_19 ( .A(w_cout_7_), .B(_149_), .C(_150_), .Y(_0__33_) );
INVX1 INVX1_19 ( .A(_45__3_), .Y(_151_) );
NAND2X1 NAND2X1_19 ( .A(w_cout_7_), .B(_46__3_), .Y(_152_) );
OAI21X1 OAI21X1_20 ( .A(w_cout_7_), .B(_151_), .C(_152_), .Y(_0__34_) );
INVX1 INVX1_20 ( .A(_49_), .Y(_153_) );
NAND2X1 NAND2X1_20 ( .A(_50_), .B(w_cout_8_), .Y(_154_) );
OAI21X1 OAI21X1_21 ( .A(w_cout_8_), .B(_153_), .C(_154_), .Y(w_cout_9_) );
INVX1 INVX1_21 ( .A(_51__0_), .Y(_155_) );
NAND2X1 NAND2X1_21 ( .A(_52__0_), .B(w_cout_8_), .Y(_156_) );
OAI21X1 OAI21X1_22 ( .A(w_cout_8_), .B(_155_), .C(_156_), .Y(_0__35_) );
INVX1 INVX1_22 ( .A(_51__1_), .Y(_157_) );
NAND2X1 NAND2X1_22 ( .A(w_cout_8_), .B(_52__1_), .Y(_158_) );
OAI21X1 OAI21X1_23 ( .A(w_cout_8_), .B(_157_), .C(_158_), .Y(_0__36_) );
INVX1 INVX1_23 ( .A(_51__2_), .Y(_159_) );
NAND2X1 NAND2X1_23 ( .A(w_cout_8_), .B(_52__2_), .Y(_160_) );
OAI21X1 OAI21X1_24 ( .A(w_cout_8_), .B(_159_), .C(_160_), .Y(_0__37_) );
INVX1 INVX1_24 ( .A(_51__3_), .Y(_161_) );
NAND2X1 NAND2X1_24 ( .A(w_cout_8_), .B(_52__3_), .Y(_162_) );
OAI21X1 OAI21X1_25 ( .A(w_cout_8_), .B(_161_), .C(_162_), .Y(_0__38_) );
INVX1 INVX1_25 ( .A(_55_), .Y(_163_) );
NAND2X1 NAND2X1_25 ( .A(_56_), .B(w_cout_9_), .Y(_164_) );
OAI21X1 OAI21X1_26 ( .A(w_cout_9_), .B(_163_), .C(_164_), .Y(w_cout_10_) );
INVX1 INVX1_26 ( .A(_57__0_), .Y(_165_) );
NAND2X1 NAND2X1_26 ( .A(_58__0_), .B(w_cout_9_), .Y(_166_) );
OAI21X1 OAI21X1_27 ( .A(w_cout_9_), .B(_165_), .C(_166_), .Y(_0__39_) );
INVX1 INVX1_27 ( .A(_57__1_), .Y(_167_) );
NAND2X1 NAND2X1_27 ( .A(w_cout_9_), .B(_58__1_), .Y(_168_) );
OAI21X1 OAI21X1_28 ( .A(w_cout_9_), .B(_167_), .C(_168_), .Y(_0__40_) );
INVX1 INVX1_28 ( .A(_57__2_), .Y(_169_) );
NAND2X1 NAND2X1_28 ( .A(w_cout_9_), .B(_58__2_), .Y(_170_) );
OAI21X1 OAI21X1_29 ( .A(w_cout_9_), .B(_169_), .C(_170_), .Y(_0__41_) );
INVX1 INVX1_29 ( .A(_57__3_), .Y(_171_) );
NAND2X1 NAND2X1_29 ( .A(w_cout_9_), .B(_58__3_), .Y(_172_) );
OAI21X1 OAI21X1_30 ( .A(w_cout_9_), .B(_171_), .C(_172_), .Y(_0__42_) );
INVX1 INVX1_30 ( .A(_61_), .Y(_173_) );
NAND2X1 NAND2X1_30 ( .A(_62_), .B(w_cout_10_), .Y(_174_) );
OAI21X1 OAI21X1_31 ( .A(w_cout_10_), .B(_173_), .C(_174_), .Y(w_cout_11_) );
INVX1 INVX1_31 ( .A(_63__0_), .Y(_175_) );
NAND2X1 NAND2X1_31 ( .A(_64__0_), .B(w_cout_10_), .Y(_176_) );
OAI21X1 OAI21X1_32 ( .A(w_cout_10_), .B(_175_), .C(_176_), .Y(_0__43_) );
INVX1 INVX1_32 ( .A(_63__1_), .Y(_177_) );
NAND2X1 NAND2X1_32 ( .A(w_cout_10_), .B(_64__1_), .Y(_178_) );
OAI21X1 OAI21X1_33 ( .A(w_cout_10_), .B(_177_), .C(_178_), .Y(_0__44_) );
INVX1 INVX1_33 ( .A(_63__2_), .Y(_179_) );
NAND2X1 NAND2X1_33 ( .A(w_cout_10_), .B(_64__2_), .Y(_180_) );
OAI21X1 OAI21X1_34 ( .A(w_cout_10_), .B(_179_), .C(_180_), .Y(_0__45_) );
INVX1 INVX1_34 ( .A(_63__3_), .Y(_181_) );
NAND2X1 NAND2X1_34 ( .A(w_cout_10_), .B(_64__3_), .Y(_182_) );
OAI21X1 OAI21X1_35 ( .A(w_cout_10_), .B(_181_), .C(_182_), .Y(_0__46_) );
INVX1 INVX1_35 ( .A(_67_), .Y(_183_) );
NAND2X1 NAND2X1_35 ( .A(_68_), .B(w_cout_11_), .Y(_184_) );
OAI21X1 OAI21X1_36 ( .A(w_cout_11_), .B(_183_), .C(_184_), .Y(w_cout_12_) );
INVX1 INVX1_36 ( .A(_69__0_), .Y(_185_) );
NAND2X1 NAND2X1_36 ( .A(_70__0_), .B(w_cout_11_), .Y(_186_) );
OAI21X1 OAI21X1_37 ( .A(w_cout_11_), .B(_185_), .C(_186_), .Y(_0__47_) );
INVX1 INVX1_37 ( .A(_69__1_), .Y(_187_) );
NAND2X1 NAND2X1_37 ( .A(w_cout_11_), .B(_70__1_), .Y(_188_) );
OAI21X1 OAI21X1_38 ( .A(w_cout_11_), .B(_187_), .C(_188_), .Y(_0__48_) );
INVX1 INVX1_38 ( .A(_69__2_), .Y(_189_) );
NAND2X1 NAND2X1_38 ( .A(w_cout_11_), .B(_70__2_), .Y(_190_) );
OAI21X1 OAI21X1_39 ( .A(w_cout_11_), .B(_189_), .C(_190_), .Y(_0__49_) );
INVX1 INVX1_39 ( .A(_69__3_), .Y(_191_) );
NAND2X1 NAND2X1_39 ( .A(w_cout_11_), .B(_70__3_), .Y(_192_) );
OAI21X1 OAI21X1_40 ( .A(w_cout_11_), .B(_191_), .C(_192_), .Y(_0__50_) );
INVX1 INVX1_40 ( .A(1'b0), .Y(_196_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_197_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_198_) );
NAND3X1 NAND3X1_1 ( .A(_196_), .B(_198_), .C(_197_), .Y(_199_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_193_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_194_) );
OAI21X1 OAI21X1_41 ( .A(_193_), .B(_194_), .C(1'b0), .Y(_195_) );
NAND2X1 NAND2X1_41 ( .A(_195_), .B(_199_), .Y(_3__0_) );
OAI21X1 OAI21X1_42 ( .A(_196_), .B(_193_), .C(_198_), .Y(_5__1_) );
INVX1 INVX1_41 ( .A(_5__1_), .Y(_203_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_204_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_205_) );
NAND3X1 NAND3X1_2 ( .A(_203_), .B(_205_), .C(_204_), .Y(_206_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_200_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_201_) );
OAI21X1 OAI21X1_43 ( .A(_200_), .B(_201_), .C(_5__1_), .Y(_202_) );
NAND2X1 NAND2X1_43 ( .A(_202_), .B(_206_), .Y(_3__1_) );
OAI21X1 OAI21X1_44 ( .A(_203_), .B(_200_), .C(_205_), .Y(_5__2_) );
INVX1 INVX1_42 ( .A(_5__2_), .Y(_210_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_211_) );
NAND2X1 NAND2X1_44 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_212_) );
NAND3X1 NAND3X1_3 ( .A(_210_), .B(_212_), .C(_211_), .Y(_213_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_207_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_208_) );
OAI21X1 OAI21X1_45 ( .A(_207_), .B(_208_), .C(_5__2_), .Y(_209_) );
NAND2X1 NAND2X1_45 ( .A(_209_), .B(_213_), .Y(_3__2_) );
OAI21X1 OAI21X1_46 ( .A(_210_), .B(_207_), .C(_212_), .Y(_5__3_) );
INVX1 INVX1_43 ( .A(_5__3_), .Y(_217_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_218_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_219_) );
NAND3X1 NAND3X1_4 ( .A(_217_), .B(_219_), .C(_218_), .Y(_220_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_214_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_215_) );
OAI21X1 OAI21X1_47 ( .A(_214_), .B(_215_), .C(_5__3_), .Y(_216_) );
NAND2X1 NAND2X1_47 ( .A(_216_), .B(_220_), .Y(_3__3_) );
OAI21X1 OAI21X1_48 ( .A(_217_), .B(_214_), .C(_219_), .Y(_1_) );
INVX1 INVX1_44 ( .A(1'b1), .Y(_224_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_225_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_226_) );
NAND3X1 NAND3X1_5 ( .A(_224_), .B(_226_), .C(_225_), .Y(_227_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_221_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_222_) );
OAI21X1 OAI21X1_49 ( .A(_221_), .B(_222_), .C(1'b1), .Y(_223_) );
NAND2X1 NAND2X1_49 ( .A(_223_), .B(_227_), .Y(_4__0_) );
OAI21X1 OAI21X1_50 ( .A(_224_), .B(_221_), .C(_226_), .Y(_6__1_) );
INVX1 INVX1_45 ( .A(_6__1_), .Y(_231_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_232_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_233_) );
NAND3X1 NAND3X1_6 ( .A(_231_), .B(_233_), .C(_232_), .Y(_234_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_228_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_229_) );
OAI21X1 OAI21X1_51 ( .A(_228_), .B(_229_), .C(_6__1_), .Y(_230_) );
NAND2X1 NAND2X1_51 ( .A(_230_), .B(_234_), .Y(_4__1_) );
OAI21X1 OAI21X1_52 ( .A(_231_), .B(_228_), .C(_233_), .Y(_6__2_) );
INVX1 INVX1_46 ( .A(_6__2_), .Y(_238_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_239_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_240_) );
NAND3X1 NAND3X1_7 ( .A(_238_), .B(_240_), .C(_239_), .Y(_241_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_235_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_236_) );
OAI21X1 OAI21X1_53 ( .A(_235_), .B(_236_), .C(_6__2_), .Y(_237_) );
NAND2X1 NAND2X1_53 ( .A(_237_), .B(_241_), .Y(_4__2_) );
OAI21X1 OAI21X1_54 ( .A(_238_), .B(_235_), .C(_240_), .Y(_6__3_) );
INVX1 INVX1_47 ( .A(_6__3_), .Y(_245_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_246_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_247_) );
NAND3X1 NAND3X1_8 ( .A(_245_), .B(_247_), .C(_246_), .Y(_248_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_242_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_243_) );
OAI21X1 OAI21X1_55 ( .A(_242_), .B(_243_), .C(_6__3_), .Y(_244_) );
NAND2X1 NAND2X1_55 ( .A(_244_), .B(_248_), .Y(_4__3_) );
OAI21X1 OAI21X1_56 ( .A(_245_), .B(_242_), .C(_247_), .Y(_2_) );
INVX1 INVX1_48 ( .A(1'b0), .Y(_252_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_253_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_254_) );
NAND3X1 NAND3X1_9 ( .A(_252_), .B(_254_), .C(_253_), .Y(_255_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_249_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_250_) );
OAI21X1 OAI21X1_57 ( .A(_249_), .B(_250_), .C(1'b0), .Y(_251_) );
NAND2X1 NAND2X1_57 ( .A(_251_), .B(_255_), .Y(_9__0_) );
OAI21X1 OAI21X1_58 ( .A(_252_), .B(_249_), .C(_254_), .Y(_11__1_) );
INVX1 INVX1_49 ( .A(_11__1_), .Y(_259_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_260_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_261_) );
NAND3X1 NAND3X1_10 ( .A(_259_), .B(_261_), .C(_260_), .Y(_262_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_256_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_257_) );
OAI21X1 OAI21X1_59 ( .A(_256_), .B(_257_), .C(_11__1_), .Y(_258_) );
NAND2X1 NAND2X1_59 ( .A(_258_), .B(_262_), .Y(_9__1_) );
OAI21X1 OAI21X1_60 ( .A(_259_), .B(_256_), .C(_261_), .Y(_11__2_) );
INVX1 INVX1_50 ( .A(_11__2_), .Y(_266_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_267_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_268_) );
NAND3X1 NAND3X1_11 ( .A(_266_), .B(_268_), .C(_267_), .Y(_269_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_263_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_264_) );
OAI21X1 OAI21X1_61 ( .A(_263_), .B(_264_), .C(_11__2_), .Y(_265_) );
NAND2X1 NAND2X1_61 ( .A(_265_), .B(_269_), .Y(_9__2_) );
OAI21X1 OAI21X1_62 ( .A(_266_), .B(_263_), .C(_268_), .Y(_11__3_) );
INVX1 INVX1_51 ( .A(_11__3_), .Y(_273_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_274_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_275_) );
NAND3X1 NAND3X1_12 ( .A(_273_), .B(_275_), .C(_274_), .Y(_276_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_270_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_271_) );
OAI21X1 OAI21X1_63 ( .A(_270_), .B(_271_), .C(_11__3_), .Y(_272_) );
NAND2X1 NAND2X1_63 ( .A(_272_), .B(_276_), .Y(_9__3_) );
OAI21X1 OAI21X1_64 ( .A(_273_), .B(_270_), .C(_275_), .Y(_7_) );
INVX1 INVX1_52 ( .A(1'b1), .Y(_280_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_281_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_282_) );
NAND3X1 NAND3X1_13 ( .A(_280_), .B(_282_), .C(_281_), .Y(_283_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_277_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_278_) );
OAI21X1 OAI21X1_65 ( .A(_277_), .B(_278_), .C(1'b1), .Y(_279_) );
NAND2X1 NAND2X1_65 ( .A(_279_), .B(_283_), .Y(_10__0_) );
OAI21X1 OAI21X1_66 ( .A(_280_), .B(_277_), .C(_282_), .Y(_12__1_) );
INVX1 INVX1_53 ( .A(_12__1_), .Y(_287_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_288_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_289_) );
NAND3X1 NAND3X1_14 ( .A(_287_), .B(_289_), .C(_288_), .Y(_290_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_284_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_285_) );
OAI21X1 OAI21X1_67 ( .A(_284_), .B(_285_), .C(_12__1_), .Y(_286_) );
NAND2X1 NAND2X1_67 ( .A(_286_), .B(_290_), .Y(_10__1_) );
OAI21X1 OAI21X1_68 ( .A(_287_), .B(_284_), .C(_289_), .Y(_12__2_) );
INVX1 INVX1_54 ( .A(_12__2_), .Y(_294_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_295_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_296_) );
NAND3X1 NAND3X1_15 ( .A(_294_), .B(_296_), .C(_295_), .Y(_297_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_291_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_292_) );
OAI21X1 OAI21X1_69 ( .A(_291_), .B(_292_), .C(_12__2_), .Y(_293_) );
NAND2X1 NAND2X1_69 ( .A(_293_), .B(_297_), .Y(_10__2_) );
OAI21X1 OAI21X1_70 ( .A(_294_), .B(_291_), .C(_296_), .Y(_12__3_) );
INVX1 INVX1_55 ( .A(_12__3_), .Y(_301_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_302_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_303_) );
NAND3X1 NAND3X1_16 ( .A(_301_), .B(_303_), .C(_302_), .Y(_304_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_298_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_299_) );
OAI21X1 OAI21X1_71 ( .A(_298_), .B(_299_), .C(_12__3_), .Y(_300_) );
NAND2X1 NAND2X1_71 ( .A(_300_), .B(_304_), .Y(_10__3_) );
OAI21X1 OAI21X1_72 ( .A(_301_), .B(_298_), .C(_303_), .Y(_8_) );
INVX1 INVX1_56 ( .A(1'b0), .Y(_308_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_309_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_310_) );
NAND3X1 NAND3X1_17 ( .A(_308_), .B(_310_), .C(_309_), .Y(_311_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_305_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_306_) );
OAI21X1 OAI21X1_73 ( .A(_305_), .B(_306_), .C(1'b0), .Y(_307_) );
NAND2X1 NAND2X1_73 ( .A(_307_), .B(_311_), .Y(_15__0_) );
OAI21X1 OAI21X1_74 ( .A(_308_), .B(_305_), .C(_310_), .Y(_17__1_) );
INVX1 INVX1_57 ( .A(_17__1_), .Y(_315_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_316_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_317_) );
NAND3X1 NAND3X1_18 ( .A(_315_), .B(_317_), .C(_316_), .Y(_318_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_312_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_313_) );
OAI21X1 OAI21X1_75 ( .A(_312_), .B(_313_), .C(_17__1_), .Y(_314_) );
NAND2X1 NAND2X1_75 ( .A(_314_), .B(_318_), .Y(_15__1_) );
OAI21X1 OAI21X1_76 ( .A(_315_), .B(_312_), .C(_317_), .Y(_17__2_) );
INVX1 INVX1_58 ( .A(_17__2_), .Y(_322_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_323_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_324_) );
NAND3X1 NAND3X1_19 ( .A(_322_), .B(_324_), .C(_323_), .Y(_325_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_319_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_320_) );
OAI21X1 OAI21X1_77 ( .A(_319_), .B(_320_), .C(_17__2_), .Y(_321_) );
NAND2X1 NAND2X1_77 ( .A(_321_), .B(_325_), .Y(_15__2_) );
OAI21X1 OAI21X1_78 ( .A(_322_), .B(_319_), .C(_324_), .Y(_17__3_) );
INVX1 INVX1_59 ( .A(_17__3_), .Y(_329_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_330_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_331_) );
NAND3X1 NAND3X1_20 ( .A(_329_), .B(_331_), .C(_330_), .Y(_332_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_326_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_327_) );
OAI21X1 OAI21X1_79 ( .A(_326_), .B(_327_), .C(_17__3_), .Y(_328_) );
NAND2X1 NAND2X1_79 ( .A(_328_), .B(_332_), .Y(_15__3_) );
OAI21X1 OAI21X1_80 ( .A(_329_), .B(_326_), .C(_331_), .Y(_13_) );
INVX1 INVX1_60 ( .A(1'b1), .Y(_336_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_337_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_338_) );
NAND3X1 NAND3X1_21 ( .A(_336_), .B(_338_), .C(_337_), .Y(_339_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_333_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_334_) );
OAI21X1 OAI21X1_81 ( .A(_333_), .B(_334_), .C(1'b1), .Y(_335_) );
NAND2X1 NAND2X1_81 ( .A(_335_), .B(_339_), .Y(_16__0_) );
OAI21X1 OAI21X1_82 ( .A(_336_), .B(_333_), .C(_338_), .Y(_18__1_) );
INVX1 INVX1_61 ( .A(_18__1_), .Y(_343_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_344_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_345_) );
NAND3X1 NAND3X1_22 ( .A(_343_), .B(_345_), .C(_344_), .Y(_346_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_340_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_341_) );
OAI21X1 OAI21X1_83 ( .A(_340_), .B(_341_), .C(_18__1_), .Y(_342_) );
NAND2X1 NAND2X1_83 ( .A(_342_), .B(_346_), .Y(_16__1_) );
OAI21X1 OAI21X1_84 ( .A(_343_), .B(_340_), .C(_345_), .Y(_18__2_) );
INVX1 INVX1_62 ( .A(_18__2_), .Y(_350_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_351_) );
NAND2X1 NAND2X1_84 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_352_) );
NAND3X1 NAND3X1_23 ( .A(_350_), .B(_352_), .C(_351_), .Y(_353_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_347_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_348_) );
OAI21X1 OAI21X1_85 ( .A(_347_), .B(_348_), .C(_18__2_), .Y(_349_) );
NAND2X1 NAND2X1_85 ( .A(_349_), .B(_353_), .Y(_16__2_) );
OAI21X1 OAI21X1_86 ( .A(_350_), .B(_347_), .C(_352_), .Y(_18__3_) );
INVX1 INVX1_63 ( .A(_18__3_), .Y(_357_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_358_) );
NAND2X1 NAND2X1_86 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_359_) );
NAND3X1 NAND3X1_24 ( .A(_357_), .B(_359_), .C(_358_), .Y(_360_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_354_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_355_) );
OAI21X1 OAI21X1_87 ( .A(_354_), .B(_355_), .C(_18__3_), .Y(_356_) );
NAND2X1 NAND2X1_87 ( .A(_356_), .B(_360_), .Y(_16__3_) );
OAI21X1 OAI21X1_88 ( .A(_357_), .B(_354_), .C(_359_), .Y(_14_) );
INVX1 INVX1_64 ( .A(1'b0), .Y(_364_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_365_) );
NAND2X1 NAND2X1_88 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_366_) );
NAND3X1 NAND3X1_25 ( .A(_364_), .B(_366_), .C(_365_), .Y(_367_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_361_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_362_) );
OAI21X1 OAI21X1_89 ( .A(_361_), .B(_362_), .C(1'b0), .Y(_363_) );
NAND2X1 NAND2X1_89 ( .A(_363_), .B(_367_), .Y(_21__0_) );
OAI21X1 OAI21X1_90 ( .A(_364_), .B(_361_), .C(_366_), .Y(_23__1_) );
INVX1 INVX1_65 ( .A(_23__1_), .Y(_371_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_372_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_373_) );
NAND3X1 NAND3X1_26 ( .A(_371_), .B(_373_), .C(_372_), .Y(_374_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_368_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_369_) );
OAI21X1 OAI21X1_91 ( .A(_368_), .B(_369_), .C(_23__1_), .Y(_370_) );
NAND2X1 NAND2X1_91 ( .A(_370_), .B(_374_), .Y(_21__1_) );
OAI21X1 OAI21X1_92 ( .A(_371_), .B(_368_), .C(_373_), .Y(_23__2_) );
INVX1 INVX1_66 ( .A(_23__2_), .Y(_378_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_379_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_380_) );
NAND3X1 NAND3X1_27 ( .A(_378_), .B(_380_), .C(_379_), .Y(_381_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_375_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_376_) );
OAI21X1 OAI21X1_93 ( .A(_375_), .B(_376_), .C(_23__2_), .Y(_377_) );
NAND2X1 NAND2X1_93 ( .A(_377_), .B(_381_), .Y(_21__2_) );
OAI21X1 OAI21X1_94 ( .A(_378_), .B(_375_), .C(_380_), .Y(_23__3_) );
INVX1 INVX1_67 ( .A(_23__3_), .Y(_385_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_386_) );
NAND2X1 NAND2X1_94 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_387_) );
NAND3X1 NAND3X1_28 ( .A(_385_), .B(_387_), .C(_386_), .Y(_388_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_382_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_383_) );
OAI21X1 OAI21X1_95 ( .A(_382_), .B(_383_), .C(_23__3_), .Y(_384_) );
NAND2X1 NAND2X1_95 ( .A(_384_), .B(_388_), .Y(_21__3_) );
OAI21X1 OAI21X1_96 ( .A(_385_), .B(_382_), .C(_387_), .Y(_19_) );
INVX1 INVX1_68 ( .A(1'b1), .Y(_392_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_393_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_394_) );
NAND3X1 NAND3X1_29 ( .A(_392_), .B(_394_), .C(_393_), .Y(_395_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_389_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_390_) );
OAI21X1 OAI21X1_97 ( .A(_389_), .B(_390_), .C(1'b1), .Y(_391_) );
NAND2X1 NAND2X1_97 ( .A(_391_), .B(_395_), .Y(_22__0_) );
OAI21X1 OAI21X1_98 ( .A(_392_), .B(_389_), .C(_394_), .Y(_24__1_) );
INVX1 INVX1_69 ( .A(_24__1_), .Y(_399_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_400_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_401_) );
NAND3X1 NAND3X1_30 ( .A(_399_), .B(_401_), .C(_400_), .Y(_402_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_396_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_397_) );
OAI21X1 OAI21X1_99 ( .A(_396_), .B(_397_), .C(_24__1_), .Y(_398_) );
NAND2X1 NAND2X1_99 ( .A(_398_), .B(_402_), .Y(_22__1_) );
OAI21X1 OAI21X1_100 ( .A(_399_), .B(_396_), .C(_401_), .Y(_24__2_) );
INVX1 INVX1_70 ( .A(_24__2_), .Y(_406_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_407_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_408_) );
NAND3X1 NAND3X1_31 ( .A(_406_), .B(_408_), .C(_407_), .Y(_409_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_403_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_404_) );
OAI21X1 OAI21X1_101 ( .A(_403_), .B(_404_), .C(_24__2_), .Y(_405_) );
NAND2X1 NAND2X1_101 ( .A(_405_), .B(_409_), .Y(_22__2_) );
OAI21X1 OAI21X1_102 ( .A(_406_), .B(_403_), .C(_408_), .Y(_24__3_) );
INVX1 INVX1_71 ( .A(_24__3_), .Y(_413_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_414_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_415_) );
NAND3X1 NAND3X1_32 ( .A(_413_), .B(_415_), .C(_414_), .Y(_416_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_410_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_411_) );
OAI21X1 OAI21X1_103 ( .A(_410_), .B(_411_), .C(_24__3_), .Y(_412_) );
NAND2X1 NAND2X1_103 ( .A(_412_), .B(_416_), .Y(_22__3_) );
OAI21X1 OAI21X1_104 ( .A(_413_), .B(_410_), .C(_415_), .Y(_20_) );
INVX1 INVX1_72 ( .A(1'b0), .Y(_420_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_421_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_422_) );
NAND3X1 NAND3X1_33 ( .A(_420_), .B(_422_), .C(_421_), .Y(_423_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_417_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_418_) );
OAI21X1 OAI21X1_105 ( .A(_417_), .B(_418_), .C(1'b0), .Y(_419_) );
NAND2X1 NAND2X1_105 ( .A(_419_), .B(_423_), .Y(_27__0_) );
OAI21X1 OAI21X1_106 ( .A(_420_), .B(_417_), .C(_422_), .Y(_29__1_) );
INVX1 INVX1_73 ( .A(_29__1_), .Y(_427_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_428_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_429_) );
NAND3X1 NAND3X1_34 ( .A(_427_), .B(_429_), .C(_428_), .Y(_430_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_424_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_425_) );
OAI21X1 OAI21X1_107 ( .A(_424_), .B(_425_), .C(_29__1_), .Y(_426_) );
NAND2X1 NAND2X1_107 ( .A(_426_), .B(_430_), .Y(_27__1_) );
OAI21X1 OAI21X1_108 ( .A(_427_), .B(_424_), .C(_429_), .Y(_29__2_) );
INVX1 INVX1_74 ( .A(_29__2_), .Y(_434_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_435_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_436_) );
NAND3X1 NAND3X1_35 ( .A(_434_), .B(_436_), .C(_435_), .Y(_437_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_431_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_432_) );
OAI21X1 OAI21X1_109 ( .A(_431_), .B(_432_), .C(_29__2_), .Y(_433_) );
NAND2X1 NAND2X1_109 ( .A(_433_), .B(_437_), .Y(_27__2_) );
OAI21X1 OAI21X1_110 ( .A(_434_), .B(_431_), .C(_436_), .Y(_29__3_) );
INVX1 INVX1_75 ( .A(_29__3_), .Y(_441_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_442_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_443_) );
NAND3X1 NAND3X1_36 ( .A(_441_), .B(_443_), .C(_442_), .Y(_444_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_438_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_439_) );
OAI21X1 OAI21X1_111 ( .A(_438_), .B(_439_), .C(_29__3_), .Y(_440_) );
NAND2X1 NAND2X1_111 ( .A(_440_), .B(_444_), .Y(_27__3_) );
OAI21X1 OAI21X1_112 ( .A(_441_), .B(_438_), .C(_443_), .Y(_25_) );
INVX1 INVX1_76 ( .A(1'b1), .Y(_448_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_449_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_450_) );
NAND3X1 NAND3X1_37 ( .A(_448_), .B(_450_), .C(_449_), .Y(_451_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_445_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_446_) );
OAI21X1 OAI21X1_113 ( .A(_445_), .B(_446_), .C(1'b1), .Y(_447_) );
NAND2X1 NAND2X1_113 ( .A(_447_), .B(_451_), .Y(_28__0_) );
OAI21X1 OAI21X1_114 ( .A(_448_), .B(_445_), .C(_450_), .Y(_30__1_) );
INVX1 INVX1_77 ( .A(_30__1_), .Y(_455_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_456_) );
NAND2X1 NAND2X1_114 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_457_) );
NAND3X1 NAND3X1_38 ( .A(_455_), .B(_457_), .C(_456_), .Y(_458_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_452_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_453_) );
OAI21X1 OAI21X1_115 ( .A(_452_), .B(_453_), .C(_30__1_), .Y(_454_) );
NAND2X1 NAND2X1_115 ( .A(_454_), .B(_458_), .Y(_28__1_) );
OAI21X1 OAI21X1_116 ( .A(_455_), .B(_452_), .C(_457_), .Y(_30__2_) );
INVX1 INVX1_78 ( .A(_30__2_), .Y(_462_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_463_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_464_) );
NAND3X1 NAND3X1_39 ( .A(_462_), .B(_464_), .C(_463_), .Y(_465_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_459_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_460_) );
OAI21X1 OAI21X1_117 ( .A(_459_), .B(_460_), .C(_30__2_), .Y(_461_) );
NAND2X1 NAND2X1_117 ( .A(_461_), .B(_465_), .Y(_28__2_) );
OAI21X1 OAI21X1_118 ( .A(_462_), .B(_459_), .C(_464_), .Y(_30__3_) );
INVX1 INVX1_79 ( .A(_30__3_), .Y(_469_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_470_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_471_) );
NAND3X1 NAND3X1_40 ( .A(_469_), .B(_471_), .C(_470_), .Y(_472_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_466_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_467_) );
OAI21X1 OAI21X1_119 ( .A(_466_), .B(_467_), .C(_30__3_), .Y(_468_) );
NAND2X1 NAND2X1_119 ( .A(_468_), .B(_472_), .Y(_28__3_) );
OAI21X1 OAI21X1_120 ( .A(_469_), .B(_466_), .C(_471_), .Y(_26_) );
INVX1 INVX1_80 ( .A(1'b0), .Y(_476_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_477_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_478_) );
NAND3X1 NAND3X1_41 ( .A(_476_), .B(_478_), .C(_477_), .Y(_479_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_473_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_474_) );
OAI21X1 OAI21X1_121 ( .A(_473_), .B(_474_), .C(1'b0), .Y(_475_) );
NAND2X1 NAND2X1_121 ( .A(_475_), .B(_479_), .Y(_33__0_) );
OAI21X1 OAI21X1_122 ( .A(_476_), .B(_473_), .C(_478_), .Y(_35__1_) );
INVX1 INVX1_81 ( .A(_35__1_), .Y(_483_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_484_) );
NAND2X1 NAND2X1_122 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_485_) );
NAND3X1 NAND3X1_42 ( .A(_483_), .B(_485_), .C(_484_), .Y(_486_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_480_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_481_) );
OAI21X1 OAI21X1_123 ( .A(_480_), .B(_481_), .C(_35__1_), .Y(_482_) );
NAND2X1 NAND2X1_123 ( .A(_482_), .B(_486_), .Y(_33__1_) );
OAI21X1 OAI21X1_124 ( .A(_483_), .B(_480_), .C(_485_), .Y(_35__2_) );
INVX1 INVX1_82 ( .A(_35__2_), .Y(_490_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_491_) );
NAND2X1 NAND2X1_124 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_492_) );
NAND3X1 NAND3X1_43 ( .A(_490_), .B(_492_), .C(_491_), .Y(_493_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_487_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_488_) );
OAI21X1 OAI21X1_125 ( .A(_487_), .B(_488_), .C(_35__2_), .Y(_489_) );
NAND2X1 NAND2X1_125 ( .A(_489_), .B(_493_), .Y(_33__2_) );
OAI21X1 OAI21X1_126 ( .A(_490_), .B(_487_), .C(_492_), .Y(_35__3_) );
INVX1 INVX1_83 ( .A(_35__3_), .Y(_497_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_498_) );
NAND2X1 NAND2X1_126 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_499_) );
NAND3X1 NAND3X1_44 ( .A(_497_), .B(_499_), .C(_498_), .Y(_500_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_494_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_495_) );
OAI21X1 OAI21X1_127 ( .A(_494_), .B(_495_), .C(_35__3_), .Y(_496_) );
NAND2X1 NAND2X1_127 ( .A(_496_), .B(_500_), .Y(_33__3_) );
OAI21X1 OAI21X1_128 ( .A(_497_), .B(_494_), .C(_499_), .Y(_31_) );
INVX1 INVX1_84 ( .A(1'b1), .Y(_504_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_505_) );
NAND2X1 NAND2X1_128 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_506_) );
NAND3X1 NAND3X1_45 ( .A(_504_), .B(_506_), .C(_505_), .Y(_507_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_501_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_502_) );
OAI21X1 OAI21X1_129 ( .A(_501_), .B(_502_), .C(1'b1), .Y(_503_) );
NAND2X1 NAND2X1_129 ( .A(_503_), .B(_507_), .Y(_34__0_) );
OAI21X1 OAI21X1_130 ( .A(_504_), .B(_501_), .C(_506_), .Y(_36__1_) );
INVX1 INVX1_85 ( .A(_36__1_), .Y(_511_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_512_) );
NAND2X1 NAND2X1_130 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_513_) );
NAND3X1 NAND3X1_46 ( .A(_511_), .B(_513_), .C(_512_), .Y(_514_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_508_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_509_) );
OAI21X1 OAI21X1_131 ( .A(_508_), .B(_509_), .C(_36__1_), .Y(_510_) );
NAND2X1 NAND2X1_131 ( .A(_510_), .B(_514_), .Y(_34__1_) );
OAI21X1 OAI21X1_132 ( .A(_511_), .B(_508_), .C(_513_), .Y(_36__2_) );
INVX1 INVX1_86 ( .A(_36__2_), .Y(_518_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_519_) );
NAND2X1 NAND2X1_132 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_520_) );
NAND3X1 NAND3X1_47 ( .A(_518_), .B(_520_), .C(_519_), .Y(_521_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_515_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_516_) );
OAI21X1 OAI21X1_133 ( .A(_515_), .B(_516_), .C(_36__2_), .Y(_517_) );
NAND2X1 NAND2X1_133 ( .A(_517_), .B(_521_), .Y(_34__2_) );
OAI21X1 OAI21X1_134 ( .A(_518_), .B(_515_), .C(_520_), .Y(_36__3_) );
INVX1 INVX1_87 ( .A(_36__3_), .Y(_525_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_526_) );
NAND2X1 NAND2X1_134 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_527_) );
NAND3X1 NAND3X1_48 ( .A(_525_), .B(_527_), .C(_526_), .Y(_528_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_522_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_523_) );
OAI21X1 OAI21X1_135 ( .A(_522_), .B(_523_), .C(_36__3_), .Y(_524_) );
NAND2X1 NAND2X1_135 ( .A(_524_), .B(_528_), .Y(_34__3_) );
OAI21X1 OAI21X1_136 ( .A(_525_), .B(_522_), .C(_527_), .Y(_32_) );
INVX1 INVX1_88 ( .A(1'b0), .Y(_532_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_533_) );
NAND2X1 NAND2X1_136 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_534_) );
NAND3X1 NAND3X1_49 ( .A(_532_), .B(_534_), .C(_533_), .Y(_535_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_529_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_530_) );
OAI21X1 OAI21X1_137 ( .A(_529_), .B(_530_), .C(1'b0), .Y(_531_) );
NAND2X1 NAND2X1_137 ( .A(_531_), .B(_535_), .Y(_39__0_) );
OAI21X1 OAI21X1_138 ( .A(_532_), .B(_529_), .C(_534_), .Y(_41__1_) );
INVX1 INVX1_89 ( .A(_41__1_), .Y(_539_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_540_) );
NAND2X1 NAND2X1_138 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_541_) );
NAND3X1 NAND3X1_50 ( .A(_539_), .B(_541_), .C(_540_), .Y(_542_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_536_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_537_) );
OAI21X1 OAI21X1_139 ( .A(_536_), .B(_537_), .C(_41__1_), .Y(_538_) );
NAND2X1 NAND2X1_139 ( .A(_538_), .B(_542_), .Y(_39__1_) );
OAI21X1 OAI21X1_140 ( .A(_539_), .B(_536_), .C(_541_), .Y(_41__2_) );
INVX1 INVX1_90 ( .A(_41__2_), .Y(_546_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_547_) );
NAND2X1 NAND2X1_140 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_548_) );
NAND3X1 NAND3X1_51 ( .A(_546_), .B(_548_), .C(_547_), .Y(_549_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_543_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_544_) );
OAI21X1 OAI21X1_141 ( .A(_543_), .B(_544_), .C(_41__2_), .Y(_545_) );
NAND2X1 NAND2X1_141 ( .A(_545_), .B(_549_), .Y(_39__2_) );
OAI21X1 OAI21X1_142 ( .A(_546_), .B(_543_), .C(_548_), .Y(_41__3_) );
INVX1 INVX1_91 ( .A(_41__3_), .Y(_553_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_554_) );
NAND2X1 NAND2X1_142 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_555_) );
NAND3X1 NAND3X1_52 ( .A(_553_), .B(_555_), .C(_554_), .Y(_556_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_550_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_551_) );
OAI21X1 OAI21X1_143 ( .A(_550_), .B(_551_), .C(_41__3_), .Y(_552_) );
NAND2X1 NAND2X1_143 ( .A(_552_), .B(_556_), .Y(_39__3_) );
OAI21X1 OAI21X1_144 ( .A(_553_), .B(_550_), .C(_555_), .Y(_37_) );
INVX1 INVX1_92 ( .A(1'b1), .Y(_560_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_561_) );
NAND2X1 NAND2X1_144 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_562_) );
NAND3X1 NAND3X1_53 ( .A(_560_), .B(_562_), .C(_561_), .Y(_563_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_557_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_558_) );
OAI21X1 OAI21X1_145 ( .A(_557_), .B(_558_), .C(1'b1), .Y(_559_) );
NAND2X1 NAND2X1_145 ( .A(_559_), .B(_563_), .Y(_40__0_) );
OAI21X1 OAI21X1_146 ( .A(_560_), .B(_557_), .C(_562_), .Y(_42__1_) );
INVX1 INVX1_93 ( .A(_42__1_), .Y(_567_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_568_) );
NAND2X1 NAND2X1_146 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_569_) );
NAND3X1 NAND3X1_54 ( .A(_567_), .B(_569_), .C(_568_), .Y(_570_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_564_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_565_) );
OAI21X1 OAI21X1_147 ( .A(_564_), .B(_565_), .C(_42__1_), .Y(_566_) );
NAND2X1 NAND2X1_147 ( .A(_566_), .B(_570_), .Y(_40__1_) );
OAI21X1 OAI21X1_148 ( .A(_567_), .B(_564_), .C(_569_), .Y(_42__2_) );
INVX1 INVX1_94 ( .A(_42__2_), .Y(_574_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_575_) );
NAND2X1 NAND2X1_148 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_576_) );
NAND3X1 NAND3X1_55 ( .A(_574_), .B(_576_), .C(_575_), .Y(_577_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_571_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_572_) );
OAI21X1 OAI21X1_149 ( .A(_571_), .B(_572_), .C(_42__2_), .Y(_573_) );
NAND2X1 NAND2X1_149 ( .A(_573_), .B(_577_), .Y(_40__2_) );
OAI21X1 OAI21X1_150 ( .A(_574_), .B(_571_), .C(_576_), .Y(_42__3_) );
INVX1 INVX1_95 ( .A(_42__3_), .Y(_581_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_582_) );
NAND2X1 NAND2X1_150 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_583_) );
NAND3X1 NAND3X1_56 ( .A(_581_), .B(_583_), .C(_582_), .Y(_584_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_578_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_579_) );
OAI21X1 OAI21X1_151 ( .A(_578_), .B(_579_), .C(_42__3_), .Y(_580_) );
NAND2X1 NAND2X1_151 ( .A(_580_), .B(_584_), .Y(_40__3_) );
OAI21X1 OAI21X1_152 ( .A(_581_), .B(_578_), .C(_583_), .Y(_38_) );
INVX1 INVX1_96 ( .A(1'b0), .Y(_588_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_589_) );
NAND2X1 NAND2X1_152 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_590_) );
NAND3X1 NAND3X1_57 ( .A(_588_), .B(_590_), .C(_589_), .Y(_591_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_585_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_586_) );
OAI21X1 OAI21X1_153 ( .A(_585_), .B(_586_), .C(1'b0), .Y(_587_) );
NAND2X1 NAND2X1_153 ( .A(_587_), .B(_591_), .Y(_45__0_) );
OAI21X1 OAI21X1_154 ( .A(_588_), .B(_585_), .C(_590_), .Y(_47__1_) );
INVX1 INVX1_97 ( .A(_47__1_), .Y(_595_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_596_) );
NAND2X1 NAND2X1_154 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_597_) );
NAND3X1 NAND3X1_58 ( .A(_595_), .B(_597_), .C(_596_), .Y(_598_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_592_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_593_) );
OAI21X1 OAI21X1_155 ( .A(_592_), .B(_593_), .C(_47__1_), .Y(_594_) );
NAND2X1 NAND2X1_155 ( .A(_594_), .B(_598_), .Y(_45__1_) );
OAI21X1 OAI21X1_156 ( .A(_595_), .B(_592_), .C(_597_), .Y(_47__2_) );
INVX1 INVX1_98 ( .A(_47__2_), .Y(_602_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_603_) );
NAND2X1 NAND2X1_156 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_604_) );
NAND3X1 NAND3X1_59 ( .A(_602_), .B(_604_), .C(_603_), .Y(_605_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_599_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_600_) );
OAI21X1 OAI21X1_157 ( .A(_599_), .B(_600_), .C(_47__2_), .Y(_601_) );
NAND2X1 NAND2X1_157 ( .A(_601_), .B(_605_), .Y(_45__2_) );
OAI21X1 OAI21X1_158 ( .A(_602_), .B(_599_), .C(_604_), .Y(_47__3_) );
INVX1 INVX1_99 ( .A(_47__3_), .Y(_609_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_610_) );
NAND2X1 NAND2X1_158 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_611_) );
NAND3X1 NAND3X1_60 ( .A(_609_), .B(_611_), .C(_610_), .Y(_612_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_606_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_607_) );
OAI21X1 OAI21X1_159 ( .A(_606_), .B(_607_), .C(_47__3_), .Y(_608_) );
NAND2X1 NAND2X1_159 ( .A(_608_), .B(_612_), .Y(_45__3_) );
OAI21X1 OAI21X1_160 ( .A(_609_), .B(_606_), .C(_611_), .Y(_43_) );
INVX1 INVX1_100 ( .A(1'b1), .Y(_616_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_617_) );
NAND2X1 NAND2X1_160 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_618_) );
NAND3X1 NAND3X1_61 ( .A(_616_), .B(_618_), .C(_617_), .Y(_619_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_613_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_614_) );
OAI21X1 OAI21X1_161 ( .A(_613_), .B(_614_), .C(1'b1), .Y(_615_) );
NAND2X1 NAND2X1_161 ( .A(_615_), .B(_619_), .Y(_46__0_) );
OAI21X1 OAI21X1_162 ( .A(_616_), .B(_613_), .C(_618_), .Y(_48__1_) );
INVX1 INVX1_101 ( .A(_48__1_), .Y(_623_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_624_) );
NAND2X1 NAND2X1_162 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_625_) );
NAND3X1 NAND3X1_62 ( .A(_623_), .B(_625_), .C(_624_), .Y(_626_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_620_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_621_) );
OAI21X1 OAI21X1_163 ( .A(_620_), .B(_621_), .C(_48__1_), .Y(_622_) );
NAND2X1 NAND2X1_163 ( .A(_622_), .B(_626_), .Y(_46__1_) );
OAI21X1 OAI21X1_164 ( .A(_623_), .B(_620_), .C(_625_), .Y(_48__2_) );
INVX1 INVX1_102 ( .A(_48__2_), .Y(_630_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_631_) );
NAND2X1 NAND2X1_164 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_632_) );
NAND3X1 NAND3X1_63 ( .A(_630_), .B(_632_), .C(_631_), .Y(_633_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_627_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_628_) );
OAI21X1 OAI21X1_165 ( .A(_627_), .B(_628_), .C(_48__2_), .Y(_629_) );
NAND2X1 NAND2X1_165 ( .A(_629_), .B(_633_), .Y(_46__2_) );
OAI21X1 OAI21X1_166 ( .A(_630_), .B(_627_), .C(_632_), .Y(_48__3_) );
INVX1 INVX1_103 ( .A(_48__3_), .Y(_637_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_638_) );
NAND2X1 NAND2X1_166 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_639_) );
NAND3X1 NAND3X1_64 ( .A(_637_), .B(_639_), .C(_638_), .Y(_640_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_634_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_635_) );
OAI21X1 OAI21X1_167 ( .A(_634_), .B(_635_), .C(_48__3_), .Y(_636_) );
NAND2X1 NAND2X1_167 ( .A(_636_), .B(_640_), .Y(_46__3_) );
OAI21X1 OAI21X1_168 ( .A(_637_), .B(_634_), .C(_639_), .Y(_44_) );
INVX1 INVX1_104 ( .A(1'b0), .Y(_644_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_645_) );
NAND2X1 NAND2X1_168 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_646_) );
NAND3X1 NAND3X1_65 ( .A(_644_), .B(_646_), .C(_645_), .Y(_647_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_641_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_642_) );
OAI21X1 OAI21X1_169 ( .A(_641_), .B(_642_), .C(1'b0), .Y(_643_) );
NAND2X1 NAND2X1_169 ( .A(_643_), .B(_647_), .Y(_51__0_) );
OAI21X1 OAI21X1_170 ( .A(_644_), .B(_641_), .C(_646_), .Y(_53__1_) );
INVX1 INVX1_105 ( .A(_53__1_), .Y(_651_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_652_) );
NAND2X1 NAND2X1_170 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_653_) );
NAND3X1 NAND3X1_66 ( .A(_651_), .B(_653_), .C(_652_), .Y(_654_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_648_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_649_) );
OAI21X1 OAI21X1_171 ( .A(_648_), .B(_649_), .C(_53__1_), .Y(_650_) );
NAND2X1 NAND2X1_171 ( .A(_650_), .B(_654_), .Y(_51__1_) );
OAI21X1 OAI21X1_172 ( .A(_651_), .B(_648_), .C(_653_), .Y(_53__2_) );
INVX1 INVX1_106 ( .A(_53__2_), .Y(_658_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_659_) );
NAND2X1 NAND2X1_172 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_660_) );
NAND3X1 NAND3X1_67 ( .A(_658_), .B(_660_), .C(_659_), .Y(_661_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_655_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_656_) );
OAI21X1 OAI21X1_173 ( .A(_655_), .B(_656_), .C(_53__2_), .Y(_657_) );
NAND2X1 NAND2X1_173 ( .A(_657_), .B(_661_), .Y(_51__2_) );
OAI21X1 OAI21X1_174 ( .A(_658_), .B(_655_), .C(_660_), .Y(_53__3_) );
INVX1 INVX1_107 ( .A(_53__3_), .Y(_665_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_666_) );
NAND2X1 NAND2X1_174 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_667_) );
NAND3X1 NAND3X1_68 ( .A(_665_), .B(_667_), .C(_666_), .Y(_668_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_662_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_663_) );
OAI21X1 OAI21X1_175 ( .A(_662_), .B(_663_), .C(_53__3_), .Y(_664_) );
NAND2X1 NAND2X1_175 ( .A(_664_), .B(_668_), .Y(_51__3_) );
OAI21X1 OAI21X1_176 ( .A(_665_), .B(_662_), .C(_667_), .Y(_49_) );
INVX1 INVX1_108 ( .A(1'b1), .Y(_672_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_673_) );
NAND2X1 NAND2X1_176 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_674_) );
NAND3X1 NAND3X1_69 ( .A(_672_), .B(_674_), .C(_673_), .Y(_675_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_669_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_670_) );
OAI21X1 OAI21X1_177 ( .A(_669_), .B(_670_), .C(1'b1), .Y(_671_) );
NAND2X1 NAND2X1_177 ( .A(_671_), .B(_675_), .Y(_52__0_) );
OAI21X1 OAI21X1_178 ( .A(_672_), .B(_669_), .C(_674_), .Y(_54__1_) );
INVX1 INVX1_109 ( .A(_54__1_), .Y(_679_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_680_) );
NAND2X1 NAND2X1_178 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_681_) );
NAND3X1 NAND3X1_70 ( .A(_679_), .B(_681_), .C(_680_), .Y(_682_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_676_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_677_) );
OAI21X1 OAI21X1_179 ( .A(_676_), .B(_677_), .C(_54__1_), .Y(_678_) );
NAND2X1 NAND2X1_179 ( .A(_678_), .B(_682_), .Y(_52__1_) );
OAI21X1 OAI21X1_180 ( .A(_679_), .B(_676_), .C(_681_), .Y(_54__2_) );
INVX1 INVX1_110 ( .A(_54__2_), .Y(_686_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_687_) );
NAND2X1 NAND2X1_180 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_688_) );
NAND3X1 NAND3X1_71 ( .A(_686_), .B(_688_), .C(_687_), .Y(_689_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_683_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_684_) );
OAI21X1 OAI21X1_181 ( .A(_683_), .B(_684_), .C(_54__2_), .Y(_685_) );
NAND2X1 NAND2X1_181 ( .A(_685_), .B(_689_), .Y(_52__2_) );
OAI21X1 OAI21X1_182 ( .A(_686_), .B(_683_), .C(_688_), .Y(_54__3_) );
INVX1 INVX1_111 ( .A(_54__3_), .Y(_693_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_694_) );
NAND2X1 NAND2X1_182 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_695_) );
NAND3X1 NAND3X1_72 ( .A(_693_), .B(_695_), .C(_694_), .Y(_696_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_690_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_691_) );
OAI21X1 OAI21X1_183 ( .A(_690_), .B(_691_), .C(_54__3_), .Y(_692_) );
NAND2X1 NAND2X1_183 ( .A(_692_), .B(_696_), .Y(_52__3_) );
OAI21X1 OAI21X1_184 ( .A(_693_), .B(_690_), .C(_695_), .Y(_50_) );
INVX1 INVX1_112 ( .A(1'b0), .Y(_700_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_701_) );
NAND2X1 NAND2X1_184 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_702_) );
NAND3X1 NAND3X1_73 ( .A(_700_), .B(_702_), .C(_701_), .Y(_703_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_697_) );
AND2X2 AND2X2_73 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_698_) );
OAI21X1 OAI21X1_185 ( .A(_697_), .B(_698_), .C(1'b0), .Y(_699_) );
NAND2X1 NAND2X1_185 ( .A(_699_), .B(_703_), .Y(_57__0_) );
OAI21X1 OAI21X1_186 ( .A(_700_), .B(_697_), .C(_702_), .Y(_59__1_) );
INVX1 INVX1_113 ( .A(_59__1_), .Y(_707_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_708_) );
NAND2X1 NAND2X1_186 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_709_) );
NAND3X1 NAND3X1_74 ( .A(_707_), .B(_709_), .C(_708_), .Y(_710_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_704_) );
AND2X2 AND2X2_74 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_705_) );
OAI21X1 OAI21X1_187 ( .A(_704_), .B(_705_), .C(_59__1_), .Y(_706_) );
NAND2X1 NAND2X1_187 ( .A(_706_), .B(_710_), .Y(_57__1_) );
OAI21X1 OAI21X1_188 ( .A(_707_), .B(_704_), .C(_709_), .Y(_59__2_) );
INVX1 INVX1_114 ( .A(_59__2_), .Y(_714_) );
OR2X2 OR2X2_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_715_) );
NAND2X1 NAND2X1_188 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_716_) );
NAND3X1 NAND3X1_75 ( .A(_714_), .B(_716_), .C(_715_), .Y(_717_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_711_) );
AND2X2 AND2X2_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_712_) );
OAI21X1 OAI21X1_189 ( .A(_711_), .B(_712_), .C(_59__2_), .Y(_713_) );
NAND2X1 NAND2X1_189 ( .A(_713_), .B(_717_), .Y(_57__2_) );
OAI21X1 OAI21X1_190 ( .A(_714_), .B(_711_), .C(_716_), .Y(_59__3_) );
INVX1 INVX1_115 ( .A(_59__3_), .Y(_721_) );
OR2X2 OR2X2_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_722_) );
NAND2X1 NAND2X1_190 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_723_) );
NAND3X1 NAND3X1_76 ( .A(_721_), .B(_723_), .C(_722_), .Y(_724_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_718_) );
AND2X2 AND2X2_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_719_) );
OAI21X1 OAI21X1_191 ( .A(_718_), .B(_719_), .C(_59__3_), .Y(_720_) );
NAND2X1 NAND2X1_191 ( .A(_720_), .B(_724_), .Y(_57__3_) );
OAI21X1 OAI21X1_192 ( .A(_721_), .B(_718_), .C(_723_), .Y(_55_) );
INVX1 INVX1_116 ( .A(1'b1), .Y(_728_) );
OR2X2 OR2X2_77 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_729_) );
NAND2X1 NAND2X1_192 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_730_) );
NAND3X1 NAND3X1_77 ( .A(_728_), .B(_730_), .C(_729_), .Y(_731_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_725_) );
AND2X2 AND2X2_77 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_726_) );
OAI21X1 OAI21X1_193 ( .A(_725_), .B(_726_), .C(1'b1), .Y(_727_) );
NAND2X1 NAND2X1_193 ( .A(_727_), .B(_731_), .Y(_58__0_) );
OAI21X1 OAI21X1_194 ( .A(_728_), .B(_725_), .C(_730_), .Y(_60__1_) );
INVX1 INVX1_117 ( .A(_60__1_), .Y(_735_) );
OR2X2 OR2X2_78 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_736_) );
NAND2X1 NAND2X1_194 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_737_) );
NAND3X1 NAND3X1_78 ( .A(_735_), .B(_737_), .C(_736_), .Y(_738_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_732_) );
AND2X2 AND2X2_78 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_733_) );
OAI21X1 OAI21X1_195 ( .A(_732_), .B(_733_), .C(_60__1_), .Y(_734_) );
NAND2X1 NAND2X1_195 ( .A(_734_), .B(_738_), .Y(_58__1_) );
OAI21X1 OAI21X1_196 ( .A(_735_), .B(_732_), .C(_737_), .Y(_60__2_) );
INVX1 INVX1_118 ( .A(_60__2_), .Y(_742_) );
OR2X2 OR2X2_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_743_) );
NAND2X1 NAND2X1_196 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_744_) );
NAND3X1 NAND3X1_79 ( .A(_742_), .B(_744_), .C(_743_), .Y(_745_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_739_) );
AND2X2 AND2X2_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_740_) );
OAI21X1 OAI21X1_197 ( .A(_739_), .B(_740_), .C(_60__2_), .Y(_741_) );
NAND2X1 NAND2X1_197 ( .A(_741_), .B(_745_), .Y(_58__2_) );
OAI21X1 OAI21X1_198 ( .A(_742_), .B(_739_), .C(_744_), .Y(_60__3_) );
INVX1 INVX1_119 ( .A(_60__3_), .Y(_749_) );
OR2X2 OR2X2_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_750_) );
NAND2X1 NAND2X1_198 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_751_) );
NAND3X1 NAND3X1_80 ( .A(_749_), .B(_751_), .C(_750_), .Y(_752_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_746_) );
AND2X2 AND2X2_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_747_) );
OAI21X1 OAI21X1_199 ( .A(_746_), .B(_747_), .C(_60__3_), .Y(_748_) );
NAND2X1 NAND2X1_199 ( .A(_748_), .B(_752_), .Y(_58__3_) );
OAI21X1 OAI21X1_200 ( .A(_749_), .B(_746_), .C(_751_), .Y(_56_) );
INVX1 INVX1_120 ( .A(1'b0), .Y(_756_) );
OR2X2 OR2X2_81 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_757_) );
NAND2X1 NAND2X1_200 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_758_) );
NAND3X1 NAND3X1_81 ( .A(_756_), .B(_758_), .C(_757_), .Y(_759_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_753_) );
AND2X2 AND2X2_81 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_754_) );
OAI21X1 OAI21X1_201 ( .A(_753_), .B(_754_), .C(1'b0), .Y(_755_) );
NAND2X1 NAND2X1_201 ( .A(_755_), .B(_759_), .Y(_63__0_) );
OAI21X1 OAI21X1_202 ( .A(_756_), .B(_753_), .C(_758_), .Y(_65__1_) );
INVX1 INVX1_121 ( .A(_65__1_), .Y(_763_) );
OR2X2 OR2X2_82 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_764_) );
NAND2X1 NAND2X1_202 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_765_) );
NAND3X1 NAND3X1_82 ( .A(_763_), .B(_765_), .C(_764_), .Y(_766_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_760_) );
AND2X2 AND2X2_82 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_761_) );
OAI21X1 OAI21X1_203 ( .A(_760_), .B(_761_), .C(_65__1_), .Y(_762_) );
NAND2X1 NAND2X1_203 ( .A(_762_), .B(_766_), .Y(_63__1_) );
OAI21X1 OAI21X1_204 ( .A(_763_), .B(_760_), .C(_765_), .Y(_65__2_) );
INVX1 INVX1_122 ( .A(_65__2_), .Y(_770_) );
OR2X2 OR2X2_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_771_) );
NAND2X1 NAND2X1_204 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_772_) );
NAND3X1 NAND3X1_83 ( .A(_770_), .B(_772_), .C(_771_), .Y(_773_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_767_) );
AND2X2 AND2X2_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_768_) );
OAI21X1 OAI21X1_205 ( .A(_767_), .B(_768_), .C(_65__2_), .Y(_769_) );
NAND2X1 NAND2X1_205 ( .A(_769_), .B(_773_), .Y(_63__2_) );
OAI21X1 OAI21X1_206 ( .A(_770_), .B(_767_), .C(_772_), .Y(_65__3_) );
INVX1 INVX1_123 ( .A(_65__3_), .Y(_777_) );
OR2X2 OR2X2_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_778_) );
NAND2X1 NAND2X1_206 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_779_) );
NAND3X1 NAND3X1_84 ( .A(_777_), .B(_779_), .C(_778_), .Y(_780_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_774_) );
AND2X2 AND2X2_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_775_) );
OAI21X1 OAI21X1_207 ( .A(_774_), .B(_775_), .C(_65__3_), .Y(_776_) );
NAND2X1 NAND2X1_207 ( .A(_776_), .B(_780_), .Y(_63__3_) );
OAI21X1 OAI21X1_208 ( .A(_777_), .B(_774_), .C(_779_), .Y(_61_) );
INVX1 INVX1_124 ( .A(1'b1), .Y(_784_) );
OR2X2 OR2X2_85 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_785_) );
NAND2X1 NAND2X1_208 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_786_) );
NAND3X1 NAND3X1_85 ( .A(_784_), .B(_786_), .C(_785_), .Y(_787_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_781_) );
AND2X2 AND2X2_85 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_782_) );
OAI21X1 OAI21X1_209 ( .A(_781_), .B(_782_), .C(1'b1), .Y(_783_) );
NAND2X1 NAND2X1_209 ( .A(_783_), .B(_787_), .Y(_64__0_) );
OAI21X1 OAI21X1_210 ( .A(_784_), .B(_781_), .C(_786_), .Y(_66__1_) );
INVX1 INVX1_125 ( .A(_66__1_), .Y(_791_) );
OR2X2 OR2X2_86 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_792_) );
NAND2X1 NAND2X1_210 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_793_) );
NAND3X1 NAND3X1_86 ( .A(_791_), .B(_793_), .C(_792_), .Y(_794_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_788_) );
AND2X2 AND2X2_86 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_789_) );
OAI21X1 OAI21X1_211 ( .A(_788_), .B(_789_), .C(_66__1_), .Y(_790_) );
NAND2X1 NAND2X1_211 ( .A(_790_), .B(_794_), .Y(_64__1_) );
OAI21X1 OAI21X1_212 ( .A(_791_), .B(_788_), .C(_793_), .Y(_66__2_) );
INVX1 INVX1_126 ( .A(_66__2_), .Y(_798_) );
OR2X2 OR2X2_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_799_) );
NAND2X1 NAND2X1_212 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_800_) );
NAND3X1 NAND3X1_87 ( .A(_798_), .B(_800_), .C(_799_), .Y(_801_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_795_) );
AND2X2 AND2X2_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_796_) );
OAI21X1 OAI21X1_213 ( .A(_795_), .B(_796_), .C(_66__2_), .Y(_797_) );
NAND2X1 NAND2X1_213 ( .A(_797_), .B(_801_), .Y(_64__2_) );
OAI21X1 OAI21X1_214 ( .A(_798_), .B(_795_), .C(_800_), .Y(_66__3_) );
INVX1 INVX1_127 ( .A(_66__3_), .Y(_805_) );
OR2X2 OR2X2_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_806_) );
NAND2X1 NAND2X1_214 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_807_) );
NAND3X1 NAND3X1_88 ( .A(_805_), .B(_807_), .C(_806_), .Y(_808_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_802_) );
AND2X2 AND2X2_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_803_) );
OAI21X1 OAI21X1_215 ( .A(_802_), .B(_803_), .C(_66__3_), .Y(_804_) );
NAND2X1 NAND2X1_215 ( .A(_804_), .B(_808_), .Y(_64__3_) );
OAI21X1 OAI21X1_216 ( .A(_805_), .B(_802_), .C(_807_), .Y(_62_) );
INVX1 INVX1_128 ( .A(1'b0), .Y(_812_) );
OR2X2 OR2X2_89 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_813_) );
NAND2X1 NAND2X1_216 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_814_) );
NAND3X1 NAND3X1_89 ( .A(_812_), .B(_814_), .C(_813_), .Y(_815_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_809_) );
AND2X2 AND2X2_89 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_810_) );
OAI21X1 OAI21X1_217 ( .A(_809_), .B(_810_), .C(1'b0), .Y(_811_) );
NAND2X1 NAND2X1_217 ( .A(_811_), .B(_815_), .Y(_69__0_) );
OAI21X1 OAI21X1_218 ( .A(_812_), .B(_809_), .C(_814_), .Y(_71__1_) );
INVX1 INVX1_129 ( .A(_71__1_), .Y(_819_) );
OR2X2 OR2X2_90 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_820_) );
NAND2X1 NAND2X1_218 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_821_) );
NAND3X1 NAND3X1_90 ( .A(_819_), .B(_821_), .C(_820_), .Y(_822_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_816_) );
AND2X2 AND2X2_90 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_817_) );
OAI21X1 OAI21X1_219 ( .A(_816_), .B(_817_), .C(_71__1_), .Y(_818_) );
NAND2X1 NAND2X1_219 ( .A(_818_), .B(_822_), .Y(_69__1_) );
OAI21X1 OAI21X1_220 ( .A(_819_), .B(_816_), .C(_821_), .Y(_71__2_) );
INVX1 INVX1_130 ( .A(_71__2_), .Y(_826_) );
OR2X2 OR2X2_91 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_827_) );
NAND2X1 NAND2X1_220 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_828_) );
NAND3X1 NAND3X1_91 ( .A(_826_), .B(_828_), .C(_827_), .Y(_829_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_823_) );
AND2X2 AND2X2_91 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_824_) );
OAI21X1 OAI21X1_221 ( .A(_823_), .B(_824_), .C(_71__2_), .Y(_825_) );
NAND2X1 NAND2X1_221 ( .A(_825_), .B(_829_), .Y(_69__2_) );
OAI21X1 OAI21X1_222 ( .A(_826_), .B(_823_), .C(_828_), .Y(_71__3_) );
INVX1 INVX1_131 ( .A(_71__3_), .Y(_833_) );
OR2X2 OR2X2_92 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_834_) );
NAND2X1 NAND2X1_222 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_835_) );
NAND3X1 NAND3X1_92 ( .A(_833_), .B(_835_), .C(_834_), .Y(_836_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_830_) );
AND2X2 AND2X2_92 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_831_) );
OAI21X1 OAI21X1_223 ( .A(_830_), .B(_831_), .C(_71__3_), .Y(_832_) );
NAND2X1 NAND2X1_223 ( .A(_832_), .B(_836_), .Y(_69__3_) );
OAI21X1 OAI21X1_224 ( .A(_833_), .B(_830_), .C(_835_), .Y(_67_) );
INVX1 INVX1_132 ( .A(1'b1), .Y(_840_) );
OR2X2 OR2X2_93 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_841_) );
NAND2X1 NAND2X1_224 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_842_) );
NAND3X1 NAND3X1_93 ( .A(_840_), .B(_842_), .C(_841_), .Y(_843_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_837_) );
AND2X2 AND2X2_93 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_838_) );
OAI21X1 OAI21X1_225 ( .A(_837_), .B(_838_), .C(1'b1), .Y(_839_) );
NAND2X1 NAND2X1_225 ( .A(_839_), .B(_843_), .Y(_70__0_) );
OAI21X1 OAI21X1_226 ( .A(_840_), .B(_837_), .C(_842_), .Y(_72__1_) );
INVX1 INVX1_133 ( .A(_72__1_), .Y(_847_) );
OR2X2 OR2X2_94 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_848_) );
NAND2X1 NAND2X1_226 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_849_) );
NAND3X1 NAND3X1_94 ( .A(_847_), .B(_849_), .C(_848_), .Y(_850_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_844_) );
AND2X2 AND2X2_94 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_845_) );
OAI21X1 OAI21X1_227 ( .A(_844_), .B(_845_), .C(_72__1_), .Y(_846_) );
NAND2X1 NAND2X1_227 ( .A(_846_), .B(_850_), .Y(_70__1_) );
OAI21X1 OAI21X1_228 ( .A(_847_), .B(_844_), .C(_849_), .Y(_72__2_) );
INVX1 INVX1_134 ( .A(_72__2_), .Y(_854_) );
OR2X2 OR2X2_95 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_855_) );
NAND2X1 NAND2X1_228 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_856_) );
NAND3X1 NAND3X1_95 ( .A(_854_), .B(_856_), .C(_855_), .Y(_857_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_851_) );
AND2X2 AND2X2_95 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_852_) );
OAI21X1 OAI21X1_229 ( .A(_851_), .B(_852_), .C(_72__2_), .Y(_853_) );
NAND2X1 NAND2X1_229 ( .A(_853_), .B(_857_), .Y(_70__2_) );
OAI21X1 OAI21X1_230 ( .A(_854_), .B(_851_), .C(_856_), .Y(_72__3_) );
INVX1 INVX1_135 ( .A(_72__3_), .Y(_861_) );
OR2X2 OR2X2_96 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_862_) );
NAND2X1 NAND2X1_230 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_863_) );
NAND3X1 NAND3X1_96 ( .A(_861_), .B(_863_), .C(_862_), .Y(_864_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_858_) );
AND2X2 AND2X2_96 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_859_) );
OAI21X1 OAI21X1_231 ( .A(_858_), .B(_859_), .C(_72__3_), .Y(_860_) );
NAND2X1 NAND2X1_231 ( .A(_860_), .B(_864_), .Y(_70__3_) );
OAI21X1 OAI21X1_232 ( .A(_861_), .B(_858_), .C(_863_), .Y(_68_) );
INVX1 INVX1_136 ( .A(1'b0), .Y(_868_) );
OR2X2 OR2X2_97 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_869_) );
NAND2X1 NAND2X1_232 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_870_) );
NAND3X1 NAND3X1_97 ( .A(_868_), .B(_870_), .C(_869_), .Y(_871_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_865_) );
AND2X2 AND2X2_97 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_866_) );
OAI21X1 OAI21X1_233 ( .A(_865_), .B(_866_), .C(1'b0), .Y(_867_) );
NAND2X1 NAND2X1_233 ( .A(_867_), .B(_871_), .Y(_0__0_) );
OAI21X1 OAI21X1_234 ( .A(_868_), .B(_865_), .C(_870_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_137 ( .A(rca_inst_w_CARRY_1_), .Y(_875_) );
OR2X2 OR2X2_98 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_876_) );
NAND2X1 NAND2X1_234 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_877_) );
NAND3X1 NAND3X1_98 ( .A(_875_), .B(_877_), .C(_876_), .Y(_878_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_872_) );
AND2X2 AND2X2_98 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_873_) );
OAI21X1 OAI21X1_235 ( .A(_872_), .B(_873_), .C(rca_inst_w_CARRY_1_), .Y(_874_) );
NAND2X1 NAND2X1_235 ( .A(_874_), .B(_878_), .Y(_0__1_) );
OAI21X1 OAI21X1_236 ( .A(_875_), .B(_872_), .C(_877_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_138 ( .A(rca_inst_w_CARRY_2_), .Y(_882_) );
OR2X2 OR2X2_99 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_883_) );
NAND2X1 NAND2X1_236 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_884_) );
NAND3X1 NAND3X1_99 ( .A(_882_), .B(_884_), .C(_883_), .Y(_885_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_879_) );
AND2X2 AND2X2_99 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_880_) );
OAI21X1 OAI21X1_237 ( .A(_879_), .B(_880_), .C(rca_inst_w_CARRY_2_), .Y(_881_) );
NAND2X1 NAND2X1_237 ( .A(_881_), .B(_885_), .Y(_0__2_) );
BUFX2 BUFX2_1 ( .A(w_cout_12_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
INVX1 INVX1_139 ( .A(_1_), .Y(_73_) );
NAND2X1 NAND2X1_238 ( .A(_2_), .B(1'b0), .Y(_74_) );
OAI21X1 OAI21X1_238 ( .A(1'b0), .B(_73_), .C(_74_), .Y(w_cout_1_) );
INVX1 INVX1_140 ( .A(_3__0_), .Y(_75_) );
NAND2X1 NAND2X1_239 ( .A(_4__0_), .B(1'b0), .Y(_76_) );
OAI21X1 OAI21X1_239 ( .A(1'b0), .B(_75_), .C(_76_), .Y(_0__3_) );
INVX1 INVX1_141 ( .A(_3__1_), .Y(_77_) );
NAND2X1 NAND2X1_240 ( .A(1'b0), .B(_4__1_), .Y(_78_) );
OAI21X1 OAI21X1_240 ( .A(1'b0), .B(_77_), .C(_78_), .Y(_0__4_) );
INVX1 INVX1_142 ( .A(_3__2_), .Y(_79_) );
NAND2X1 NAND2X1_241 ( .A(1'b0), .B(_4__2_), .Y(_80_) );
OAI21X1 OAI21X1_241 ( .A(1'b0), .B(_79_), .C(_80_), .Y(_0__5_) );
INVX1 INVX1_143 ( .A(_3__3_), .Y(_81_) );
NAND2X1 NAND2X1_242 ( .A(1'b0), .B(_4__3_), .Y(_82_) );
OAI21X1 OAI21X1_242 ( .A(1'b0), .B(_81_), .C(_82_), .Y(_0__6_) );
INVX1 INVX1_144 ( .A(_7_), .Y(_83_) );
NAND2X1 NAND2X1_243 ( .A(_8_), .B(w_cout_1_), .Y(_84_) );
OAI21X1 OAI21X1_243 ( .A(w_cout_1_), .B(_83_), .C(_84_), .Y(w_cout_2_) );
INVX1 INVX1_145 ( .A(_9__0_), .Y(_85_) );
NAND2X1 NAND2X1_244 ( .A(_10__0_), .B(w_cout_1_), .Y(_86_) );
OAI21X1 OAI21X1_244 ( .A(w_cout_1_), .B(_85_), .C(_86_), .Y(_0__7_) );
INVX1 INVX1_146 ( .A(_9__1_), .Y(_87_) );
NAND2X1 NAND2X1_245 ( .A(w_cout_1_), .B(_10__1_), .Y(_88_) );
OAI21X1 OAI21X1_245 ( .A(w_cout_1_), .B(_87_), .C(_88_), .Y(_0__8_) );
INVX1 INVX1_147 ( .A(_9__2_), .Y(_89_) );
NAND2X1 NAND2X1_246 ( .A(w_cout_1_), .B(_10__2_), .Y(_90_) );
OAI21X1 OAI21X1_246 ( .A(w_cout_1_), .B(_89_), .C(_90_), .Y(_0__9_) );
INVX1 INVX1_148 ( .A(_9__3_), .Y(_91_) );
NAND2X1 NAND2X1_247 ( .A(w_cout_1_), .B(_10__3_), .Y(_92_) );
OAI21X1 OAI21X1_247 ( .A(w_cout_1_), .B(_91_), .C(_92_), .Y(_0__10_) );
INVX1 INVX1_149 ( .A(_13_), .Y(_93_) );
NAND2X1 NAND2X1_248 ( .A(_14_), .B(w_cout_2_), .Y(_94_) );
OAI21X1 OAI21X1_248 ( .A(w_cout_2_), .B(_93_), .C(_94_), .Y(w_cout_3_) );
INVX1 INVX1_150 ( .A(_15__0_), .Y(_95_) );
NAND2X1 NAND2X1_249 ( .A(_16__0_), .B(w_cout_2_), .Y(_96_) );
OAI21X1 OAI21X1_249 ( .A(w_cout_2_), .B(_95_), .C(_96_), .Y(_0__11_) );
INVX1 INVX1_151 ( .A(_15__1_), .Y(_97_) );
NAND2X1 NAND2X1_250 ( .A(w_cout_2_), .B(_16__1_), .Y(_98_) );
OAI21X1 OAI21X1_250 ( .A(w_cout_2_), .B(_97_), .C(_98_), .Y(_0__12_) );
INVX1 INVX1_152 ( .A(_15__2_), .Y(_99_) );
NAND2X1 NAND2X1_251 ( .A(w_cout_2_), .B(_16__2_), .Y(_100_) );
OAI21X1 OAI21X1_251 ( .A(w_cout_2_), .B(_99_), .C(_100_), .Y(_0__13_) );
INVX1 INVX1_153 ( .A(_15__3_), .Y(_101_) );
NAND2X1 NAND2X1_252 ( .A(w_cout_2_), .B(_16__3_), .Y(_102_) );
OAI21X1 OAI21X1_252 ( .A(w_cout_2_), .B(_101_), .C(_102_), .Y(_0__14_) );
INVX1 INVX1_154 ( .A(_19_), .Y(_103_) );
NAND2X1 NAND2X1_253 ( .A(_20_), .B(w_cout_3_), .Y(_104_) );
OAI21X1 OAI21X1_253 ( .A(w_cout_3_), .B(_103_), .C(_104_), .Y(w_cout_4_) );
INVX1 INVX1_155 ( .A(_21__0_), .Y(_105_) );
NAND2X1 NAND2X1_254 ( .A(_22__0_), .B(w_cout_3_), .Y(_106_) );
OAI21X1 OAI21X1_254 ( .A(w_cout_3_), .B(_105_), .C(_106_), .Y(_0__15_) );
INVX1 INVX1_156 ( .A(_21__1_), .Y(_107_) );
NAND2X1 NAND2X1_255 ( .A(w_cout_3_), .B(_22__1_), .Y(_108_) );
OAI21X1 OAI21X1_255 ( .A(w_cout_3_), .B(_107_), .C(_108_), .Y(_0__16_) );
INVX1 INVX1_157 ( .A(_21__2_), .Y(_109_) );
NAND2X1 NAND2X1_256 ( .A(w_cout_3_), .B(_22__2_), .Y(_110_) );
OAI21X1 OAI21X1_256 ( .A(w_cout_3_), .B(_109_), .C(_110_), .Y(_0__17_) );
INVX1 INVX1_158 ( .A(_21__3_), .Y(_111_) );
NAND2X1 NAND2X1_257 ( .A(w_cout_3_), .B(_22__3_), .Y(_112_) );
OAI21X1 OAI21X1_257 ( .A(w_cout_3_), .B(_111_), .C(_112_), .Y(_0__18_) );
INVX1 INVX1_159 ( .A(_25_), .Y(_113_) );
NAND2X1 NAND2X1_258 ( .A(_26_), .B(w_cout_4_), .Y(_114_) );
BUFX2 BUFX2_53 ( .A(1'b0), .Y(_5__0_) );
BUFX2 BUFX2_54 ( .A(_1_), .Y(_5__4_) );
BUFX2 BUFX2_55 ( .A(1'b1), .Y(_6__0_) );
BUFX2 BUFX2_56 ( .A(_2_), .Y(_6__4_) );
BUFX2 BUFX2_57 ( .A(1'b0), .Y(_11__0_) );
BUFX2 BUFX2_58 ( .A(_7_), .Y(_11__4_) );
BUFX2 BUFX2_59 ( .A(1'b1), .Y(_12__0_) );
BUFX2 BUFX2_60 ( .A(_8_), .Y(_12__4_) );
BUFX2 BUFX2_61 ( .A(1'b0), .Y(_17__0_) );
BUFX2 BUFX2_62 ( .A(_13_), .Y(_17__4_) );
BUFX2 BUFX2_63 ( .A(1'b1), .Y(_18__0_) );
BUFX2 BUFX2_64 ( .A(_14_), .Y(_18__4_) );
BUFX2 BUFX2_65 ( .A(1'b0), .Y(_23__0_) );
BUFX2 BUFX2_66 ( .A(_19_), .Y(_23__4_) );
BUFX2 BUFX2_67 ( .A(1'b1), .Y(_24__0_) );
BUFX2 BUFX2_68 ( .A(_20_), .Y(_24__4_) );
BUFX2 BUFX2_69 ( .A(1'b0), .Y(_29__0_) );
BUFX2 BUFX2_70 ( .A(_25_), .Y(_29__4_) );
BUFX2 BUFX2_71 ( .A(1'b1), .Y(_30__0_) );
BUFX2 BUFX2_72 ( .A(_26_), .Y(_30__4_) );
BUFX2 BUFX2_73 ( .A(1'b0), .Y(_35__0_) );
BUFX2 BUFX2_74 ( .A(_31_), .Y(_35__4_) );
BUFX2 BUFX2_75 ( .A(1'b1), .Y(_36__0_) );
BUFX2 BUFX2_76 ( .A(_32_), .Y(_36__4_) );
BUFX2 BUFX2_77 ( .A(1'b0), .Y(_41__0_) );
BUFX2 BUFX2_78 ( .A(_37_), .Y(_41__4_) );
BUFX2 BUFX2_79 ( .A(1'b1), .Y(_42__0_) );
BUFX2 BUFX2_80 ( .A(_38_), .Y(_42__4_) );
BUFX2 BUFX2_81 ( .A(1'b0), .Y(_47__0_) );
BUFX2 BUFX2_82 ( .A(_43_), .Y(_47__4_) );
BUFX2 BUFX2_83 ( .A(1'b1), .Y(_48__0_) );
BUFX2 BUFX2_84 ( .A(_44_), .Y(_48__4_) );
BUFX2 BUFX2_85 ( .A(1'b0), .Y(_53__0_) );
BUFX2 BUFX2_86 ( .A(_49_), .Y(_53__4_) );
BUFX2 BUFX2_87 ( .A(1'b1), .Y(_54__0_) );
BUFX2 BUFX2_88 ( .A(_50_), .Y(_54__4_) );
BUFX2 BUFX2_89 ( .A(1'b0), .Y(_59__0_) );
BUFX2 BUFX2_90 ( .A(_55_), .Y(_59__4_) );
BUFX2 BUFX2_91 ( .A(1'b1), .Y(_60__0_) );
BUFX2 BUFX2_92 ( .A(_56_), .Y(_60__4_) );
BUFX2 BUFX2_93 ( .A(1'b0), .Y(_65__0_) );
BUFX2 BUFX2_94 ( .A(_61_), .Y(_65__4_) );
BUFX2 BUFX2_95 ( .A(1'b1), .Y(_66__0_) );
BUFX2 BUFX2_96 ( .A(_62_), .Y(_66__4_) );
BUFX2 BUFX2_97 ( .A(1'b0), .Y(_71__0_) );
BUFX2 BUFX2_98 ( .A(_67_), .Y(_71__4_) );
BUFX2 BUFX2_99 ( .A(1'b1), .Y(_72__0_) );
BUFX2 BUFX2_100 ( .A(_68_), .Y(_72__4_) );
BUFX2 BUFX2_101 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_102 ( .A(1'b0), .Y(w_cout_0_) );
endmodule
