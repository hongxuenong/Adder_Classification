module cla_26bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add1[19], i_add1[20], i_add1[21], i_add1[22], i_add1[23], i_add1[24], i_add1[25], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], i_add2[19], i_add2[20], i_add2[21], i_add2[22], i_add2[23], i_add2[24], i_add2[25], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19], o_result[20], o_result[21], o_result[22], o_result[23], o_result[24], o_result[25], o_result[26]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add1[19];
input i_add1[20];
input i_add1[21];
input i_add1[22];
input i_add1[23];
input i_add1[24];
input i_add1[25];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
input i_add2[19];
input i_add2[20];
input i_add2[21];
input i_add2[22];
input i_add2[23];
input i_add2[24];
input i_add2[25];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];
output o_result[20];
output o_result[21];
output o_result[22];
output o_result[23];
output o_result[24];
output o_result[25];
output o_result[26];

NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_117_) );
INVX1 INVX1_1 ( .A(_117_), .Y(w_C_1_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_118_) );
AOI22X1 AOI22X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_119_) );
NOR2X1 NOR2X1_2 ( .A(_118_), .B(_119_), .Y(w_C_2_) );
INVX1 INVX1_2 ( .A(i_add2[2]), .Y(_120_) );
INVX1 INVX1_3 ( .A(i_add1[2]), .Y(_121_) );
NAND2X1 NAND2X1_2 ( .A(_120_), .B(_121_), .Y(_122_) );
NAND2X1 NAND2X1_3 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_123_) );
OAI21X1 OAI21X1_1 ( .A(_118_), .B(_119_), .C(_123_), .Y(_124_) );
AND2X2 AND2X2_1 ( .A(_124_), .B(_122_), .Y(w_C_3_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_125_) );
OR2X2 OR2X2_1 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_126_) );
NAND3X1 NAND3X1_1 ( .A(_122_), .B(_126_), .C(_124_), .Y(_127_) );
NAND2X1 NAND2X1_5 ( .A(_125_), .B(_127_), .Y(w_C_4_) );
NOR2X1 NOR2X1_3 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_128_) );
INVX1 INVX1_4 ( .A(_128_), .Y(_129_) );
NAND2X1 NAND2X1_6 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_130_) );
NAND3X1 NAND3X1_2 ( .A(_125_), .B(_130_), .C(_127_), .Y(_131_) );
AND2X2 AND2X2_2 ( .A(_131_), .B(_129_), .Y(w_C_5_) );
INVX1 INVX1_5 ( .A(i_add2[5]), .Y(_132_) );
INVX1 INVX1_6 ( .A(i_add1[5]), .Y(_0_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_1_) );
INVX1 INVX1_7 ( .A(_1_), .Y(_2_) );
NAND3X1 NAND3X1_3 ( .A(_129_), .B(_2_), .C(_131_), .Y(_3_) );
OAI21X1 OAI21X1_2 ( .A(_132_), .B(_0_), .C(_3_), .Y(w_C_6_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_4_) );
INVX1 INVX1_8 ( .A(_4_), .Y(_5_) );
NOR2X1 NOR2X1_6 ( .A(_132_), .B(_0_), .Y(_6_) );
INVX1 INVX1_9 ( .A(_6_), .Y(_7_) );
AND2X2 AND2X2_3 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_8_) );
INVX1 INVX1_10 ( .A(_8_), .Y(_9_) );
NAND3X1 NAND3X1_4 ( .A(_7_), .B(_9_), .C(_3_), .Y(_10_) );
AND2X2 AND2X2_4 ( .A(_10_), .B(_5_), .Y(w_C_7_) );
AND2X2 AND2X2_5 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_11_) );
INVX1 INVX1_11 ( .A(_11_), .Y(_12_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_13_) );
INVX1 INVX1_12 ( .A(_13_), .Y(_14_) );
NAND3X1 NAND3X1_5 ( .A(_5_), .B(_14_), .C(_10_), .Y(_15_) );
AND2X2 AND2X2_6 ( .A(_15_), .B(_12_), .Y(_16_) );
INVX1 INVX1_13 ( .A(_16_), .Y(w_C_8_) );
AND2X2 AND2X2_7 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_17_) );
INVX1 INVX1_14 ( .A(_17_), .Y(_18_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_19_) );
OAI21X1 OAI21X1_3 ( .A(_19_), .B(_16_), .C(_18_), .Y(w_C_9_) );
AND2X2 AND2X2_8 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_20_) );
INVX1 INVX1_15 ( .A(_20_), .Y(_21_) );
INVX1 INVX1_16 ( .A(_19_), .Y(_22_) );
NAND3X1 NAND3X1_6 ( .A(_12_), .B(_18_), .C(_15_), .Y(_23_) );
NOR2X1 NOR2X1_9 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_24_) );
INVX1 INVX1_17 ( .A(_24_), .Y(_25_) );
NAND3X1 NAND3X1_7 ( .A(_22_), .B(_25_), .C(_23_), .Y(_26_) );
AND2X2 AND2X2_9 ( .A(_26_), .B(_21_), .Y(_27_) );
INVX1 INVX1_18 ( .A(_27_), .Y(w_C_10_) );
AND2X2 AND2X2_10 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_28_) );
INVX1 INVX1_19 ( .A(_28_), .Y(_29_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_30_) );
OAI21X1 OAI21X1_4 ( .A(_30_), .B(_27_), .C(_29_), .Y(w_C_11_) );
INVX1 INVX1_20 ( .A(i_add2[11]), .Y(_31_) );
INVX1 INVX1_21 ( .A(i_add1[11]), .Y(_32_) );
INVX1 INVX1_22 ( .A(_30_), .Y(_33_) );
NAND3X1 NAND3X1_8 ( .A(_21_), .B(_29_), .C(_26_), .Y(_34_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_35_) );
INVX1 INVX1_23 ( .A(_35_), .Y(_36_) );
NAND3X1 NAND3X1_9 ( .A(_33_), .B(_36_), .C(_34_), .Y(_37_) );
OAI21X1 OAI21X1_5 ( .A(_31_), .B(_32_), .C(_37_), .Y(w_C_12_) );
NOR2X1 NOR2X1_12 ( .A(_31_), .B(_32_), .Y(_38_) );
INVX1 INVX1_24 ( .A(_38_), .Y(_39_) );
AND2X2 AND2X2_11 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_40_) );
INVX1 INVX1_25 ( .A(_40_), .Y(_41_) );
NAND3X1 NAND3X1_10 ( .A(_39_), .B(_41_), .C(_37_), .Y(_42_) );
OAI21X1 OAI21X1_6 ( .A(i_add2[12]), .B(i_add1[12]), .C(_42_), .Y(_43_) );
INVX1 INVX1_26 ( .A(_43_), .Y(w_C_13_) );
INVX1 INVX1_27 ( .A(i_add2[13]), .Y(_44_) );
INVX1 INVX1_28 ( .A(i_add1[13]), .Y(_45_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_46_) );
INVX1 INVX1_29 ( .A(_46_), .Y(_47_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_48_) );
INVX1 INVX1_30 ( .A(_48_), .Y(_49_) );
NAND3X1 NAND3X1_11 ( .A(_47_), .B(_49_), .C(_42_), .Y(_50_) );
OAI21X1 OAI21X1_7 ( .A(_44_), .B(_45_), .C(_50_), .Y(w_C_14_) );
NOR2X1 NOR2X1_15 ( .A(_44_), .B(_45_), .Y(_51_) );
INVX1 INVX1_31 ( .A(_51_), .Y(_52_) );
AND2X2 AND2X2_12 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_53_) );
INVX1 INVX1_32 ( .A(_53_), .Y(_54_) );
NAND3X1 NAND3X1_12 ( .A(_52_), .B(_54_), .C(_50_), .Y(_55_) );
OAI21X1 OAI21X1_8 ( .A(i_add2[14]), .B(i_add1[14]), .C(_55_), .Y(_56_) );
INVX1 INVX1_33 ( .A(_56_), .Y(w_C_15_) );
INVX1 INVX1_34 ( .A(i_add2[15]), .Y(_57_) );
INVX1 INVX1_35 ( .A(i_add1[15]), .Y(_58_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_59_) );
INVX1 INVX1_36 ( .A(_59_), .Y(_60_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_61_) );
INVX1 INVX1_37 ( .A(_61_), .Y(_62_) );
NAND3X1 NAND3X1_13 ( .A(_60_), .B(_62_), .C(_55_), .Y(_63_) );
OAI21X1 OAI21X1_9 ( .A(_57_), .B(_58_), .C(_63_), .Y(w_C_16_) );
NOR2X1 NOR2X1_18 ( .A(_57_), .B(_58_), .Y(_64_) );
INVX1 INVX1_38 ( .A(_64_), .Y(_65_) );
AND2X2 AND2X2_13 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_66_) );
INVX1 INVX1_39 ( .A(_66_), .Y(_67_) );
NAND3X1 NAND3X1_14 ( .A(_65_), .B(_67_), .C(_63_), .Y(_68_) );
OAI21X1 OAI21X1_10 ( .A(i_add2[16]), .B(i_add1[16]), .C(_68_), .Y(_69_) );
INVX1 INVX1_40 ( .A(_69_), .Y(w_C_17_) );
INVX1 INVX1_41 ( .A(i_add2[17]), .Y(_70_) );
INVX1 INVX1_42 ( .A(i_add1[17]), .Y(_71_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_72_) );
INVX1 INVX1_43 ( .A(_72_), .Y(_73_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_74_) );
INVX1 INVX1_44 ( .A(_74_), .Y(_75_) );
NAND3X1 NAND3X1_15 ( .A(_73_), .B(_75_), .C(_68_), .Y(_76_) );
OAI21X1 OAI21X1_11 ( .A(_70_), .B(_71_), .C(_76_), .Y(w_C_18_) );
NOR2X1 NOR2X1_21 ( .A(_70_), .B(_71_), .Y(_77_) );
INVX1 INVX1_45 ( .A(_77_), .Y(_78_) );
AND2X2 AND2X2_14 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_79_) );
INVX1 INVX1_46 ( .A(_79_), .Y(_80_) );
NAND3X1 NAND3X1_16 ( .A(_78_), .B(_80_), .C(_76_), .Y(_81_) );
OAI21X1 OAI21X1_12 ( .A(i_add2[18]), .B(i_add1[18]), .C(_81_), .Y(_82_) );
INVX1 INVX1_47 ( .A(_82_), .Y(w_C_19_) );
INVX1 INVX1_48 ( .A(i_add2[19]), .Y(_83_) );
INVX1 INVX1_49 ( .A(i_add1[19]), .Y(_84_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_85_) );
INVX1 INVX1_50 ( .A(_85_), .Y(_86_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_87_) );
INVX1 INVX1_51 ( .A(_87_), .Y(_88_) );
NAND3X1 NAND3X1_17 ( .A(_86_), .B(_88_), .C(_81_), .Y(_89_) );
OAI21X1 OAI21X1_13 ( .A(_83_), .B(_84_), .C(_89_), .Y(w_C_20_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_90_) );
INVX1 INVX1_52 ( .A(_90_), .Y(_91_) );
NOR2X1 NOR2X1_25 ( .A(_83_), .B(_84_), .Y(_92_) );
INVX1 INVX1_53 ( .A(_92_), .Y(_93_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_94_) );
NAND3X1 NAND3X1_18 ( .A(_93_), .B(_94_), .C(_89_), .Y(_95_) );
AND2X2 AND2X2_15 ( .A(_95_), .B(_91_), .Y(w_C_21_) );
INVX1 INVX1_54 ( .A(i_add2[21]), .Y(_96_) );
INVX1 INVX1_55 ( .A(i_add1[21]), .Y(_97_) );
NAND2X1 NAND2X1_8 ( .A(_96_), .B(_97_), .Y(_98_) );
NAND3X1 NAND3X1_19 ( .A(_91_), .B(_98_), .C(_95_), .Y(_99_) );
OAI21X1 OAI21X1_14 ( .A(_96_), .B(_97_), .C(_99_), .Y(w_C_22_) );
INVX1 INVX1_56 ( .A(i_add2[22]), .Y(_100_) );
INVX1 INVX1_57 ( .A(i_add1[22]), .Y(_101_) );
NAND2X1 NAND2X1_9 ( .A(_100_), .B(_101_), .Y(_102_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_103_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_104_) );
NAND3X1 NAND3X1_20 ( .A(_103_), .B(_104_), .C(_99_), .Y(_105_) );
AND2X2 AND2X2_16 ( .A(_105_), .B(_102_), .Y(w_C_23_) );
INVX1 INVX1_58 ( .A(i_add2[23]), .Y(_106_) );
INVX1 INVX1_59 ( .A(i_add1[23]), .Y(_107_) );
NAND2X1 NAND2X1_12 ( .A(_106_), .B(_107_), .Y(_108_) );
NAND3X1 NAND3X1_21 ( .A(_102_), .B(_108_), .C(_105_), .Y(_109_) );
OAI21X1 OAI21X1_15 ( .A(_106_), .B(_107_), .C(_109_), .Y(w_C_24_) );
OR2X2 OR2X2_2 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_110_) );
NAND2X1 NAND2X1_13 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_111_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_112_) );
NAND3X1 NAND3X1_22 ( .A(_111_), .B(_112_), .C(_109_), .Y(_113_) );
AND2X2 AND2X2_17 ( .A(_113_), .B(_110_), .Y(w_C_25_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_114_) );
OR2X2 OR2X2_3 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_115_) );
NAND3X1 NAND3X1_23 ( .A(_110_), .B(_115_), .C(_113_), .Y(_116_) );
NAND2X1 NAND2X1_16 ( .A(_114_), .B(_116_), .Y(w_C_26_) );
BUFX2 BUFX2_1 ( .A(_133__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_133__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_133__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_133__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_133__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_133__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_133__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_133__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_133__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_133__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_133__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_133__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_133__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_133__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_133__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_133__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_133__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_133__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_133__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(_133__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .A(_133__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .A(_133__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .A(_133__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .A(_133__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .A(_133__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .A(_133__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .A(w_C_26_), .Y(o_result[26]) );
INVX1 INVX1_60 ( .A(w_C_4_), .Y(_137_) );
OR2X2 OR2X2_4 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_138_) );
NAND2X1 NAND2X1_17 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_139_) );
NAND3X1 NAND3X1_24 ( .A(_137_), .B(_139_), .C(_138_), .Y(_140_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_134_) );
AND2X2 AND2X2_18 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_135_) );
OAI21X1 OAI21X1_16 ( .A(_134_), .B(_135_), .C(w_C_4_), .Y(_136_) );
NAND2X1 NAND2X1_18 ( .A(_136_), .B(_140_), .Y(_133__4_) );
INVX1 INVX1_61 ( .A(w_C_5_), .Y(_144_) );
OR2X2 OR2X2_5 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_145_) );
NAND2X1 NAND2X1_19 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_146_) );
NAND3X1 NAND3X1_25 ( .A(_144_), .B(_146_), .C(_145_), .Y(_147_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_141_) );
AND2X2 AND2X2_19 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_142_) );
OAI21X1 OAI21X1_17 ( .A(_141_), .B(_142_), .C(w_C_5_), .Y(_143_) );
NAND2X1 NAND2X1_20 ( .A(_143_), .B(_147_), .Y(_133__5_) );
INVX1 INVX1_62 ( .A(w_C_6_), .Y(_151_) );
OR2X2 OR2X2_6 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_152_) );
NAND2X1 NAND2X1_21 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_153_) );
NAND3X1 NAND3X1_26 ( .A(_151_), .B(_153_), .C(_152_), .Y(_154_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_148_) );
AND2X2 AND2X2_20 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_149_) );
OAI21X1 OAI21X1_18 ( .A(_148_), .B(_149_), .C(w_C_6_), .Y(_150_) );
NAND2X1 NAND2X1_22 ( .A(_150_), .B(_154_), .Y(_133__6_) );
INVX1 INVX1_63 ( .A(w_C_7_), .Y(_158_) );
OR2X2 OR2X2_7 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_159_) );
NAND2X1 NAND2X1_23 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_160_) );
NAND3X1 NAND3X1_27 ( .A(_158_), .B(_160_), .C(_159_), .Y(_161_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_155_) );
AND2X2 AND2X2_21 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_156_) );
OAI21X1 OAI21X1_19 ( .A(_155_), .B(_156_), .C(w_C_7_), .Y(_157_) );
NAND2X1 NAND2X1_24 ( .A(_157_), .B(_161_), .Y(_133__7_) );
INVX1 INVX1_64 ( .A(w_C_8_), .Y(_165_) );
OR2X2 OR2X2_8 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_166_) );
NAND2X1 NAND2X1_25 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_167_) );
NAND3X1 NAND3X1_28 ( .A(_165_), .B(_167_), .C(_166_), .Y(_168_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_162_) );
AND2X2 AND2X2_22 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_163_) );
OAI21X1 OAI21X1_20 ( .A(_162_), .B(_163_), .C(w_C_8_), .Y(_164_) );
NAND2X1 NAND2X1_26 ( .A(_164_), .B(_168_), .Y(_133__8_) );
INVX1 INVX1_65 ( .A(w_C_9_), .Y(_172_) );
OR2X2 OR2X2_9 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_173_) );
NAND2X1 NAND2X1_27 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_174_) );
NAND3X1 NAND3X1_29 ( .A(_172_), .B(_174_), .C(_173_), .Y(_175_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_169_) );
AND2X2 AND2X2_23 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_170_) );
OAI21X1 OAI21X1_21 ( .A(_169_), .B(_170_), .C(w_C_9_), .Y(_171_) );
NAND2X1 NAND2X1_28 ( .A(_171_), .B(_175_), .Y(_133__9_) );
INVX1 INVX1_66 ( .A(w_C_10_), .Y(_179_) );
OR2X2 OR2X2_10 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_180_) );
NAND2X1 NAND2X1_29 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_181_) );
NAND3X1 NAND3X1_30 ( .A(_179_), .B(_181_), .C(_180_), .Y(_182_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_176_) );
AND2X2 AND2X2_24 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_177_) );
OAI21X1 OAI21X1_22 ( .A(_176_), .B(_177_), .C(w_C_10_), .Y(_178_) );
NAND2X1 NAND2X1_30 ( .A(_178_), .B(_182_), .Y(_133__10_) );
INVX1 INVX1_67 ( .A(w_C_11_), .Y(_186_) );
OR2X2 OR2X2_11 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_187_) );
NAND2X1 NAND2X1_31 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_188_) );
NAND3X1 NAND3X1_31 ( .A(_186_), .B(_188_), .C(_187_), .Y(_189_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_183_) );
AND2X2 AND2X2_25 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_184_) );
OAI21X1 OAI21X1_23 ( .A(_183_), .B(_184_), .C(w_C_11_), .Y(_185_) );
NAND2X1 NAND2X1_32 ( .A(_185_), .B(_189_), .Y(_133__11_) );
INVX1 INVX1_68 ( .A(w_C_12_), .Y(_193_) );
OR2X2 OR2X2_12 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_194_) );
NAND2X1 NAND2X1_33 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_195_) );
NAND3X1 NAND3X1_32 ( .A(_193_), .B(_195_), .C(_194_), .Y(_196_) );
NOR2X1 NOR2X1_34 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_190_) );
AND2X2 AND2X2_26 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_191_) );
OAI21X1 OAI21X1_24 ( .A(_190_), .B(_191_), .C(w_C_12_), .Y(_192_) );
NAND2X1 NAND2X1_34 ( .A(_192_), .B(_196_), .Y(_133__12_) );
INVX1 INVX1_69 ( .A(w_C_13_), .Y(_200_) );
OR2X2 OR2X2_13 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_201_) );
NAND2X1 NAND2X1_35 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_202_) );
NAND3X1 NAND3X1_33 ( .A(_200_), .B(_202_), .C(_201_), .Y(_203_) );
NOR2X1 NOR2X1_35 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_197_) );
AND2X2 AND2X2_27 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_198_) );
OAI21X1 OAI21X1_25 ( .A(_197_), .B(_198_), .C(w_C_13_), .Y(_199_) );
NAND2X1 NAND2X1_36 ( .A(_199_), .B(_203_), .Y(_133__13_) );
INVX1 INVX1_70 ( .A(w_C_14_), .Y(_207_) );
OR2X2 OR2X2_14 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_208_) );
NAND2X1 NAND2X1_37 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_209_) );
NAND3X1 NAND3X1_34 ( .A(_207_), .B(_209_), .C(_208_), .Y(_210_) );
NOR2X1 NOR2X1_36 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_204_) );
AND2X2 AND2X2_28 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_205_) );
OAI21X1 OAI21X1_26 ( .A(_204_), .B(_205_), .C(w_C_14_), .Y(_206_) );
NAND2X1 NAND2X1_38 ( .A(_206_), .B(_210_), .Y(_133__14_) );
INVX1 INVX1_71 ( .A(w_C_15_), .Y(_214_) );
OR2X2 OR2X2_15 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_215_) );
NAND2X1 NAND2X1_39 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_216_) );
NAND3X1 NAND3X1_35 ( .A(_214_), .B(_216_), .C(_215_), .Y(_217_) );
NOR2X1 NOR2X1_37 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_211_) );
AND2X2 AND2X2_29 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_212_) );
OAI21X1 OAI21X1_27 ( .A(_211_), .B(_212_), .C(w_C_15_), .Y(_213_) );
NAND2X1 NAND2X1_40 ( .A(_213_), .B(_217_), .Y(_133__15_) );
INVX1 INVX1_72 ( .A(w_C_16_), .Y(_221_) );
OR2X2 OR2X2_16 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_222_) );
NAND2X1 NAND2X1_41 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_223_) );
NAND3X1 NAND3X1_36 ( .A(_221_), .B(_223_), .C(_222_), .Y(_224_) );
NOR2X1 NOR2X1_38 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_218_) );
AND2X2 AND2X2_30 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_219_) );
OAI21X1 OAI21X1_28 ( .A(_218_), .B(_219_), .C(w_C_16_), .Y(_220_) );
NAND2X1 NAND2X1_42 ( .A(_220_), .B(_224_), .Y(_133__16_) );
INVX1 INVX1_73 ( .A(w_C_17_), .Y(_228_) );
OR2X2 OR2X2_17 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_229_) );
NAND2X1 NAND2X1_43 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_230_) );
NAND3X1 NAND3X1_37 ( .A(_228_), .B(_230_), .C(_229_), .Y(_231_) );
NOR2X1 NOR2X1_39 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_225_) );
AND2X2 AND2X2_31 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_226_) );
OAI21X1 OAI21X1_29 ( .A(_225_), .B(_226_), .C(w_C_17_), .Y(_227_) );
NAND2X1 NAND2X1_44 ( .A(_227_), .B(_231_), .Y(_133__17_) );
INVX1 INVX1_74 ( .A(w_C_18_), .Y(_235_) );
OR2X2 OR2X2_18 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_236_) );
NAND2X1 NAND2X1_45 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_237_) );
NAND3X1 NAND3X1_38 ( .A(_235_), .B(_237_), .C(_236_), .Y(_238_) );
NOR2X1 NOR2X1_40 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_232_) );
AND2X2 AND2X2_32 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_233_) );
OAI21X1 OAI21X1_30 ( .A(_232_), .B(_233_), .C(w_C_18_), .Y(_234_) );
NAND2X1 NAND2X1_46 ( .A(_234_), .B(_238_), .Y(_133__18_) );
INVX1 INVX1_75 ( .A(w_C_19_), .Y(_242_) );
OR2X2 OR2X2_19 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_243_) );
NAND2X1 NAND2X1_47 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_244_) );
NAND3X1 NAND3X1_39 ( .A(_242_), .B(_244_), .C(_243_), .Y(_245_) );
NOR2X1 NOR2X1_41 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_239_) );
AND2X2 AND2X2_33 ( .A(i_add2[19]), .B(i_add1[19]), .Y(_240_) );
OAI21X1 OAI21X1_31 ( .A(_239_), .B(_240_), .C(w_C_19_), .Y(_241_) );
NAND2X1 NAND2X1_48 ( .A(_241_), .B(_245_), .Y(_133__19_) );
INVX1 INVX1_76 ( .A(w_C_20_), .Y(_249_) );
OR2X2 OR2X2_20 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_250_) );
NAND2X1 NAND2X1_49 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_251_) );
NAND3X1 NAND3X1_40 ( .A(_249_), .B(_251_), .C(_250_), .Y(_252_) );
NOR2X1 NOR2X1_42 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_246_) );
AND2X2 AND2X2_34 ( .A(i_add2[20]), .B(i_add1[20]), .Y(_247_) );
OAI21X1 OAI21X1_32 ( .A(_246_), .B(_247_), .C(w_C_20_), .Y(_248_) );
NAND2X1 NAND2X1_50 ( .A(_248_), .B(_252_), .Y(_133__20_) );
INVX1 INVX1_77 ( .A(w_C_21_), .Y(_256_) );
OR2X2 OR2X2_21 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_257_) );
NAND2X1 NAND2X1_51 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_258_) );
NAND3X1 NAND3X1_41 ( .A(_256_), .B(_258_), .C(_257_), .Y(_259_) );
NOR2X1 NOR2X1_43 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_253_) );
AND2X2 AND2X2_35 ( .A(i_add2[21]), .B(i_add1[21]), .Y(_254_) );
OAI21X1 OAI21X1_33 ( .A(_253_), .B(_254_), .C(w_C_21_), .Y(_255_) );
NAND2X1 NAND2X1_52 ( .A(_255_), .B(_259_), .Y(_133__21_) );
INVX1 INVX1_78 ( .A(w_C_22_), .Y(_263_) );
OR2X2 OR2X2_22 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_264_) );
NAND2X1 NAND2X1_53 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_265_) );
NAND3X1 NAND3X1_42 ( .A(_263_), .B(_265_), .C(_264_), .Y(_266_) );
NOR2X1 NOR2X1_44 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_260_) );
AND2X2 AND2X2_36 ( .A(i_add2[22]), .B(i_add1[22]), .Y(_261_) );
OAI21X1 OAI21X1_34 ( .A(_260_), .B(_261_), .C(w_C_22_), .Y(_262_) );
NAND2X1 NAND2X1_54 ( .A(_262_), .B(_266_), .Y(_133__22_) );
INVX1 INVX1_79 ( .A(w_C_23_), .Y(_270_) );
OR2X2 OR2X2_23 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_271_) );
NAND2X1 NAND2X1_55 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_272_) );
NAND3X1 NAND3X1_43 ( .A(_270_), .B(_272_), .C(_271_), .Y(_273_) );
NOR2X1 NOR2X1_45 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_267_) );
AND2X2 AND2X2_37 ( .A(i_add2[23]), .B(i_add1[23]), .Y(_268_) );
OAI21X1 OAI21X1_35 ( .A(_267_), .B(_268_), .C(w_C_23_), .Y(_269_) );
NAND2X1 NAND2X1_56 ( .A(_269_), .B(_273_), .Y(_133__23_) );
INVX1 INVX1_80 ( .A(w_C_24_), .Y(_277_) );
OR2X2 OR2X2_24 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_278_) );
NAND2X1 NAND2X1_57 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_279_) );
NAND3X1 NAND3X1_44 ( .A(_277_), .B(_279_), .C(_278_), .Y(_280_) );
NOR2X1 NOR2X1_46 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_274_) );
AND2X2 AND2X2_38 ( .A(i_add2[24]), .B(i_add1[24]), .Y(_275_) );
OAI21X1 OAI21X1_36 ( .A(_274_), .B(_275_), .C(w_C_24_), .Y(_276_) );
NAND2X1 NAND2X1_58 ( .A(_276_), .B(_280_), .Y(_133__24_) );
INVX1 INVX1_81 ( .A(w_C_25_), .Y(_284_) );
OR2X2 OR2X2_25 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_285_) );
NAND2X1 NAND2X1_59 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_286_) );
NAND3X1 NAND3X1_45 ( .A(_284_), .B(_286_), .C(_285_), .Y(_287_) );
NOR2X1 NOR2X1_47 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_281_) );
AND2X2 AND2X2_39 ( .A(i_add2[25]), .B(i_add1[25]), .Y(_282_) );
OAI21X1 OAI21X1_37 ( .A(_281_), .B(_282_), .C(w_C_25_), .Y(_283_) );
NAND2X1 NAND2X1_60 ( .A(_283_), .B(_287_), .Y(_133__25_) );
INVX1 INVX1_82 ( .A(1'b0), .Y(_291_) );
OR2X2 OR2X2_26 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_292_) );
NAND2X1 NAND2X1_61 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_293_) );
NAND3X1 NAND3X1_46 ( .A(_291_), .B(_293_), .C(_292_), .Y(_294_) );
NOR2X1 NOR2X1_48 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_288_) );
AND2X2 AND2X2_40 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_289_) );
OAI21X1 OAI21X1_38 ( .A(_288_), .B(_289_), .C(1'b0), .Y(_290_) );
NAND2X1 NAND2X1_62 ( .A(_290_), .B(_294_), .Y(_133__0_) );
INVX1 INVX1_83 ( .A(w_C_1_), .Y(_298_) );
OR2X2 OR2X2_27 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_299_) );
NAND2X1 NAND2X1_63 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_300_) );
NAND3X1 NAND3X1_47 ( .A(_298_), .B(_300_), .C(_299_), .Y(_301_) );
NOR2X1 NOR2X1_49 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_295_) );
AND2X2 AND2X2_41 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_296_) );
OAI21X1 OAI21X1_39 ( .A(_295_), .B(_296_), .C(w_C_1_), .Y(_297_) );
NAND2X1 NAND2X1_64 ( .A(_297_), .B(_301_), .Y(_133__1_) );
INVX1 INVX1_84 ( .A(w_C_2_), .Y(_305_) );
OR2X2 OR2X2_28 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_306_) );
NAND2X1 NAND2X1_65 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_307_) );
NAND3X1 NAND3X1_48 ( .A(_305_), .B(_307_), .C(_306_), .Y(_308_) );
NOR2X1 NOR2X1_50 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_302_) );
AND2X2 AND2X2_42 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_303_) );
OAI21X1 OAI21X1_40 ( .A(_302_), .B(_303_), .C(w_C_2_), .Y(_304_) );
NAND2X1 NAND2X1_66 ( .A(_304_), .B(_308_), .Y(_133__2_) );
INVX1 INVX1_85 ( .A(w_C_3_), .Y(_312_) );
OR2X2 OR2X2_29 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_313_) );
NAND2X1 NAND2X1_67 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_314_) );
NAND3X1 NAND3X1_49 ( .A(_312_), .B(_314_), .C(_313_), .Y(_315_) );
NOR2X1 NOR2X1_51 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_309_) );
AND2X2 AND2X2_43 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_310_) );
OAI21X1 OAI21X1_41 ( .A(_309_), .B(_310_), .C(w_C_3_), .Y(_311_) );
NAND2X1 NAND2X1_68 ( .A(_311_), .B(_315_), .Y(_133__3_) );
BUFX2 BUFX2_28 ( .A(w_C_26_), .Y(_133__26_) );
BUFX2 BUFX2_29 ( .A(1'b0), .Y(w_C_0_) );
endmodule
