module CSkipA_18bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [17:0] i_add_term1;
input [17:0] i_add_term2;
output [17:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX2 BUFX2_1 ( .A(w_cout_5_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
INVX1 INVX1_1 ( .A(i_add_term1[0]), .Y(_13_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[0]), .B(_13_), .Y(_14_) );
INVX1 INVX1_2 ( .A(i_add_term2[0]), .Y(_15_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term1[0]), .B(_15_), .Y(_16_) );
INVX1 INVX1_3 ( .A(i_add_term1[1]), .Y(_17_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[1]), .B(_17_), .Y(_18_) );
INVX1 INVX1_4 ( .A(i_add_term2[1]), .Y(_19_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term1[1]), .B(_19_), .Y(_20_) );
OAI22X1 OAI22X1_1 ( .A(_14_), .B(_16_), .C(_18_), .D(_20_), .Y(_21_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_22_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_23_) );
NOR2X1 NOR2X1_6 ( .A(_22_), .B(_23_), .Y(_24_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_25_) );
NAND2X1 NAND2X1_1 ( .A(_24_), .B(_25_), .Y(_26_) );
NOR2X1 NOR2X1_7 ( .A(_21_), .B(_26_), .Y(_3_) );
INVX1 INVX1_5 ( .A(_1_), .Y(_27_) );
NAND2X1 NAND2X1_2 ( .A(gnd), .B(_3_), .Y(_28_) );
OAI21X1 OAI21X1_1 ( .A(_3_), .B(_27_), .C(_28_), .Y(w_cout_1_) );
INVX1 INVX1_6 ( .A(i_add_term1[4]), .Y(_29_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[4]), .B(_29_), .Y(_30_) );
INVX1 INVX1_7 ( .A(i_add_term2[4]), .Y(_31_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term1[4]), .B(_31_), .Y(_32_) );
INVX1 INVX1_8 ( .A(i_add_term1[5]), .Y(_33_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[5]), .B(_33_), .Y(_34_) );
INVX1 INVX1_9 ( .A(i_add_term2[5]), .Y(_35_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term1[5]), .B(_35_), .Y(_36_) );
OAI22X1 OAI22X1_2 ( .A(_30_), .B(_32_), .C(_34_), .D(_36_), .Y(_37_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_38_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_39_) );
NOR2X1 NOR2X1_13 ( .A(_38_), .B(_39_), .Y(_40_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_41_) );
NAND2X1 NAND2X1_3 ( .A(_40_), .B(_41_), .Y(_42_) );
NOR2X1 NOR2X1_14 ( .A(_37_), .B(_42_), .Y(_6_) );
INVX1 INVX1_10 ( .A(_4_), .Y(_43_) );
NAND2X1 NAND2X1_4 ( .A(gnd), .B(_6_), .Y(_44_) );
OAI21X1 OAI21X1_2 ( .A(_6_), .B(_43_), .C(_44_), .Y(w_cout_2_) );
INVX1 INVX1_11 ( .A(i_add_term1[8]), .Y(_45_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[8]), .B(_45_), .Y(_46_) );
INVX1 INVX1_12 ( .A(i_add_term2[8]), .Y(_47_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term1[8]), .B(_47_), .Y(_48_) );
INVX1 INVX1_13 ( .A(i_add_term1[9]), .Y(_49_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[9]), .B(_49_), .Y(_50_) );
INVX1 INVX1_14 ( .A(i_add_term2[9]), .Y(_51_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term1[9]), .B(_51_), .Y(_52_) );
OAI22X1 OAI22X1_3 ( .A(_46_), .B(_48_), .C(_50_), .D(_52_), .Y(_53_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_54_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_55_) );
NOR2X1 NOR2X1_20 ( .A(_54_), .B(_55_), .Y(_56_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_57_) );
NAND2X1 NAND2X1_5 ( .A(_56_), .B(_57_), .Y(_58_) );
NOR2X1 NOR2X1_21 ( .A(_53_), .B(_58_), .Y(_9_) );
INVX1 INVX1_15 ( .A(_7_), .Y(_59_) );
NAND2X1 NAND2X1_6 ( .A(gnd), .B(_9_), .Y(_60_) );
OAI21X1 OAI21X1_3 ( .A(_9_), .B(_59_), .C(_60_), .Y(w_cout_3_) );
INVX1 INVX1_16 ( .A(i_add_term1[12]), .Y(_61_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[12]), .B(_61_), .Y(_62_) );
INVX1 INVX1_17 ( .A(i_add_term2[12]), .Y(_63_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term1[12]), .B(_63_), .Y(_64_) );
INVX1 INVX1_18 ( .A(i_add_term1[13]), .Y(_65_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[13]), .B(_65_), .Y(_66_) );
INVX1 INVX1_19 ( .A(i_add_term2[13]), .Y(_67_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term1[13]), .B(_67_), .Y(_68_) );
OAI22X1 OAI22X1_4 ( .A(_62_), .B(_64_), .C(_66_), .D(_68_), .Y(_69_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_70_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_71_) );
NOR2X1 NOR2X1_27 ( .A(_70_), .B(_71_), .Y(_72_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_73_) );
NAND2X1 NAND2X1_7 ( .A(_72_), .B(_73_), .Y(_74_) );
NOR2X1 NOR2X1_28 ( .A(_69_), .B(_74_), .Y(_12_) );
INVX1 INVX1_20 ( .A(_10_), .Y(_75_) );
NAND2X1 NAND2X1_8 ( .A(gnd), .B(_12_), .Y(_76_) );
OAI21X1 OAI21X1_4 ( .A(_12_), .B(_75_), .C(_76_), .Y(cskip2_inst_cin) );
INVX1 INVX1_21 ( .A(gnd), .Y(_80_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_81_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_82_) );
NAND3X1 NAND3X1_1 ( .A(_80_), .B(_82_), .C(_81_), .Y(_83_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_77_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_78_) );
OAI21X1 OAI21X1_5 ( .A(_77_), .B(_78_), .C(gnd), .Y(_79_) );
NAND2X1 NAND2X1_10 ( .A(_79_), .B(_83_), .Y(_0__0_) );
OAI21X1 OAI21X1_6 ( .A(_80_), .B(_77_), .C(_82_), .Y(_2__1_) );
INVX1 INVX1_22 ( .A(_2__1_), .Y(_87_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_88_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_89_) );
NAND3X1 NAND3X1_2 ( .A(_87_), .B(_89_), .C(_88_), .Y(_90_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_84_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_85_) );
OAI21X1 OAI21X1_7 ( .A(_84_), .B(_85_), .C(_2__1_), .Y(_86_) );
NAND2X1 NAND2X1_12 ( .A(_86_), .B(_90_), .Y(_0__1_) );
OAI21X1 OAI21X1_8 ( .A(_87_), .B(_84_), .C(_89_), .Y(_2__2_) );
INVX1 INVX1_23 ( .A(_2__2_), .Y(_94_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_95_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_96_) );
NAND3X1 NAND3X1_3 ( .A(_94_), .B(_96_), .C(_95_), .Y(_97_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_91_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_92_) );
OAI21X1 OAI21X1_9 ( .A(_91_), .B(_92_), .C(_2__2_), .Y(_93_) );
NAND2X1 NAND2X1_14 ( .A(_93_), .B(_97_), .Y(_0__2_) );
OAI21X1 OAI21X1_10 ( .A(_94_), .B(_91_), .C(_96_), .Y(_2__3_) );
INVX1 INVX1_24 ( .A(_2__3_), .Y(_101_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_102_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_103_) );
NAND3X1 NAND3X1_4 ( .A(_101_), .B(_103_), .C(_102_), .Y(_104_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_98_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_99_) );
OAI21X1 OAI21X1_11 ( .A(_98_), .B(_99_), .C(_2__3_), .Y(_100_) );
NAND2X1 NAND2X1_16 ( .A(_100_), .B(_104_), .Y(_0__3_) );
OAI21X1 OAI21X1_12 ( .A(_101_), .B(_98_), .C(_103_), .Y(_1_) );
INVX1 INVX1_25 ( .A(w_cout_1_), .Y(_108_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_109_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_110_) );
NAND3X1 NAND3X1_5 ( .A(_108_), .B(_110_), .C(_109_), .Y(_111_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_105_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_106_) );
OAI21X1 OAI21X1_13 ( .A(_105_), .B(_106_), .C(w_cout_1_), .Y(_107_) );
NAND2X1 NAND2X1_18 ( .A(_107_), .B(_111_), .Y(_0__4_) );
OAI21X1 OAI21X1_14 ( .A(_108_), .B(_105_), .C(_110_), .Y(_5__1_) );
INVX1 INVX1_26 ( .A(_5__1_), .Y(_115_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_116_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_117_) );
NAND3X1 NAND3X1_6 ( .A(_115_), .B(_117_), .C(_116_), .Y(_118_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_112_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_113_) );
OAI21X1 OAI21X1_15 ( .A(_112_), .B(_113_), .C(_5__1_), .Y(_114_) );
NAND2X1 NAND2X1_20 ( .A(_114_), .B(_118_), .Y(_0__5_) );
OAI21X1 OAI21X1_16 ( .A(_115_), .B(_112_), .C(_117_), .Y(_5__2_) );
INVX1 INVX1_27 ( .A(_5__2_), .Y(_122_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_123_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_124_) );
NAND3X1 NAND3X1_7 ( .A(_122_), .B(_124_), .C(_123_), .Y(_125_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_119_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_120_) );
OAI21X1 OAI21X1_17 ( .A(_119_), .B(_120_), .C(_5__2_), .Y(_121_) );
NAND2X1 NAND2X1_22 ( .A(_121_), .B(_125_), .Y(_0__6_) );
OAI21X1 OAI21X1_18 ( .A(_122_), .B(_119_), .C(_124_), .Y(_5__3_) );
INVX1 INVX1_28 ( .A(_5__3_), .Y(_129_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_130_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_131_) );
NAND3X1 NAND3X1_8 ( .A(_129_), .B(_131_), .C(_130_), .Y(_132_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_126_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_127_) );
OAI21X1 OAI21X1_19 ( .A(_126_), .B(_127_), .C(_5__3_), .Y(_128_) );
NAND2X1 NAND2X1_24 ( .A(_128_), .B(_132_), .Y(_0__7_) );
OAI21X1 OAI21X1_20 ( .A(_129_), .B(_126_), .C(_131_), .Y(_4_) );
INVX1 INVX1_29 ( .A(w_cout_2_), .Y(_136_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_137_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_138_) );
NAND3X1 NAND3X1_9 ( .A(_136_), .B(_138_), .C(_137_), .Y(_139_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_133_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_134_) );
OAI21X1 OAI21X1_21 ( .A(_133_), .B(_134_), .C(w_cout_2_), .Y(_135_) );
NAND2X1 NAND2X1_26 ( .A(_135_), .B(_139_), .Y(_0__8_) );
OAI21X1 OAI21X1_22 ( .A(_136_), .B(_133_), .C(_138_), .Y(_8__1_) );
INVX1 INVX1_30 ( .A(_8__1_), .Y(_143_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_144_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_145_) );
NAND3X1 NAND3X1_10 ( .A(_143_), .B(_145_), .C(_144_), .Y(_146_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_140_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_141_) );
OAI21X1 OAI21X1_23 ( .A(_140_), .B(_141_), .C(_8__1_), .Y(_142_) );
NAND2X1 NAND2X1_28 ( .A(_142_), .B(_146_), .Y(_0__9_) );
OAI21X1 OAI21X1_24 ( .A(_143_), .B(_140_), .C(_145_), .Y(_8__2_) );
INVX1 INVX1_31 ( .A(_8__2_), .Y(_150_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_151_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_152_) );
NAND3X1 NAND3X1_11 ( .A(_150_), .B(_152_), .C(_151_), .Y(_153_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_147_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_148_) );
OAI21X1 OAI21X1_25 ( .A(_147_), .B(_148_), .C(_8__2_), .Y(_149_) );
NAND2X1 NAND2X1_30 ( .A(_149_), .B(_153_), .Y(_0__10_) );
OAI21X1 OAI21X1_26 ( .A(_150_), .B(_147_), .C(_152_), .Y(_8__3_) );
INVX1 INVX1_32 ( .A(_8__3_), .Y(_157_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_158_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_159_) );
NAND3X1 NAND3X1_12 ( .A(_157_), .B(_159_), .C(_158_), .Y(_160_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_154_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_155_) );
OAI21X1 OAI21X1_27 ( .A(_154_), .B(_155_), .C(_8__3_), .Y(_156_) );
NAND2X1 NAND2X1_32 ( .A(_156_), .B(_160_), .Y(_0__11_) );
OAI21X1 OAI21X1_28 ( .A(_157_), .B(_154_), .C(_159_), .Y(_7_) );
INVX1 INVX1_33 ( .A(w_cout_3_), .Y(_164_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_165_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_166_) );
NAND3X1 NAND3X1_13 ( .A(_164_), .B(_166_), .C(_165_), .Y(_167_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_161_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_162_) );
OAI21X1 OAI21X1_29 ( .A(_161_), .B(_162_), .C(w_cout_3_), .Y(_163_) );
NAND2X1 NAND2X1_34 ( .A(_163_), .B(_167_), .Y(_0__12_) );
OAI21X1 OAI21X1_30 ( .A(_164_), .B(_161_), .C(_166_), .Y(_11__1_) );
INVX1 INVX1_34 ( .A(_11__1_), .Y(_171_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_172_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_173_) );
NAND3X1 NAND3X1_14 ( .A(_171_), .B(_173_), .C(_172_), .Y(_174_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_168_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_169_) );
OAI21X1 OAI21X1_31 ( .A(_168_), .B(_169_), .C(_11__1_), .Y(_170_) );
NAND2X1 NAND2X1_36 ( .A(_170_), .B(_174_), .Y(_0__13_) );
OAI21X1 OAI21X1_32 ( .A(_171_), .B(_168_), .C(_173_), .Y(_11__2_) );
INVX1 INVX1_35 ( .A(_11__2_), .Y(_178_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_179_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_180_) );
NAND3X1 NAND3X1_15 ( .A(_178_), .B(_180_), .C(_179_), .Y(_181_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_175_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_176_) );
OAI21X1 OAI21X1_33 ( .A(_175_), .B(_176_), .C(_11__2_), .Y(_177_) );
NAND2X1 NAND2X1_38 ( .A(_177_), .B(_181_), .Y(_0__14_) );
OAI21X1 OAI21X1_34 ( .A(_178_), .B(_175_), .C(_180_), .Y(_11__3_) );
INVX1 INVX1_36 ( .A(_11__3_), .Y(_185_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_186_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_187_) );
NAND3X1 NAND3X1_16 ( .A(_185_), .B(_187_), .C(_186_), .Y(_188_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_182_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_183_) );
OAI21X1 OAI21X1_35 ( .A(_182_), .B(_183_), .C(_11__3_), .Y(_184_) );
NAND2X1 NAND2X1_40 ( .A(_184_), .B(_188_), .Y(_0__15_) );
OAI21X1 OAI21X1_36 ( .A(_185_), .B(_182_), .C(_187_), .Y(_10_) );
INVX1 INVX1_37 ( .A(cskip2_inst_cin), .Y(_192_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_193_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_194_) );
NAND3X1 NAND3X1_17 ( .A(_192_), .B(_194_), .C(_193_), .Y(_195_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_189_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_190_) );
OAI21X1 OAI21X1_37 ( .A(_189_), .B(_190_), .C(cskip2_inst_cin), .Y(_191_) );
NAND2X1 NAND2X1_42 ( .A(_191_), .B(_195_), .Y(_0__16_) );
OAI21X1 OAI21X1_38 ( .A(_192_), .B(_189_), .C(_194_), .Y(cskip2_inst_rca0_w_CARRY_1_) );
INVX1 INVX1_38 ( .A(cskip2_inst_rca0_w_CARRY_1_), .Y(_199_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_200_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_201_) );
NAND3X1 NAND3X1_18 ( .A(_199_), .B(_201_), .C(_200_), .Y(_202_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_196_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_197_) );
OAI21X1 OAI21X1_39 ( .A(_196_), .B(_197_), .C(cskip2_inst_rca0_w_CARRY_1_), .Y(_198_) );
NAND2X1 NAND2X1_44 ( .A(_198_), .B(_202_), .Y(_0__17_) );
OAI21X1 OAI21X1_40 ( .A(_199_), .B(_196_), .C(_201_), .Y(cskip2_inst_rca0_w_CARRY_2_) );
INVX1 INVX1_39 ( .A(cskip2_inst_rca0_w_CARRY_2_), .Y(_204_) );
NAND2X1 NAND2X1_45 ( .A(gnd), .B(gnd), .Y(_205_) );
NOR2X1 NOR2X1_47 ( .A(gnd), .B(gnd), .Y(_203_) );
OAI21X1 OAI21X1_41 ( .A(_204_), .B(_203_), .C(_205_), .Y(cskip2_inst_rca0_w_CARRY_3_) );
INVX1 INVX1_40 ( .A(cskip2_inst_rca0_w_CARRY_3_), .Y(_207_) );
NAND2X1 NAND2X1_46 ( .A(gnd), .B(gnd), .Y(_208_) );
NOR2X1 NOR2X1_48 ( .A(gnd), .B(gnd), .Y(_206_) );
OAI21X1 OAI21X1_42 ( .A(_207_), .B(_206_), .C(_208_), .Y(cskip2_inst_cout0) );
INVX1 INVX1_41 ( .A(i_add_term1[17]), .Y(_213_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[17]), .B(_213_), .Y(_214_) );
INVX1 INVX1_42 ( .A(i_add_term2[17]), .Y(_215_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term1[17]), .B(_215_), .Y(_216_) );
INVX1 INVX1_43 ( .A(i_add_term1[16]), .Y(_209_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[16]), .B(_209_), .Y(_210_) );
INVX1 INVX1_44 ( .A(i_add_term2[16]), .Y(_211_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term1[16]), .B(_211_), .Y(_212_) );
AOI22X1 AOI22X1_1 ( .A(_214_), .B(_216_), .C(_210_), .D(_212_), .Y(cskip2_inst_skip0_P) );
INVX1 INVX1_45 ( .A(cskip2_inst_cout0), .Y(_217_) );
NAND2X1 NAND2X1_51 ( .A(gnd), .B(cskip2_inst_skip0_P), .Y(_218_) );
OAI21X1 OAI21X1_43 ( .A(cskip2_inst_skip0_P), .B(_217_), .C(_218_), .Y(w_cout_5_) );
BUFX2 BUFX2_20 ( .A(gnd), .Y(_2__0_) );
BUFX2 BUFX2_21 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_22 ( .A(w_cout_1_), .Y(_5__0_) );
BUFX2 BUFX2_23 ( .A(_4_), .Y(_5__4_) );
BUFX2 BUFX2_24 ( .A(w_cout_2_), .Y(_8__0_) );
BUFX2 BUFX2_25 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_26 ( .A(w_cout_3_), .Y(_11__0_) );
BUFX2 BUFX2_27 ( .A(_10_), .Y(_11__4_) );
BUFX2 BUFX2_28 ( .A(cskip2_inst_cin), .Y(cskip2_inst_rca0_w_CARRY_0_) );
BUFX2 BUFX2_29 ( .A(cskip2_inst_cout0), .Y(cskip2_inst_rca0_w_CARRY_4_) );
BUFX2 BUFX2_30 ( .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_31 ( .A(cskip2_inst_cin), .Y(w_cout_4_) );
endmodule
