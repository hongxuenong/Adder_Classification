module CSkipA_61bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term1[26], i_add_term1[27], i_add_term1[28], i_add_term1[29], i_add_term1[30], i_add_term1[31], i_add_term1[32], i_add_term1[33], i_add_term1[34], i_add_term1[35], i_add_term1[36], i_add_term1[37], i_add_term1[38], i_add_term1[39], i_add_term1[40], i_add_term1[41], i_add_term1[42], i_add_term1[43], i_add_term1[44], i_add_term1[45], i_add_term1[46], i_add_term1[47], i_add_term1[48], i_add_term1[49], i_add_term1[50], i_add_term1[51], i_add_term1[52], i_add_term1[53], i_add_term1[54], i_add_term1[55], i_add_term1[56], i_add_term1[57], i_add_term1[58], i_add_term1[59], i_add_term1[60], i_add_term1[61], i_add_term1[62], i_add_term1[63], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], i_add_term2[26], i_add_term2[27], i_add_term2[28], i_add_term2[29], i_add_term2[30], i_add_term2[31], i_add_term2[32], i_add_term2[33], i_add_term2[34], i_add_term2[35], i_add_term2[36], i_add_term2[37], i_add_term2[38], i_add_term2[39], i_add_term2[40], i_add_term2[41], i_add_term2[42], i_add_term2[43], i_add_term2[44], i_add_term2[45], i_add_term2[46], i_add_term2[47], i_add_term2[48], i_add_term2[49], i_add_term2[50], i_add_term2[51], i_add_term2[52], i_add_term2[53], i_add_term2[54], i_add_term2[55], i_add_term2[56], i_add_term2[57], i_add_term2[58], i_add_term2[59], i_add_term2[60], i_add_term2[61], i_add_term2[62], i_add_term2[63], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], sum[26], sum[27], sum[28], sum[29], sum[30], sum[31], sum[32], sum[33], sum[34], sum[35], sum[36], sum[37], sum[38], sum[39], sum[40], sum[41], sum[42], sum[43], sum[44], sum[45], sum[46], sum[47], sum[48], sum[49], sum[50], sum[51], sum[52], sum[53], sum[54], sum[55], sum[56], sum[57], sum[58], sum[59], sum[60], sum[61], sum[62], sum[63], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term1[26];
input i_add_term1[27];
input i_add_term1[28];
input i_add_term1[29];
input i_add_term1[30];
input i_add_term1[31];
input i_add_term1[32];
input i_add_term1[33];
input i_add_term1[34];
input i_add_term1[35];
input i_add_term1[36];
input i_add_term1[37];
input i_add_term1[38];
input i_add_term1[39];
input i_add_term1[40];
input i_add_term1[41];
input i_add_term1[42];
input i_add_term1[43];
input i_add_term1[44];
input i_add_term1[45];
input i_add_term1[46];
input i_add_term1[47];
input i_add_term1[48];
input i_add_term1[49];
input i_add_term1[50];
input i_add_term1[51];
input i_add_term1[52];
input i_add_term1[53];
input i_add_term1[54];
input i_add_term1[55];
input i_add_term1[56];
input i_add_term1[57];
input i_add_term1[58];
input i_add_term1[59];
input i_add_term1[60];
input i_add_term1[61];
input i_add_term1[62];
input i_add_term1[63];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
input i_add_term2[26];
input i_add_term2[27];
input i_add_term2[28];
input i_add_term2[29];
input i_add_term2[30];
input i_add_term2[31];
input i_add_term2[32];
input i_add_term2[33];
input i_add_term2[34];
input i_add_term2[35];
input i_add_term2[36];
input i_add_term2[37];
input i_add_term2[38];
input i_add_term2[39];
input i_add_term2[40];
input i_add_term2[41];
input i_add_term2[42];
input i_add_term2[43];
input i_add_term2[44];
input i_add_term2[45];
input i_add_term2[46];
input i_add_term2[47];
input i_add_term2[48];
input i_add_term2[49];
input i_add_term2[50];
input i_add_term2[51];
input i_add_term2[52];
input i_add_term2[53];
input i_add_term2[54];
input i_add_term2[55];
input i_add_term2[56];
input i_add_term2[57];
input i_add_term2[58];
input i_add_term2[59];
input i_add_term2[60];
input i_add_term2[61];
input i_add_term2[62];
input i_add_term2[63];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output sum[26];
output sum[27];
output sum[28];
output sum[29];
output sum[30];
output sum[31];
output sum[32];
output sum[33];
output sum[34];
output sum[35];
output sum[36];
output sum[37];
output sum[38];
output sum[39];
output sum[40];
output sum[41];
output sum[42];
output sum[43];
output sum[44];
output sum[45];
output sum[46];
output sum[47];
output sum[48];
output sum[49];
output sum[50];
output sum[51];
output sum[52];
output sum[53];
output sum[54];
output sum[55];
output sum[56];
output sum[57];
output sum[58];
output sum[59];
output sum[60];
output sum[61];
output sum[62];
output sum[63];
output cout;

NAND3X1 NAND3X1_1 ( .A(_320_), .B(_322_), .C(_321_), .Y(_323_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_317_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_318_) );
OAI21X1 OAI21X1_1 ( .A(_317_), .B(_318_), .C(w_cout_7_), .Y(_319_) );
NAND2X1 NAND2X1_1 ( .A(_319_), .B(_323_), .Y(_0__32_) );
OAI21X1 OAI21X1_2 ( .A(_320_), .B(_317_), .C(_322_), .Y(_16__1_) );
INVX1 INVX1_1 ( .A(_16__1_), .Y(_327_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_328_) );
NAND2X1 NAND2X1_2 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_329_) );
NAND3X1 NAND3X1_2 ( .A(_327_), .B(_329_), .C(_328_), .Y(_330_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_324_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_325_) );
OAI21X1 OAI21X1_3 ( .A(_324_), .B(_325_), .C(_16__1_), .Y(_326_) );
NAND2X1 NAND2X1_3 ( .A(_326_), .B(_330_), .Y(_0__33_) );
OAI21X1 OAI21X1_4 ( .A(_327_), .B(_324_), .C(_329_), .Y(_16__2_) );
INVX1 INVX1_2 ( .A(_16__2_), .Y(_334_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_335_) );
NAND2X1 NAND2X1_4 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_336_) );
NAND3X1 NAND3X1_3 ( .A(_334_), .B(_336_), .C(_335_), .Y(_337_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_331_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_332_) );
OAI21X1 OAI21X1_5 ( .A(_331_), .B(_332_), .C(_16__2_), .Y(_333_) );
NAND2X1 NAND2X1_5 ( .A(_333_), .B(_337_), .Y(_0__34_) );
OAI21X1 OAI21X1_6 ( .A(_334_), .B(_331_), .C(_336_), .Y(_16__3_) );
INVX1 INVX1_3 ( .A(_16__3_), .Y(_341_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_342_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_343_) );
NAND3X1 NAND3X1_4 ( .A(_341_), .B(_343_), .C(_342_), .Y(_344_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_338_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_339_) );
OAI21X1 OAI21X1_7 ( .A(_338_), .B(_339_), .C(_16__3_), .Y(_340_) );
NAND2X1 NAND2X1_7 ( .A(_340_), .B(_344_), .Y(_0__35_) );
OAI21X1 OAI21X1_8 ( .A(_341_), .B(_338_), .C(_343_), .Y(_15_) );
INVX1 INVX1_4 ( .A(w_cout_8_), .Y(_348_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_349_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_350_) );
NAND3X1 NAND3X1_5 ( .A(_348_), .B(_350_), .C(_349_), .Y(_351_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_345_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_346_) );
OAI21X1 OAI21X1_9 ( .A(_345_), .B(_346_), .C(w_cout_8_), .Y(_347_) );
NAND2X1 NAND2X1_9 ( .A(_347_), .B(_351_), .Y(_0__36_) );
OAI21X1 OAI21X1_10 ( .A(_348_), .B(_345_), .C(_350_), .Y(_18__1_) );
INVX1 INVX1_5 ( .A(_18__1_), .Y(_355_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_356_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_357_) );
NAND3X1 NAND3X1_6 ( .A(_355_), .B(_357_), .C(_356_), .Y(_358_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_352_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_353_) );
OAI21X1 OAI21X1_11 ( .A(_352_), .B(_353_), .C(_18__1_), .Y(_354_) );
NAND2X1 NAND2X1_11 ( .A(_354_), .B(_358_), .Y(_0__37_) );
OAI21X1 OAI21X1_12 ( .A(_355_), .B(_352_), .C(_357_), .Y(_18__2_) );
INVX1 INVX1_6 ( .A(_18__2_), .Y(_362_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_363_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_364_) );
NAND3X1 NAND3X1_7 ( .A(_362_), .B(_364_), .C(_363_), .Y(_365_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_359_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_360_) );
OAI21X1 OAI21X1_13 ( .A(_359_), .B(_360_), .C(_18__2_), .Y(_361_) );
NAND2X1 NAND2X1_13 ( .A(_361_), .B(_365_), .Y(_0__38_) );
OAI21X1 OAI21X1_14 ( .A(_362_), .B(_359_), .C(_364_), .Y(_18__3_) );
INVX1 INVX1_7 ( .A(_18__3_), .Y(_369_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_370_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_371_) );
NAND3X1 NAND3X1_8 ( .A(_369_), .B(_371_), .C(_370_), .Y(_372_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_366_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_367_) );
OAI21X1 OAI21X1_15 ( .A(_366_), .B(_367_), .C(_18__3_), .Y(_368_) );
NAND2X1 NAND2X1_15 ( .A(_368_), .B(_372_), .Y(_0__39_) );
OAI21X1 OAI21X1_16 ( .A(_369_), .B(_366_), .C(_371_), .Y(_17_) );
INVX1 INVX1_8 ( .A(w_cout_9_), .Y(_376_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_377_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_378_) );
NAND3X1 NAND3X1_9 ( .A(_376_), .B(_378_), .C(_377_), .Y(_379_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_373_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_374_) );
OAI21X1 OAI21X1_17 ( .A(_373_), .B(_374_), .C(w_cout_9_), .Y(_375_) );
NAND2X1 NAND2X1_17 ( .A(_375_), .B(_379_), .Y(_0__40_) );
OAI21X1 OAI21X1_18 ( .A(_376_), .B(_373_), .C(_378_), .Y(_20__1_) );
INVX1 INVX1_9 ( .A(_20__1_), .Y(_383_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_384_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_385_) );
NAND3X1 NAND3X1_10 ( .A(_383_), .B(_385_), .C(_384_), .Y(_386_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_380_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_381_) );
OAI21X1 OAI21X1_19 ( .A(_380_), .B(_381_), .C(_20__1_), .Y(_382_) );
NAND2X1 NAND2X1_19 ( .A(_382_), .B(_386_), .Y(_0__41_) );
OAI21X1 OAI21X1_20 ( .A(_383_), .B(_380_), .C(_385_), .Y(_20__2_) );
INVX1 INVX1_10 ( .A(_20__2_), .Y(_390_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_391_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_392_) );
NAND3X1 NAND3X1_11 ( .A(_390_), .B(_392_), .C(_391_), .Y(_393_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_387_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_388_) );
OAI21X1 OAI21X1_21 ( .A(_387_), .B(_388_), .C(_20__2_), .Y(_389_) );
NAND2X1 NAND2X1_21 ( .A(_389_), .B(_393_), .Y(_0__42_) );
OAI21X1 OAI21X1_22 ( .A(_390_), .B(_387_), .C(_392_), .Y(_20__3_) );
INVX1 INVX1_11 ( .A(_20__3_), .Y(_397_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_398_) );
NAND2X1 NAND2X1_22 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_399_) );
NAND3X1 NAND3X1_12 ( .A(_397_), .B(_399_), .C(_398_), .Y(_400_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_394_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_395_) );
OAI21X1 OAI21X1_23 ( .A(_394_), .B(_395_), .C(_20__3_), .Y(_396_) );
NAND2X1 NAND2X1_23 ( .A(_396_), .B(_400_), .Y(_0__43_) );
OAI21X1 OAI21X1_24 ( .A(_397_), .B(_394_), .C(_399_), .Y(_19_) );
INVX1 INVX1_12 ( .A(w_cout_10_), .Y(_404_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_405_) );
NAND2X1 NAND2X1_24 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_406_) );
NAND3X1 NAND3X1_13 ( .A(_404_), .B(_406_), .C(_405_), .Y(_407_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_401_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_402_) );
OAI21X1 OAI21X1_25 ( .A(_401_), .B(_402_), .C(w_cout_10_), .Y(_403_) );
NAND2X1 NAND2X1_25 ( .A(_403_), .B(_407_), .Y(_0__44_) );
OAI21X1 OAI21X1_26 ( .A(_404_), .B(_401_), .C(_406_), .Y(_22__1_) );
INVX1 INVX1_13 ( .A(_22__1_), .Y(_411_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_412_) );
NAND2X1 NAND2X1_26 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_413_) );
NAND3X1 NAND3X1_14 ( .A(_411_), .B(_413_), .C(_412_), .Y(_414_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_408_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_409_) );
OAI21X1 OAI21X1_27 ( .A(_408_), .B(_409_), .C(_22__1_), .Y(_410_) );
NAND2X1 NAND2X1_27 ( .A(_410_), .B(_414_), .Y(_0__45_) );
OAI21X1 OAI21X1_28 ( .A(_411_), .B(_408_), .C(_413_), .Y(_22__2_) );
INVX1 INVX1_14 ( .A(_22__2_), .Y(_418_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_419_) );
NAND2X1 NAND2X1_28 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_420_) );
NAND3X1 NAND3X1_15 ( .A(_418_), .B(_420_), .C(_419_), .Y(_421_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_415_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_416_) );
OAI21X1 OAI21X1_29 ( .A(_415_), .B(_416_), .C(_22__2_), .Y(_417_) );
NAND2X1 NAND2X1_29 ( .A(_417_), .B(_421_), .Y(_0__46_) );
OAI21X1 OAI21X1_30 ( .A(_418_), .B(_415_), .C(_420_), .Y(_22__3_) );
INVX1 INVX1_15 ( .A(_22__3_), .Y(_425_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_426_) );
NAND2X1 NAND2X1_30 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_427_) );
NAND3X1 NAND3X1_16 ( .A(_425_), .B(_427_), .C(_426_), .Y(_428_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_422_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_423_) );
OAI21X1 OAI21X1_31 ( .A(_422_), .B(_423_), .C(_22__3_), .Y(_424_) );
NAND2X1 NAND2X1_31 ( .A(_424_), .B(_428_), .Y(_0__47_) );
OAI21X1 OAI21X1_32 ( .A(_425_), .B(_422_), .C(_427_), .Y(_21_) );
INVX1 INVX1_16 ( .A(w_cout_11_), .Y(_432_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_433_) );
NAND2X1 NAND2X1_32 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_434_) );
NAND3X1 NAND3X1_17 ( .A(_432_), .B(_434_), .C(_433_), .Y(_435_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_429_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_430_) );
OAI21X1 OAI21X1_33 ( .A(_429_), .B(_430_), .C(w_cout_11_), .Y(_431_) );
NAND2X1 NAND2X1_33 ( .A(_431_), .B(_435_), .Y(_0__48_) );
OAI21X1 OAI21X1_34 ( .A(_432_), .B(_429_), .C(_434_), .Y(_24__1_) );
INVX1 INVX1_17 ( .A(_24__1_), .Y(_439_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_440_) );
NAND2X1 NAND2X1_34 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_441_) );
NAND3X1 NAND3X1_18 ( .A(_439_), .B(_441_), .C(_440_), .Y(_442_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_436_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_437_) );
OAI21X1 OAI21X1_35 ( .A(_436_), .B(_437_), .C(_24__1_), .Y(_438_) );
NAND2X1 NAND2X1_35 ( .A(_438_), .B(_442_), .Y(_0__49_) );
OAI21X1 OAI21X1_36 ( .A(_439_), .B(_436_), .C(_441_), .Y(_24__2_) );
INVX1 INVX1_18 ( .A(_24__2_), .Y(_446_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_447_) );
NAND2X1 NAND2X1_36 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_448_) );
NAND3X1 NAND3X1_19 ( .A(_446_), .B(_448_), .C(_447_), .Y(_449_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_443_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_444_) );
OAI21X1 OAI21X1_37 ( .A(_443_), .B(_444_), .C(_24__2_), .Y(_445_) );
NAND2X1 NAND2X1_37 ( .A(_445_), .B(_449_), .Y(_0__50_) );
OAI21X1 OAI21X1_38 ( .A(_446_), .B(_443_), .C(_448_), .Y(_24__3_) );
INVX1 INVX1_19 ( .A(_24__3_), .Y(_453_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_454_) );
NAND2X1 NAND2X1_38 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_455_) );
NAND3X1 NAND3X1_20 ( .A(_453_), .B(_455_), .C(_454_), .Y(_456_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_450_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_451_) );
OAI21X1 OAI21X1_39 ( .A(_450_), .B(_451_), .C(_24__3_), .Y(_452_) );
NAND2X1 NAND2X1_39 ( .A(_452_), .B(_456_), .Y(_0__51_) );
OAI21X1 OAI21X1_40 ( .A(_453_), .B(_450_), .C(_455_), .Y(_23_) );
INVX1 INVX1_20 ( .A(w_cout_12_), .Y(_460_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_461_) );
NAND2X1 NAND2X1_40 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_462_) );
NAND3X1 NAND3X1_21 ( .A(_460_), .B(_462_), .C(_461_), .Y(_463_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_457_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_458_) );
OAI21X1 OAI21X1_41 ( .A(_457_), .B(_458_), .C(w_cout_12_), .Y(_459_) );
NAND2X1 NAND2X1_41 ( .A(_459_), .B(_463_), .Y(_0__52_) );
OAI21X1 OAI21X1_42 ( .A(_460_), .B(_457_), .C(_462_), .Y(_26__1_) );
INVX1 INVX1_21 ( .A(_26__1_), .Y(_467_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_468_) );
NAND2X1 NAND2X1_42 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_469_) );
NAND3X1 NAND3X1_22 ( .A(_467_), .B(_469_), .C(_468_), .Y(_470_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_464_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_465_) );
OAI21X1 OAI21X1_43 ( .A(_464_), .B(_465_), .C(_26__1_), .Y(_466_) );
NAND2X1 NAND2X1_43 ( .A(_466_), .B(_470_), .Y(_0__53_) );
OAI21X1 OAI21X1_44 ( .A(_467_), .B(_464_), .C(_469_), .Y(_26__2_) );
INVX1 INVX1_22 ( .A(_26__2_), .Y(_474_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_475_) );
NAND2X1 NAND2X1_44 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_476_) );
NAND3X1 NAND3X1_23 ( .A(_474_), .B(_476_), .C(_475_), .Y(_477_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_471_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_472_) );
OAI21X1 OAI21X1_45 ( .A(_471_), .B(_472_), .C(_26__2_), .Y(_473_) );
NAND2X1 NAND2X1_45 ( .A(_473_), .B(_477_), .Y(_0__54_) );
OAI21X1 OAI21X1_46 ( .A(_474_), .B(_471_), .C(_476_), .Y(_26__3_) );
INVX1 INVX1_23 ( .A(_26__3_), .Y(_481_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_482_) );
NAND2X1 NAND2X1_46 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_483_) );
NAND3X1 NAND3X1_24 ( .A(_481_), .B(_483_), .C(_482_), .Y(_484_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_478_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_479_) );
OAI21X1 OAI21X1_47 ( .A(_478_), .B(_479_), .C(_26__3_), .Y(_480_) );
NAND2X1 NAND2X1_47 ( .A(_480_), .B(_484_), .Y(_0__55_) );
OAI21X1 OAI21X1_48 ( .A(_481_), .B(_478_), .C(_483_), .Y(_25_) );
INVX1 INVX1_24 ( .A(w_cout_13_), .Y(_488_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_489_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_490_) );
NAND3X1 NAND3X1_25 ( .A(_488_), .B(_490_), .C(_489_), .Y(_491_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_485_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_486_) );
OAI21X1 OAI21X1_49 ( .A(_485_), .B(_486_), .C(w_cout_13_), .Y(_487_) );
NAND2X1 NAND2X1_49 ( .A(_487_), .B(_491_), .Y(_0__56_) );
OAI21X1 OAI21X1_50 ( .A(_488_), .B(_485_), .C(_490_), .Y(_28__1_) );
INVX1 INVX1_25 ( .A(_28__1_), .Y(_495_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_496_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_497_) );
NAND3X1 NAND3X1_26 ( .A(_495_), .B(_497_), .C(_496_), .Y(_498_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_492_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_493_) );
OAI21X1 OAI21X1_51 ( .A(_492_), .B(_493_), .C(_28__1_), .Y(_494_) );
NAND2X1 NAND2X1_51 ( .A(_494_), .B(_498_), .Y(_0__57_) );
OAI21X1 OAI21X1_52 ( .A(_495_), .B(_492_), .C(_497_), .Y(_28__2_) );
INVX1 INVX1_26 ( .A(_28__2_), .Y(_502_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_503_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_504_) );
NAND3X1 NAND3X1_27 ( .A(_502_), .B(_504_), .C(_503_), .Y(_505_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_499_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_500_) );
OAI21X1 OAI21X1_53 ( .A(_499_), .B(_500_), .C(_28__2_), .Y(_501_) );
NAND2X1 NAND2X1_53 ( .A(_501_), .B(_505_), .Y(_0__58_) );
OAI21X1 OAI21X1_54 ( .A(_502_), .B(_499_), .C(_504_), .Y(_28__3_) );
INVX1 INVX1_27 ( .A(_28__3_), .Y(_509_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_510_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_511_) );
NAND3X1 NAND3X1_28 ( .A(_509_), .B(_511_), .C(_510_), .Y(_512_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_506_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_507_) );
OAI21X1 OAI21X1_55 ( .A(_506_), .B(_507_), .C(_28__3_), .Y(_508_) );
NAND2X1 NAND2X1_55 ( .A(_508_), .B(_512_), .Y(_0__59_) );
OAI21X1 OAI21X1_56 ( .A(_509_), .B(_506_), .C(_511_), .Y(_27_) );
INVX1 INVX1_28 ( .A(w_cout_14_), .Y(_516_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_517_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_518_) );
NAND3X1 NAND3X1_29 ( .A(_516_), .B(_518_), .C(_517_), .Y(_519_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_513_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .Y(_514_) );
OAI21X1 OAI21X1_57 ( .A(_513_), .B(_514_), .C(w_cout_14_), .Y(_515_) );
NAND2X1 NAND2X1_57 ( .A(_515_), .B(_519_), .Y(_0__60_) );
OAI21X1 OAI21X1_58 ( .A(_516_), .B(_513_), .C(_518_), .Y(_30__1_) );
INVX1 INVX1_29 ( .A(_30__1_), .Y(_523_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_524_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_525_) );
NAND3X1 NAND3X1_30 ( .A(_523_), .B(_525_), .C(_524_), .Y(_526_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_520_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_521_) );
OAI21X1 OAI21X1_59 ( .A(_520_), .B(_521_), .C(_30__1_), .Y(_522_) );
NAND2X1 NAND2X1_59 ( .A(_522_), .B(_526_), .Y(_0__61_) );
OAI21X1 OAI21X1_60 ( .A(_523_), .B(_520_), .C(_525_), .Y(_30__2_) );
INVX1 INVX1_30 ( .A(_30__2_), .Y(_530_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_531_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_532_) );
NAND3X1 NAND3X1_31 ( .A(_530_), .B(_532_), .C(_531_), .Y(_533_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_527_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_528_) );
OAI21X1 OAI21X1_61 ( .A(_527_), .B(_528_), .C(_30__2_), .Y(_529_) );
NAND2X1 NAND2X1_61 ( .A(_529_), .B(_533_), .Y(_0__62_) );
OAI21X1 OAI21X1_62 ( .A(_530_), .B(_527_), .C(_532_), .Y(_30__3_) );
INVX1 INVX1_31 ( .A(_30__3_), .Y(_537_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_538_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_539_) );
NAND3X1 NAND3X1_32 ( .A(_537_), .B(_539_), .C(_538_), .Y(_540_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_534_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_535_) );
OAI21X1 OAI21X1_63 ( .A(_534_), .B(_535_), .C(_30__3_), .Y(_536_) );
NAND2X1 NAND2X1_63 ( .A(_536_), .B(_540_), .Y(_0__63_) );
OAI21X1 OAI21X1_64 ( .A(_537_), .B(_534_), .C(_539_), .Y(_29_) );
INVX1 INVX1_32 ( .A(1'b0), .Y(_544_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_545_) );
NAND2X1 NAND2X1_64 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_546_) );
NAND3X1 NAND3X1_33 ( .A(_544_), .B(_546_), .C(_545_), .Y(_547_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_541_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_542_) );
OAI21X1 OAI21X1_65 ( .A(_541_), .B(_542_), .C(1'b0), .Y(_543_) );
NAND2X1 NAND2X1_65 ( .A(_543_), .B(_547_), .Y(_0__0_) );
OAI21X1 OAI21X1_66 ( .A(_544_), .B(_541_), .C(_546_), .Y(rca_inst_w_CARRY_1_) );
INVX1 INVX1_33 ( .A(rca_inst_w_CARRY_1_), .Y(_551_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_552_) );
NAND2X1 NAND2X1_66 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_553_) );
NAND3X1 NAND3X1_34 ( .A(_551_), .B(_553_), .C(_552_), .Y(_554_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_548_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_549_) );
OAI21X1 OAI21X1_67 ( .A(_548_), .B(_549_), .C(rca_inst_w_CARRY_1_), .Y(_550_) );
NAND2X1 NAND2X1_67 ( .A(_550_), .B(_554_), .Y(_0__1_) );
OAI21X1 OAI21X1_68 ( .A(_551_), .B(_548_), .C(_553_), .Y(rca_inst_w_CARRY_2_) );
INVX1 INVX1_34 ( .A(rca_inst_w_CARRY_2_), .Y(_558_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_559_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_560_) );
NAND3X1 NAND3X1_35 ( .A(_558_), .B(_560_), .C(_559_), .Y(_561_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_555_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_556_) );
OAI21X1 OAI21X1_69 ( .A(_555_), .B(_556_), .C(rca_inst_w_CARRY_2_), .Y(_557_) );
NAND2X1 NAND2X1_69 ( .A(_557_), .B(_561_), .Y(_0__2_) );
OAI21X1 OAI21X1_70 ( .A(_558_), .B(_555_), .C(_560_), .Y(rca_inst_w_CARRY_3_) );
INVX1 INVX1_35 ( .A(rca_inst_w_CARRY_3_), .Y(_565_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_566_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_567_) );
NAND3X1 NAND3X1_36 ( .A(_565_), .B(_567_), .C(_566_), .Y(_568_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_562_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_563_) );
OAI21X1 OAI21X1_71 ( .A(_562_), .B(_563_), .C(rca_inst_w_CARRY_3_), .Y(_564_) );
NAND2X1 NAND2X1_71 ( .A(_564_), .B(_568_), .Y(_0__3_) );
OAI21X1 OAI21X1_72 ( .A(_565_), .B(_562_), .C(_567_), .Y(cout0) );
INVX1 INVX1_36 ( .A(cout0), .Y(_569_) );
OAI21X1 OAI21X1_73 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .C(1'b0), .Y(_570_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_571_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_572_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_573_) );
NAND3X1 NAND3X1_37 ( .A(_571_), .B(_572_), .C(_573_), .Y(_574_) );
OAI21X1 OAI21X1_74 ( .A(_570_), .B(_574_), .C(_569_), .Y(skip0_cin_next) );
BUFX2 BUFX2_1 ( .A(w_cout_15_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .A(_0__54_), .Y(sum[54]) );
BUFX2 BUFX2_57 ( .A(_0__55_), .Y(sum[55]) );
BUFX2 BUFX2_58 ( .A(_0__56_), .Y(sum[56]) );
BUFX2 BUFX2_59 ( .A(_0__57_), .Y(sum[57]) );
BUFX2 BUFX2_60 ( .A(_0__58_), .Y(sum[58]) );
BUFX2 BUFX2_61 ( .A(_0__59_), .Y(sum[59]) );
BUFX2 BUFX2_62 ( .A(_0__60_), .Y(sum[60]) );
BUFX2 BUFX2_63 ( .A(_0__61_), .Y(sum[61]) );
BUFX2 BUFX2_64 ( .A(_0__62_), .Y(sum[62]) );
BUFX2 BUFX2_65 ( .A(_0__63_), .Y(sum[63]) );
INVX1 INVX1_37 ( .A(_1_), .Y(_31_) );
OAI21X1 OAI21X1_75 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .C(1'b0), .Y(_32_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_33_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_34_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_35_) );
NAND3X1 NAND3X1_38 ( .A(_33_), .B(_34_), .C(_35_), .Y(_36_) );
OAI21X1 OAI21X1_76 ( .A(_32_), .B(_36_), .C(_31_), .Y(w_cout_1_) );
INVX1 INVX1_38 ( .A(_3_), .Y(_37_) );
OAI21X1 OAI21X1_77 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .C(1'b0), .Y(_38_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_39_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_40_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_41_) );
NAND3X1 NAND3X1_39 ( .A(_39_), .B(_40_), .C(_41_), .Y(_42_) );
OAI21X1 OAI21X1_78 ( .A(_38_), .B(_42_), .C(_37_), .Y(w_cout_2_) );
INVX1 INVX1_39 ( .A(_5_), .Y(_43_) );
OAI21X1 OAI21X1_79 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .C(1'b0), .Y(_44_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_45_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_46_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_47_) );
NAND3X1 NAND3X1_40 ( .A(_45_), .B(_46_), .C(_47_), .Y(_48_) );
OAI21X1 OAI21X1_80 ( .A(_44_), .B(_48_), .C(_43_), .Y(w_cout_3_) );
INVX1 INVX1_40 ( .A(_7_), .Y(_49_) );
OAI21X1 OAI21X1_81 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .C(1'b0), .Y(_50_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_51_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_52_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_53_) );
NAND3X1 NAND3X1_41 ( .A(_51_), .B(_52_), .C(_53_), .Y(_54_) );
OAI21X1 OAI21X1_82 ( .A(_50_), .B(_54_), .C(_49_), .Y(w_cout_4_) );
INVX1 INVX1_41 ( .A(_9_), .Y(_55_) );
OAI21X1 OAI21X1_83 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .C(1'b0), .Y(_56_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_57_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_58_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_59_) );
NAND3X1 NAND3X1_42 ( .A(_57_), .B(_58_), .C(_59_), .Y(_60_) );
OAI21X1 OAI21X1_84 ( .A(_56_), .B(_60_), .C(_55_), .Y(w_cout_5_) );
INVX1 INVX1_42 ( .A(_11_), .Y(_61_) );
OAI21X1 OAI21X1_85 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .C(1'b0), .Y(_62_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_63_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_64_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_65_) );
NAND3X1 NAND3X1_43 ( .A(_63_), .B(_64_), .C(_65_), .Y(_66_) );
OAI21X1 OAI21X1_86 ( .A(_62_), .B(_66_), .C(_61_), .Y(w_cout_6_) );
INVX1 INVX1_43 ( .A(_13_), .Y(_67_) );
OAI21X1 OAI21X1_87 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .C(1'b0), .Y(_68_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_69_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_70_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_71_) );
NAND3X1 NAND3X1_44 ( .A(_69_), .B(_70_), .C(_71_), .Y(_72_) );
OAI21X1 OAI21X1_88 ( .A(_68_), .B(_72_), .C(_67_), .Y(w_cout_7_) );
INVX1 INVX1_44 ( .A(_15_), .Y(_73_) );
OAI21X1 OAI21X1_89 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .C(1'b0), .Y(_74_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_75_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_76_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_77_) );
NAND3X1 NAND3X1_45 ( .A(_75_), .B(_76_), .C(_77_), .Y(_78_) );
OAI21X1 OAI21X1_90 ( .A(_74_), .B(_78_), .C(_73_), .Y(w_cout_8_) );
INVX1 INVX1_45 ( .A(_17_), .Y(_79_) );
OAI21X1 OAI21X1_91 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .C(1'b0), .Y(_80_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_81_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_82_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_83_) );
NAND3X1 NAND3X1_46 ( .A(_81_), .B(_82_), .C(_83_), .Y(_84_) );
OAI21X1 OAI21X1_92 ( .A(_80_), .B(_84_), .C(_79_), .Y(w_cout_9_) );
INVX1 INVX1_46 ( .A(_19_), .Y(_85_) );
OAI21X1 OAI21X1_93 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .C(1'b0), .Y(_86_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_87_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_88_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_89_) );
NAND3X1 NAND3X1_47 ( .A(_87_), .B(_88_), .C(_89_), .Y(_90_) );
OAI21X1 OAI21X1_94 ( .A(_86_), .B(_90_), .C(_85_), .Y(w_cout_10_) );
INVX1 INVX1_47 ( .A(_21_), .Y(_91_) );
OAI21X1 OAI21X1_95 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .C(1'b0), .Y(_92_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_93_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_94_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_95_) );
NAND3X1 NAND3X1_48 ( .A(_93_), .B(_94_), .C(_95_), .Y(_96_) );
OAI21X1 OAI21X1_96 ( .A(_92_), .B(_96_), .C(_91_), .Y(w_cout_11_) );
INVX1 INVX1_48 ( .A(_23_), .Y(_97_) );
OAI21X1 OAI21X1_97 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .C(1'b0), .Y(_98_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_99_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_100_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_101_) );
NAND3X1 NAND3X1_49 ( .A(_99_), .B(_100_), .C(_101_), .Y(_102_) );
OAI21X1 OAI21X1_98 ( .A(_98_), .B(_102_), .C(_97_), .Y(w_cout_12_) );
INVX1 INVX1_49 ( .A(_25_), .Y(_103_) );
OAI21X1 OAI21X1_99 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .C(1'b0), .Y(_104_) );
OR2X2 OR2X2_75 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_105_) );
OR2X2 OR2X2_76 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_106_) );
OR2X2 OR2X2_77 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_107_) );
NAND3X1 NAND3X1_50 ( .A(_105_), .B(_106_), .C(_107_), .Y(_108_) );
OAI21X1 OAI21X1_100 ( .A(_104_), .B(_108_), .C(_103_), .Y(w_cout_13_) );
INVX1 INVX1_50 ( .A(_27_), .Y(_109_) );
OAI21X1 OAI21X1_101 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .C(1'b0), .Y(_110_) );
OR2X2 OR2X2_78 ( .A(i_add_term2[59]), .B(i_add_term1[59]), .Y(_111_) );
OR2X2 OR2X2_79 ( .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_112_) );
OR2X2 OR2X2_80 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_113_) );
NAND3X1 NAND3X1_51 ( .A(_111_), .B(_112_), .C(_113_), .Y(_114_) );
OAI21X1 OAI21X1_102 ( .A(_110_), .B(_114_), .C(_109_), .Y(w_cout_14_) );
INVX1 INVX1_51 ( .A(_29_), .Y(_115_) );
OAI21X1 OAI21X1_103 ( .A(i_add_term2[60]), .B(i_add_term1[60]), .C(1'b0), .Y(_116_) );
OR2X2 OR2X2_81 ( .A(i_add_term2[63]), .B(i_add_term1[63]), .Y(_117_) );
OR2X2 OR2X2_82 ( .A(i_add_term2[62]), .B(i_add_term1[62]), .Y(_118_) );
OR2X2 OR2X2_83 ( .A(i_add_term2[61]), .B(i_add_term1[61]), .Y(_119_) );
NAND3X1 NAND3X1_52 ( .A(_117_), .B(_118_), .C(_119_), .Y(_120_) );
OAI21X1 OAI21X1_104 ( .A(_116_), .B(_120_), .C(_115_), .Y(w_cout_15_) );
INVX1 INVX1_52 ( .A(skip0_cin_next), .Y(_124_) );
OR2X2 OR2X2_84 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_125_) );
NAND2X1 NAND2X1_72 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_126_) );
NAND3X1 NAND3X1_53 ( .A(_124_), .B(_126_), .C(_125_), .Y(_127_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_121_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_122_) );
OAI21X1 OAI21X1_105 ( .A(_121_), .B(_122_), .C(skip0_cin_next), .Y(_123_) );
NAND2X1 NAND2X1_73 ( .A(_123_), .B(_127_), .Y(_0__4_) );
OAI21X1 OAI21X1_106 ( .A(_124_), .B(_121_), .C(_126_), .Y(_2__1_) );
INVX1 INVX1_53 ( .A(_2__1_), .Y(_131_) );
OR2X2 OR2X2_85 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_132_) );
NAND2X1 NAND2X1_74 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_133_) );
NAND3X1 NAND3X1_54 ( .A(_131_), .B(_133_), .C(_132_), .Y(_134_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_128_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_129_) );
OAI21X1 OAI21X1_107 ( .A(_128_), .B(_129_), .C(_2__1_), .Y(_130_) );
NAND2X1 NAND2X1_75 ( .A(_130_), .B(_134_), .Y(_0__5_) );
OAI21X1 OAI21X1_108 ( .A(_131_), .B(_128_), .C(_133_), .Y(_2__2_) );
INVX1 INVX1_54 ( .A(_2__2_), .Y(_138_) );
OR2X2 OR2X2_86 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_139_) );
NAND2X1 NAND2X1_76 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_140_) );
NAND3X1 NAND3X1_55 ( .A(_138_), .B(_140_), .C(_139_), .Y(_141_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_135_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_136_) );
OAI21X1 OAI21X1_109 ( .A(_135_), .B(_136_), .C(_2__2_), .Y(_137_) );
NAND2X1 NAND2X1_77 ( .A(_137_), .B(_141_), .Y(_0__6_) );
OAI21X1 OAI21X1_110 ( .A(_138_), .B(_135_), .C(_140_), .Y(_2__3_) );
INVX1 INVX1_55 ( .A(_2__3_), .Y(_145_) );
OR2X2 OR2X2_87 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_146_) );
NAND2X1 NAND2X1_78 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_147_) );
NAND3X1 NAND3X1_56 ( .A(_145_), .B(_147_), .C(_146_), .Y(_148_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_142_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_143_) );
OAI21X1 OAI21X1_111 ( .A(_142_), .B(_143_), .C(_2__3_), .Y(_144_) );
NAND2X1 NAND2X1_79 ( .A(_144_), .B(_148_), .Y(_0__7_) );
OAI21X1 OAI21X1_112 ( .A(_145_), .B(_142_), .C(_147_), .Y(_1_) );
INVX1 INVX1_56 ( .A(w_cout_1_), .Y(_152_) );
OR2X2 OR2X2_88 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_153_) );
NAND2X1 NAND2X1_80 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_154_) );
NAND3X1 NAND3X1_57 ( .A(_152_), .B(_154_), .C(_153_), .Y(_155_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_149_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_150_) );
OAI21X1 OAI21X1_113 ( .A(_149_), .B(_150_), .C(w_cout_1_), .Y(_151_) );
NAND2X1 NAND2X1_81 ( .A(_151_), .B(_155_), .Y(_0__8_) );
OAI21X1 OAI21X1_114 ( .A(_152_), .B(_149_), .C(_154_), .Y(_4__1_) );
INVX1 INVX1_57 ( .A(_4__1_), .Y(_159_) );
OR2X2 OR2X2_89 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_160_) );
NAND2X1 NAND2X1_82 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_161_) );
NAND3X1 NAND3X1_58 ( .A(_159_), .B(_161_), .C(_160_), .Y(_162_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_156_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_157_) );
OAI21X1 OAI21X1_115 ( .A(_156_), .B(_157_), .C(_4__1_), .Y(_158_) );
NAND2X1 NAND2X1_83 ( .A(_158_), .B(_162_), .Y(_0__9_) );
OAI21X1 OAI21X1_116 ( .A(_159_), .B(_156_), .C(_161_), .Y(_4__2_) );
INVX1 INVX1_58 ( .A(_4__2_), .Y(_166_) );
OR2X2 OR2X2_90 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_167_) );
NAND2X1 NAND2X1_84 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_168_) );
NAND3X1 NAND3X1_59 ( .A(_166_), .B(_168_), .C(_167_), .Y(_169_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_163_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_164_) );
OAI21X1 OAI21X1_117 ( .A(_163_), .B(_164_), .C(_4__2_), .Y(_165_) );
NAND2X1 NAND2X1_85 ( .A(_165_), .B(_169_), .Y(_0__10_) );
OAI21X1 OAI21X1_118 ( .A(_166_), .B(_163_), .C(_168_), .Y(_4__3_) );
INVX1 INVX1_59 ( .A(_4__3_), .Y(_173_) );
OR2X2 OR2X2_91 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_174_) );
NAND2X1 NAND2X1_86 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_175_) );
NAND3X1 NAND3X1_60 ( .A(_173_), .B(_175_), .C(_174_), .Y(_176_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_170_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_171_) );
OAI21X1 OAI21X1_119 ( .A(_170_), .B(_171_), .C(_4__3_), .Y(_172_) );
NAND2X1 NAND2X1_87 ( .A(_172_), .B(_176_), .Y(_0__11_) );
OAI21X1 OAI21X1_120 ( .A(_173_), .B(_170_), .C(_175_), .Y(_3_) );
INVX1 INVX1_60 ( .A(w_cout_2_), .Y(_180_) );
OR2X2 OR2X2_92 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_181_) );
NAND2X1 NAND2X1_88 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_182_) );
NAND3X1 NAND3X1_61 ( .A(_180_), .B(_182_), .C(_181_), .Y(_183_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_177_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_178_) );
OAI21X1 OAI21X1_121 ( .A(_177_), .B(_178_), .C(w_cout_2_), .Y(_179_) );
NAND2X1 NAND2X1_89 ( .A(_179_), .B(_183_), .Y(_0__12_) );
OAI21X1 OAI21X1_122 ( .A(_180_), .B(_177_), .C(_182_), .Y(_6__1_) );
INVX1 INVX1_61 ( .A(_6__1_), .Y(_187_) );
OR2X2 OR2X2_93 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_188_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_189_) );
NAND3X1 NAND3X1_62 ( .A(_187_), .B(_189_), .C(_188_), .Y(_190_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_184_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_185_) );
OAI21X1 OAI21X1_123 ( .A(_184_), .B(_185_), .C(_6__1_), .Y(_186_) );
NAND2X1 NAND2X1_91 ( .A(_186_), .B(_190_), .Y(_0__13_) );
OAI21X1 OAI21X1_124 ( .A(_187_), .B(_184_), .C(_189_), .Y(_6__2_) );
INVX1 INVX1_62 ( .A(_6__2_), .Y(_194_) );
OR2X2 OR2X2_94 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_195_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_196_) );
NAND3X1 NAND3X1_63 ( .A(_194_), .B(_196_), .C(_195_), .Y(_197_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_191_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_192_) );
OAI21X1 OAI21X1_125 ( .A(_191_), .B(_192_), .C(_6__2_), .Y(_193_) );
NAND2X1 NAND2X1_93 ( .A(_193_), .B(_197_), .Y(_0__14_) );
OAI21X1 OAI21X1_126 ( .A(_194_), .B(_191_), .C(_196_), .Y(_6__3_) );
INVX1 INVX1_63 ( .A(_6__3_), .Y(_201_) );
OR2X2 OR2X2_95 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_202_) );
NAND2X1 NAND2X1_94 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_203_) );
NAND3X1 NAND3X1_64 ( .A(_201_), .B(_203_), .C(_202_), .Y(_204_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_198_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_199_) );
OAI21X1 OAI21X1_127 ( .A(_198_), .B(_199_), .C(_6__3_), .Y(_200_) );
NAND2X1 NAND2X1_95 ( .A(_200_), .B(_204_), .Y(_0__15_) );
OAI21X1 OAI21X1_128 ( .A(_201_), .B(_198_), .C(_203_), .Y(_5_) );
INVX1 INVX1_64 ( .A(w_cout_3_), .Y(_208_) );
OR2X2 OR2X2_96 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_209_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_210_) );
NAND3X1 NAND3X1_65 ( .A(_208_), .B(_210_), .C(_209_), .Y(_211_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_205_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_206_) );
OAI21X1 OAI21X1_129 ( .A(_205_), .B(_206_), .C(w_cout_3_), .Y(_207_) );
NAND2X1 NAND2X1_97 ( .A(_207_), .B(_211_), .Y(_0__16_) );
OAI21X1 OAI21X1_130 ( .A(_208_), .B(_205_), .C(_210_), .Y(_8__1_) );
INVX1 INVX1_65 ( .A(_8__1_), .Y(_215_) );
OR2X2 OR2X2_97 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_216_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_217_) );
NAND3X1 NAND3X1_66 ( .A(_215_), .B(_217_), .C(_216_), .Y(_218_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_212_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_213_) );
OAI21X1 OAI21X1_131 ( .A(_212_), .B(_213_), .C(_8__1_), .Y(_214_) );
NAND2X1 NAND2X1_99 ( .A(_214_), .B(_218_), .Y(_0__17_) );
OAI21X1 OAI21X1_132 ( .A(_215_), .B(_212_), .C(_217_), .Y(_8__2_) );
INVX1 INVX1_66 ( .A(_8__2_), .Y(_222_) );
OR2X2 OR2X2_98 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_223_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_224_) );
NAND3X1 NAND3X1_67 ( .A(_222_), .B(_224_), .C(_223_), .Y(_225_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_219_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_220_) );
OAI21X1 OAI21X1_133 ( .A(_219_), .B(_220_), .C(_8__2_), .Y(_221_) );
NAND2X1 NAND2X1_101 ( .A(_221_), .B(_225_), .Y(_0__18_) );
OAI21X1 OAI21X1_134 ( .A(_222_), .B(_219_), .C(_224_), .Y(_8__3_) );
INVX1 INVX1_67 ( .A(_8__3_), .Y(_229_) );
OR2X2 OR2X2_99 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_230_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_231_) );
NAND3X1 NAND3X1_68 ( .A(_229_), .B(_231_), .C(_230_), .Y(_232_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_226_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_227_) );
OAI21X1 OAI21X1_135 ( .A(_226_), .B(_227_), .C(_8__3_), .Y(_228_) );
NAND2X1 NAND2X1_103 ( .A(_228_), .B(_232_), .Y(_0__19_) );
OAI21X1 OAI21X1_136 ( .A(_229_), .B(_226_), .C(_231_), .Y(_7_) );
INVX1 INVX1_68 ( .A(w_cout_4_), .Y(_236_) );
OR2X2 OR2X2_100 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_237_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_238_) );
NAND3X1 NAND3X1_69 ( .A(_236_), .B(_238_), .C(_237_), .Y(_239_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_233_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_234_) );
OAI21X1 OAI21X1_137 ( .A(_233_), .B(_234_), .C(w_cout_4_), .Y(_235_) );
NAND2X1 NAND2X1_105 ( .A(_235_), .B(_239_), .Y(_0__20_) );
OAI21X1 OAI21X1_138 ( .A(_236_), .B(_233_), .C(_238_), .Y(_10__1_) );
INVX1 INVX1_69 ( .A(_10__1_), .Y(_243_) );
OR2X2 OR2X2_101 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_244_) );
NAND2X1 NAND2X1_106 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_245_) );
NAND3X1 NAND3X1_70 ( .A(_243_), .B(_245_), .C(_244_), .Y(_246_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_240_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_241_) );
OAI21X1 OAI21X1_139 ( .A(_240_), .B(_241_), .C(_10__1_), .Y(_242_) );
NAND2X1 NAND2X1_107 ( .A(_242_), .B(_246_), .Y(_0__21_) );
OAI21X1 OAI21X1_140 ( .A(_243_), .B(_240_), .C(_245_), .Y(_10__2_) );
INVX1 INVX1_70 ( .A(_10__2_), .Y(_250_) );
OR2X2 OR2X2_102 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_251_) );
NAND2X1 NAND2X1_108 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_252_) );
NAND3X1 NAND3X1_71 ( .A(_250_), .B(_252_), .C(_251_), .Y(_253_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_247_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_248_) );
OAI21X1 OAI21X1_141 ( .A(_247_), .B(_248_), .C(_10__2_), .Y(_249_) );
NAND2X1 NAND2X1_109 ( .A(_249_), .B(_253_), .Y(_0__22_) );
OAI21X1 OAI21X1_142 ( .A(_250_), .B(_247_), .C(_252_), .Y(_10__3_) );
INVX1 INVX1_71 ( .A(_10__3_), .Y(_257_) );
OR2X2 OR2X2_103 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_258_) );
NAND2X1 NAND2X1_110 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_259_) );
NAND3X1 NAND3X1_72 ( .A(_257_), .B(_259_), .C(_258_), .Y(_260_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_254_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_255_) );
OAI21X1 OAI21X1_143 ( .A(_254_), .B(_255_), .C(_10__3_), .Y(_256_) );
NAND2X1 NAND2X1_111 ( .A(_256_), .B(_260_), .Y(_0__23_) );
OAI21X1 OAI21X1_144 ( .A(_257_), .B(_254_), .C(_259_), .Y(_9_) );
INVX1 INVX1_72 ( .A(w_cout_5_), .Y(_264_) );
OR2X2 OR2X2_104 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_265_) );
NAND2X1 NAND2X1_112 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_266_) );
NAND3X1 NAND3X1_73 ( .A(_264_), .B(_266_), .C(_265_), .Y(_267_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_261_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_262_) );
OAI21X1 OAI21X1_145 ( .A(_261_), .B(_262_), .C(w_cout_5_), .Y(_263_) );
NAND2X1 NAND2X1_113 ( .A(_263_), .B(_267_), .Y(_0__24_) );
OAI21X1 OAI21X1_146 ( .A(_264_), .B(_261_), .C(_266_), .Y(_12__1_) );
INVX1 INVX1_73 ( .A(_12__1_), .Y(_271_) );
OR2X2 OR2X2_105 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_272_) );
NAND2X1 NAND2X1_114 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_273_) );
NAND3X1 NAND3X1_74 ( .A(_271_), .B(_273_), .C(_272_), .Y(_274_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_268_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_269_) );
OAI21X1 OAI21X1_147 ( .A(_268_), .B(_269_), .C(_12__1_), .Y(_270_) );
NAND2X1 NAND2X1_115 ( .A(_270_), .B(_274_), .Y(_0__25_) );
OAI21X1 OAI21X1_148 ( .A(_271_), .B(_268_), .C(_273_), .Y(_12__2_) );
INVX1 INVX1_74 ( .A(_12__2_), .Y(_278_) );
OR2X2 OR2X2_106 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_279_) );
NAND2X1 NAND2X1_116 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_280_) );
NAND3X1 NAND3X1_75 ( .A(_278_), .B(_280_), .C(_279_), .Y(_281_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_275_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_276_) );
OAI21X1 OAI21X1_149 ( .A(_275_), .B(_276_), .C(_12__2_), .Y(_277_) );
NAND2X1 NAND2X1_117 ( .A(_277_), .B(_281_), .Y(_0__26_) );
OAI21X1 OAI21X1_150 ( .A(_278_), .B(_275_), .C(_280_), .Y(_12__3_) );
INVX1 INVX1_75 ( .A(_12__3_), .Y(_285_) );
OR2X2 OR2X2_107 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_286_) );
NAND2X1 NAND2X1_118 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_287_) );
NAND3X1 NAND3X1_76 ( .A(_285_), .B(_287_), .C(_286_), .Y(_288_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_282_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_283_) );
OAI21X1 OAI21X1_151 ( .A(_282_), .B(_283_), .C(_12__3_), .Y(_284_) );
NAND2X1 NAND2X1_119 ( .A(_284_), .B(_288_), .Y(_0__27_) );
OAI21X1 OAI21X1_152 ( .A(_285_), .B(_282_), .C(_287_), .Y(_11_) );
INVX1 INVX1_76 ( .A(w_cout_6_), .Y(_292_) );
OR2X2 OR2X2_108 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_293_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_294_) );
NAND3X1 NAND3X1_77 ( .A(_292_), .B(_294_), .C(_293_), .Y(_295_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_289_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_290_) );
OAI21X1 OAI21X1_153 ( .A(_289_), .B(_290_), .C(w_cout_6_), .Y(_291_) );
NAND2X1 NAND2X1_121 ( .A(_291_), .B(_295_), .Y(_0__28_) );
OAI21X1 OAI21X1_154 ( .A(_292_), .B(_289_), .C(_294_), .Y(_14__1_) );
INVX1 INVX1_77 ( .A(_14__1_), .Y(_299_) );
OR2X2 OR2X2_109 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_300_) );
NAND2X1 NAND2X1_122 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_301_) );
NAND3X1 NAND3X1_78 ( .A(_299_), .B(_301_), .C(_300_), .Y(_302_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_296_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_297_) );
OAI21X1 OAI21X1_155 ( .A(_296_), .B(_297_), .C(_14__1_), .Y(_298_) );
NAND2X1 NAND2X1_123 ( .A(_298_), .B(_302_), .Y(_0__29_) );
OAI21X1 OAI21X1_156 ( .A(_299_), .B(_296_), .C(_301_), .Y(_14__2_) );
INVX1 INVX1_78 ( .A(_14__2_), .Y(_306_) );
OR2X2 OR2X2_110 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_307_) );
NAND2X1 NAND2X1_124 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_308_) );
NAND3X1 NAND3X1_79 ( .A(_306_), .B(_308_), .C(_307_), .Y(_309_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_303_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_304_) );
OAI21X1 OAI21X1_157 ( .A(_303_), .B(_304_), .C(_14__2_), .Y(_305_) );
NAND2X1 NAND2X1_125 ( .A(_305_), .B(_309_), .Y(_0__30_) );
OAI21X1 OAI21X1_158 ( .A(_306_), .B(_303_), .C(_308_), .Y(_14__3_) );
INVX1 INVX1_79 ( .A(_14__3_), .Y(_313_) );
OR2X2 OR2X2_111 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_314_) );
NAND2X1 NAND2X1_126 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_315_) );
NAND3X1 NAND3X1_80 ( .A(_313_), .B(_315_), .C(_314_), .Y(_316_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_310_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_311_) );
OAI21X1 OAI21X1_159 ( .A(_310_), .B(_311_), .C(_14__3_), .Y(_312_) );
NAND2X1 NAND2X1_127 ( .A(_312_), .B(_316_), .Y(_0__31_) );
OAI21X1 OAI21X1_160 ( .A(_313_), .B(_310_), .C(_315_), .Y(_13_) );
INVX1 INVX1_80 ( .A(w_cout_7_), .Y(_320_) );
OR2X2 OR2X2_112 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_321_) );
NAND2X1 NAND2X1_128 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_322_) );
BUFX2 BUFX2_66 ( .A(skip0_cin_next), .Y(_2__0_) );
BUFX2 BUFX2_67 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_68 ( .A(w_cout_1_), .Y(_4__0_) );
BUFX2 BUFX2_69 ( .A(_3_), .Y(_4__4_) );
BUFX2 BUFX2_70 ( .A(w_cout_2_), .Y(_6__0_) );
BUFX2 BUFX2_71 ( .A(_5_), .Y(_6__4_) );
BUFX2 BUFX2_72 ( .A(w_cout_3_), .Y(_8__0_) );
BUFX2 BUFX2_73 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_74 ( .A(w_cout_4_), .Y(_10__0_) );
BUFX2 BUFX2_75 ( .A(_9_), .Y(_10__4_) );
BUFX2 BUFX2_76 ( .A(w_cout_5_), .Y(_12__0_) );
BUFX2 BUFX2_77 ( .A(_11_), .Y(_12__4_) );
BUFX2 BUFX2_78 ( .A(w_cout_6_), .Y(_14__0_) );
BUFX2 BUFX2_79 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_80 ( .A(w_cout_7_), .Y(_16__0_) );
BUFX2 BUFX2_81 ( .A(_15_), .Y(_16__4_) );
BUFX2 BUFX2_82 ( .A(w_cout_8_), .Y(_18__0_) );
BUFX2 BUFX2_83 ( .A(_17_), .Y(_18__4_) );
BUFX2 BUFX2_84 ( .A(w_cout_9_), .Y(_20__0_) );
BUFX2 BUFX2_85 ( .A(_19_), .Y(_20__4_) );
BUFX2 BUFX2_86 ( .A(w_cout_10_), .Y(_22__0_) );
BUFX2 BUFX2_87 ( .A(_21_), .Y(_22__4_) );
BUFX2 BUFX2_88 ( .A(w_cout_11_), .Y(_24__0_) );
BUFX2 BUFX2_89 ( .A(_23_), .Y(_24__4_) );
BUFX2 BUFX2_90 ( .A(w_cout_12_), .Y(_26__0_) );
BUFX2 BUFX2_91 ( .A(_25_), .Y(_26__4_) );
BUFX2 BUFX2_92 ( .A(w_cout_13_), .Y(_28__0_) );
BUFX2 BUFX2_93 ( .A(_27_), .Y(_28__4_) );
BUFX2 BUFX2_94 ( .A(w_cout_14_), .Y(_30__0_) );
BUFX2 BUFX2_95 ( .A(_29_), .Y(_30__4_) );
BUFX2 BUFX2_96 ( .A(1'b0), .Y(rca_inst_w_CARRY_0_) );
BUFX2 BUFX2_97 ( .A(cout0), .Y(rca_inst_w_CARRY_4_) );
BUFX2 BUFX2_98 ( .A(skip0_cin_next), .Y(w_cout_0_) );
endmodule
