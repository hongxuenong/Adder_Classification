module CSkipA_26bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term1[6], i_add_term1[7], i_add_term1[8], i_add_term1[9], i_add_term1[10], i_add_term1[11], i_add_term1[12], i_add_term1[13], i_add_term1[14], i_add_term1[15], i_add_term1[16], i_add_term1[17], i_add_term1[18], i_add_term1[19], i_add_term1[20], i_add_term1[21], i_add_term1[22], i_add_term1[23], i_add_term1[24], i_add_term1[25], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], i_add_term2[6], i_add_term2[7], i_add_term2[8], i_add_term2[9], i_add_term2[10], i_add_term2[11], i_add_term2[12], i_add_term2[13], i_add_term2[14], i_add_term2[15], i_add_term2[16], i_add_term2[17], i_add_term2[18], i_add_term2[19], i_add_term2[20], i_add_term2[21], i_add_term2[22], i_add_term2[23], i_add_term2[24], i_add_term2[25], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], sum[6], sum[7], sum[8], sum[9], sum[10], sum[11], sum[12], sum[13], sum[14], sum[15], sum[16], sum[17], sum[18], sum[19], sum[20], sum[21], sum[22], sum[23], sum[24], sum[25], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term1[6];
input i_add_term1[7];
input i_add_term1[8];
input i_add_term1[9];
input i_add_term1[10];
input i_add_term1[11];
input i_add_term1[12];
input i_add_term1[13];
input i_add_term1[14];
input i_add_term1[15];
input i_add_term1[16];
input i_add_term1[17];
input i_add_term1[18];
input i_add_term1[19];
input i_add_term1[20];
input i_add_term1[21];
input i_add_term1[22];
input i_add_term1[23];
input i_add_term1[24];
input i_add_term1[25];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
input i_add_term2[6];
input i_add_term2[7];
input i_add_term2[8];
input i_add_term2[9];
input i_add_term2[10];
input i_add_term2[11];
input i_add_term2[12];
input i_add_term2[13];
input i_add_term2[14];
input i_add_term2[15];
input i_add_term2[16];
input i_add_term2[17];
input i_add_term2[18];
input i_add_term2[19];
input i_add_term2[20];
input i_add_term2[21];
input i_add_term2[22];
input i_add_term2[23];
input i_add_term2[24];
input i_add_term2[25];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output sum[6];
output sum[7];
output sum[8];
output sum[9];
output sum[10];
output sum[11];
output sum[12];
output sum[13];
output sum[14];
output sum[15];
output sum[16];
output sum[17];
output sum[18];
output sum[19];
output sum[20];
output sum[21];
output sum[22];
output sum[23];
output sum[24];
output sum[25];
output cout;

BUFX2 BUFX2_1 ( .A(w_cout_7_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
INVX1 INVX1_1 ( .A(i_add_term1[0]), .Y(_19_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[0]), .B(_19_), .Y(_20_) );
INVX1 INVX1_2 ( .A(i_add_term2[0]), .Y(_21_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term1[0]), .B(_21_), .Y(_22_) );
INVX1 INVX1_3 ( .A(i_add_term1[1]), .Y(_23_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[1]), .B(_23_), .Y(_24_) );
INVX1 INVX1_4 ( .A(i_add_term2[1]), .Y(_25_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term1[1]), .B(_25_), .Y(_26_) );
OAI22X1 OAI22X1_1 ( .A(_20_), .B(_22_), .C(_24_), .D(_26_), .Y(_27_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_28_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_29_) );
NOR2X1 NOR2X1_6 ( .A(_28_), .B(_29_), .Y(_30_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_31_) );
NAND2X1 NAND2X1_1 ( .A(_30_), .B(_31_), .Y(_32_) );
NOR2X1 NOR2X1_7 ( .A(_27_), .B(_32_), .Y(_3_) );
INVX1 INVX1_5 ( .A(_1_), .Y(_33_) );
NAND2X1 NAND2X1_2 ( .A(1'b0), .B(_3_), .Y(_34_) );
OAI21X1 OAI21X1_1 ( .A(_3_), .B(_33_), .C(_34_), .Y(w_cout_1_) );
INVX1 INVX1_6 ( .A(i_add_term1[4]), .Y(_35_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[4]), .B(_35_), .Y(_36_) );
INVX1 INVX1_7 ( .A(i_add_term2[4]), .Y(_37_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term1[4]), .B(_37_), .Y(_38_) );
INVX1 INVX1_8 ( .A(i_add_term1[5]), .Y(_39_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[5]), .B(_39_), .Y(_40_) );
INVX1 INVX1_9 ( .A(i_add_term2[5]), .Y(_41_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term1[5]), .B(_41_), .Y(_42_) );
OAI22X1 OAI22X1_2 ( .A(_36_), .B(_38_), .C(_40_), .D(_42_), .Y(_43_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_44_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_45_) );
NOR2X1 NOR2X1_13 ( .A(_44_), .B(_45_), .Y(_46_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_47_) );
NAND2X1 NAND2X1_3 ( .A(_46_), .B(_47_), .Y(_48_) );
NOR2X1 NOR2X1_14 ( .A(_43_), .B(_48_), .Y(_6_) );
INVX1 INVX1_10 ( .A(_4_), .Y(_49_) );
NAND2X1 NAND2X1_4 ( .A(1'b0), .B(_6_), .Y(_50_) );
OAI21X1 OAI21X1_2 ( .A(_6_), .B(_49_), .C(_50_), .Y(w_cout_2_) );
INVX1 INVX1_11 ( .A(i_add_term1[8]), .Y(_51_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[8]), .B(_51_), .Y(_52_) );
INVX1 INVX1_12 ( .A(i_add_term2[8]), .Y(_53_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term1[8]), .B(_53_), .Y(_54_) );
INVX1 INVX1_13 ( .A(i_add_term1[9]), .Y(_55_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[9]), .B(_55_), .Y(_56_) );
INVX1 INVX1_14 ( .A(i_add_term2[9]), .Y(_57_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term1[9]), .B(_57_), .Y(_58_) );
OAI22X1 OAI22X1_3 ( .A(_52_), .B(_54_), .C(_56_), .D(_58_), .Y(_59_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_60_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_61_) );
NOR2X1 NOR2X1_20 ( .A(_60_), .B(_61_), .Y(_62_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_63_) );
NAND2X1 NAND2X1_5 ( .A(_62_), .B(_63_), .Y(_64_) );
NOR2X1 NOR2X1_21 ( .A(_59_), .B(_64_), .Y(_9_) );
INVX1 INVX1_15 ( .A(_7_), .Y(_65_) );
NAND2X1 NAND2X1_6 ( .A(1'b0), .B(_9_), .Y(_66_) );
OAI21X1 OAI21X1_3 ( .A(_9_), .B(_65_), .C(_66_), .Y(w_cout_3_) );
INVX1 INVX1_16 ( .A(i_add_term1[12]), .Y(_67_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[12]), .B(_67_), .Y(_68_) );
INVX1 INVX1_17 ( .A(i_add_term2[12]), .Y(_69_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term1[12]), .B(_69_), .Y(_70_) );
INVX1 INVX1_18 ( .A(i_add_term1[13]), .Y(_71_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[13]), .B(_71_), .Y(_72_) );
INVX1 INVX1_19 ( .A(i_add_term2[13]), .Y(_73_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term1[13]), .B(_73_), .Y(_74_) );
OAI22X1 OAI22X1_4 ( .A(_68_), .B(_70_), .C(_72_), .D(_74_), .Y(_75_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_76_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_77_) );
NOR2X1 NOR2X1_27 ( .A(_76_), .B(_77_), .Y(_78_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_79_) );
NAND2X1 NAND2X1_7 ( .A(_78_), .B(_79_), .Y(_80_) );
NOR2X1 NOR2X1_28 ( .A(_75_), .B(_80_), .Y(_12_) );
INVX1 INVX1_20 ( .A(_10_), .Y(_81_) );
NAND2X1 NAND2X1_8 ( .A(1'b0), .B(_12_), .Y(_82_) );
OAI21X1 OAI21X1_4 ( .A(_12_), .B(_81_), .C(_82_), .Y(w_cout_4_) );
INVX1 INVX1_21 ( .A(i_add_term1[16]), .Y(_83_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[16]), .B(_83_), .Y(_84_) );
INVX1 INVX1_22 ( .A(i_add_term2[16]), .Y(_85_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term1[16]), .B(_85_), .Y(_86_) );
INVX1 INVX1_23 ( .A(i_add_term1[17]), .Y(_87_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[17]), .B(_87_), .Y(_88_) );
INVX1 INVX1_24 ( .A(i_add_term2[17]), .Y(_89_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term1[17]), .B(_89_), .Y(_90_) );
OAI22X1 OAI22X1_5 ( .A(_84_), .B(_86_), .C(_88_), .D(_90_), .Y(_91_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_92_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_93_) );
NOR2X1 NOR2X1_34 ( .A(_92_), .B(_93_), .Y(_94_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_95_) );
NAND2X1 NAND2X1_9 ( .A(_94_), .B(_95_), .Y(_96_) );
NOR2X1 NOR2X1_35 ( .A(_91_), .B(_96_), .Y(_15_) );
INVX1 INVX1_25 ( .A(_13_), .Y(_97_) );
NAND2X1 NAND2X1_10 ( .A(1'b0), .B(_15_), .Y(_98_) );
OAI21X1 OAI21X1_5 ( .A(_15_), .B(_97_), .C(_98_), .Y(w_cout_5_) );
INVX1 INVX1_26 ( .A(i_add_term1[20]), .Y(_99_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[20]), .B(_99_), .Y(_100_) );
INVX1 INVX1_27 ( .A(i_add_term2[20]), .Y(_101_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term1[20]), .B(_101_), .Y(_102_) );
INVX1 INVX1_28 ( .A(i_add_term1[21]), .Y(_103_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[21]), .B(_103_), .Y(_104_) );
INVX1 INVX1_29 ( .A(i_add_term2[21]), .Y(_105_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term1[21]), .B(_105_), .Y(_106_) );
OAI22X1 OAI22X1_6 ( .A(_100_), .B(_102_), .C(_104_), .D(_106_), .Y(_107_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_108_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_109_) );
NOR2X1 NOR2X1_41 ( .A(_108_), .B(_109_), .Y(_110_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_111_) );
NAND2X1 NAND2X1_11 ( .A(_110_), .B(_111_), .Y(_112_) );
NOR2X1 NOR2X1_42 ( .A(_107_), .B(_112_), .Y(_18_) );
INVX1 INVX1_30 ( .A(_16_), .Y(_113_) );
NAND2X1 NAND2X1_12 ( .A(1'b0), .B(_18_), .Y(_114_) );
OAI21X1 OAI21X1_6 ( .A(_18_), .B(_113_), .C(_114_), .Y(cskip2_inst_cin) );
INVX1 INVX1_31 ( .A(1'b0), .Y(_118_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_119_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_120_) );
NAND3X1 NAND3X1_1 ( .A(_118_), .B(_120_), .C(_119_), .Y(_121_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_115_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_116_) );
OAI21X1 OAI21X1_7 ( .A(_115_), .B(_116_), .C(1'b0), .Y(_117_) );
NAND2X1 NAND2X1_14 ( .A(_117_), .B(_121_), .Y(_0__0_) );
OAI21X1 OAI21X1_8 ( .A(_118_), .B(_115_), .C(_120_), .Y(_2__1_) );
INVX1 INVX1_32 ( .A(_2__1_), .Y(_125_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_126_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_127_) );
NAND3X1 NAND3X1_2 ( .A(_125_), .B(_127_), .C(_126_), .Y(_128_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_122_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_123_) );
OAI21X1 OAI21X1_9 ( .A(_122_), .B(_123_), .C(_2__1_), .Y(_124_) );
NAND2X1 NAND2X1_16 ( .A(_124_), .B(_128_), .Y(_0__1_) );
OAI21X1 OAI21X1_10 ( .A(_125_), .B(_122_), .C(_127_), .Y(_2__2_) );
INVX1 INVX1_33 ( .A(_2__2_), .Y(_132_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_133_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_134_) );
NAND3X1 NAND3X1_3 ( .A(_132_), .B(_134_), .C(_133_), .Y(_135_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_129_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_130_) );
OAI21X1 OAI21X1_11 ( .A(_129_), .B(_130_), .C(_2__2_), .Y(_131_) );
NAND2X1 NAND2X1_18 ( .A(_131_), .B(_135_), .Y(_0__2_) );
OAI21X1 OAI21X1_12 ( .A(_132_), .B(_129_), .C(_134_), .Y(_2__3_) );
INVX1 INVX1_34 ( .A(_2__3_), .Y(_139_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_140_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_141_) );
NAND3X1 NAND3X1_4 ( .A(_139_), .B(_141_), .C(_140_), .Y(_142_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_136_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_137_) );
OAI21X1 OAI21X1_13 ( .A(_136_), .B(_137_), .C(_2__3_), .Y(_138_) );
NAND2X1 NAND2X1_20 ( .A(_138_), .B(_142_), .Y(_0__3_) );
OAI21X1 OAI21X1_14 ( .A(_139_), .B(_136_), .C(_141_), .Y(_1_) );
INVX1 INVX1_35 ( .A(w_cout_1_), .Y(_146_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_147_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_148_) );
NAND3X1 NAND3X1_5 ( .A(_146_), .B(_148_), .C(_147_), .Y(_149_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_143_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_144_) );
OAI21X1 OAI21X1_15 ( .A(_143_), .B(_144_), .C(w_cout_1_), .Y(_145_) );
NAND2X1 NAND2X1_22 ( .A(_145_), .B(_149_), .Y(_0__4_) );
OAI21X1 OAI21X1_16 ( .A(_146_), .B(_143_), .C(_148_), .Y(_5__1_) );
INVX1 INVX1_36 ( .A(_5__1_), .Y(_153_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_154_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_155_) );
NAND3X1 NAND3X1_6 ( .A(_153_), .B(_155_), .C(_154_), .Y(_156_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_150_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_151_) );
OAI21X1 OAI21X1_17 ( .A(_150_), .B(_151_), .C(_5__1_), .Y(_152_) );
NAND2X1 NAND2X1_24 ( .A(_152_), .B(_156_), .Y(_0__5_) );
OAI21X1 OAI21X1_18 ( .A(_153_), .B(_150_), .C(_155_), .Y(_5__2_) );
INVX1 INVX1_37 ( .A(_5__2_), .Y(_160_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_161_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_162_) );
NAND3X1 NAND3X1_7 ( .A(_160_), .B(_162_), .C(_161_), .Y(_163_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_157_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_158_) );
OAI21X1 OAI21X1_19 ( .A(_157_), .B(_158_), .C(_5__2_), .Y(_159_) );
NAND2X1 NAND2X1_26 ( .A(_159_), .B(_163_), .Y(_0__6_) );
OAI21X1 OAI21X1_20 ( .A(_160_), .B(_157_), .C(_162_), .Y(_5__3_) );
INVX1 INVX1_38 ( .A(_5__3_), .Y(_167_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_168_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_169_) );
NAND3X1 NAND3X1_8 ( .A(_167_), .B(_169_), .C(_168_), .Y(_170_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_164_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_165_) );
OAI21X1 OAI21X1_21 ( .A(_164_), .B(_165_), .C(_5__3_), .Y(_166_) );
NAND2X1 NAND2X1_28 ( .A(_166_), .B(_170_), .Y(_0__7_) );
OAI21X1 OAI21X1_22 ( .A(_167_), .B(_164_), .C(_169_), .Y(_4_) );
INVX1 INVX1_39 ( .A(w_cout_2_), .Y(_174_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_175_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_176_) );
NAND3X1 NAND3X1_9 ( .A(_174_), .B(_176_), .C(_175_), .Y(_177_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_171_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_172_) );
OAI21X1 OAI21X1_23 ( .A(_171_), .B(_172_), .C(w_cout_2_), .Y(_173_) );
NAND2X1 NAND2X1_30 ( .A(_173_), .B(_177_), .Y(_0__8_) );
OAI21X1 OAI21X1_24 ( .A(_174_), .B(_171_), .C(_176_), .Y(_8__1_) );
INVX1 INVX1_40 ( .A(_8__1_), .Y(_181_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_182_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_183_) );
NAND3X1 NAND3X1_10 ( .A(_181_), .B(_183_), .C(_182_), .Y(_184_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_178_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_179_) );
OAI21X1 OAI21X1_25 ( .A(_178_), .B(_179_), .C(_8__1_), .Y(_180_) );
NAND2X1 NAND2X1_32 ( .A(_180_), .B(_184_), .Y(_0__9_) );
OAI21X1 OAI21X1_26 ( .A(_181_), .B(_178_), .C(_183_), .Y(_8__2_) );
INVX1 INVX1_41 ( .A(_8__2_), .Y(_188_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_189_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_190_) );
NAND3X1 NAND3X1_11 ( .A(_188_), .B(_190_), .C(_189_), .Y(_191_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_185_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_186_) );
OAI21X1 OAI21X1_27 ( .A(_185_), .B(_186_), .C(_8__2_), .Y(_187_) );
NAND2X1 NAND2X1_34 ( .A(_187_), .B(_191_), .Y(_0__10_) );
OAI21X1 OAI21X1_28 ( .A(_188_), .B(_185_), .C(_190_), .Y(_8__3_) );
INVX1 INVX1_42 ( .A(_8__3_), .Y(_195_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_196_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_197_) );
NAND3X1 NAND3X1_12 ( .A(_195_), .B(_197_), .C(_196_), .Y(_198_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_192_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_193_) );
OAI21X1 OAI21X1_29 ( .A(_192_), .B(_193_), .C(_8__3_), .Y(_194_) );
NAND2X1 NAND2X1_36 ( .A(_194_), .B(_198_), .Y(_0__11_) );
OAI21X1 OAI21X1_30 ( .A(_195_), .B(_192_), .C(_197_), .Y(_7_) );
INVX1 INVX1_43 ( .A(w_cout_3_), .Y(_202_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_203_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_204_) );
NAND3X1 NAND3X1_13 ( .A(_202_), .B(_204_), .C(_203_), .Y(_205_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_199_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_200_) );
OAI21X1 OAI21X1_31 ( .A(_199_), .B(_200_), .C(w_cout_3_), .Y(_201_) );
NAND2X1 NAND2X1_38 ( .A(_201_), .B(_205_), .Y(_0__12_) );
OAI21X1 OAI21X1_32 ( .A(_202_), .B(_199_), .C(_204_), .Y(_11__1_) );
INVX1 INVX1_44 ( .A(_11__1_), .Y(_209_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_210_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_211_) );
NAND3X1 NAND3X1_14 ( .A(_209_), .B(_211_), .C(_210_), .Y(_212_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_206_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_207_) );
OAI21X1 OAI21X1_33 ( .A(_206_), .B(_207_), .C(_11__1_), .Y(_208_) );
NAND2X1 NAND2X1_40 ( .A(_208_), .B(_212_), .Y(_0__13_) );
OAI21X1 OAI21X1_34 ( .A(_209_), .B(_206_), .C(_211_), .Y(_11__2_) );
INVX1 INVX1_45 ( .A(_11__2_), .Y(_216_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_217_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_218_) );
NAND3X1 NAND3X1_15 ( .A(_216_), .B(_218_), .C(_217_), .Y(_219_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_213_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_214_) );
OAI21X1 OAI21X1_35 ( .A(_213_), .B(_214_), .C(_11__2_), .Y(_215_) );
NAND2X1 NAND2X1_42 ( .A(_215_), .B(_219_), .Y(_0__14_) );
OAI21X1 OAI21X1_36 ( .A(_216_), .B(_213_), .C(_218_), .Y(_11__3_) );
INVX1 INVX1_46 ( .A(_11__3_), .Y(_223_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_224_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_225_) );
NAND3X1 NAND3X1_16 ( .A(_223_), .B(_225_), .C(_224_), .Y(_226_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_220_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_221_) );
OAI21X1 OAI21X1_37 ( .A(_220_), .B(_221_), .C(_11__3_), .Y(_222_) );
NAND2X1 NAND2X1_44 ( .A(_222_), .B(_226_), .Y(_0__15_) );
OAI21X1 OAI21X1_38 ( .A(_223_), .B(_220_), .C(_225_), .Y(_10_) );
INVX1 INVX1_47 ( .A(w_cout_4_), .Y(_230_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_231_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_232_) );
NAND3X1 NAND3X1_17 ( .A(_230_), .B(_232_), .C(_231_), .Y(_233_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_227_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_228_) );
OAI21X1 OAI21X1_39 ( .A(_227_), .B(_228_), .C(w_cout_4_), .Y(_229_) );
NAND2X1 NAND2X1_46 ( .A(_229_), .B(_233_), .Y(_0__16_) );
OAI21X1 OAI21X1_40 ( .A(_230_), .B(_227_), .C(_232_), .Y(_14__1_) );
INVX1 INVX1_48 ( .A(_14__1_), .Y(_237_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_238_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_239_) );
NAND3X1 NAND3X1_18 ( .A(_237_), .B(_239_), .C(_238_), .Y(_240_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_234_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_235_) );
OAI21X1 OAI21X1_41 ( .A(_234_), .B(_235_), .C(_14__1_), .Y(_236_) );
NAND2X1 NAND2X1_48 ( .A(_236_), .B(_240_), .Y(_0__17_) );
OAI21X1 OAI21X1_42 ( .A(_237_), .B(_234_), .C(_239_), .Y(_14__2_) );
INVX1 INVX1_49 ( .A(_14__2_), .Y(_244_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_245_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_246_) );
NAND3X1 NAND3X1_19 ( .A(_244_), .B(_246_), .C(_245_), .Y(_247_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_241_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_242_) );
OAI21X1 OAI21X1_43 ( .A(_241_), .B(_242_), .C(_14__2_), .Y(_243_) );
NAND2X1 NAND2X1_50 ( .A(_243_), .B(_247_), .Y(_0__18_) );
OAI21X1 OAI21X1_44 ( .A(_244_), .B(_241_), .C(_246_), .Y(_14__3_) );
INVX1 INVX1_50 ( .A(_14__3_), .Y(_251_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_252_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_253_) );
NAND3X1 NAND3X1_20 ( .A(_251_), .B(_253_), .C(_252_), .Y(_254_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_248_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_249_) );
OAI21X1 OAI21X1_45 ( .A(_248_), .B(_249_), .C(_14__3_), .Y(_250_) );
NAND2X1 NAND2X1_52 ( .A(_250_), .B(_254_), .Y(_0__19_) );
OAI21X1 OAI21X1_46 ( .A(_251_), .B(_248_), .C(_253_), .Y(_13_) );
INVX1 INVX1_51 ( .A(w_cout_5_), .Y(_258_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_259_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_260_) );
NAND3X1 NAND3X1_21 ( .A(_258_), .B(_260_), .C(_259_), .Y(_261_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_255_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_256_) );
OAI21X1 OAI21X1_47 ( .A(_255_), .B(_256_), .C(w_cout_5_), .Y(_257_) );
NAND2X1 NAND2X1_54 ( .A(_257_), .B(_261_), .Y(_0__20_) );
OAI21X1 OAI21X1_48 ( .A(_258_), .B(_255_), .C(_260_), .Y(_17__1_) );
INVX1 INVX1_52 ( .A(_17__1_), .Y(_265_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_266_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_267_) );
NAND3X1 NAND3X1_22 ( .A(_265_), .B(_267_), .C(_266_), .Y(_268_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_262_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_263_) );
OAI21X1 OAI21X1_49 ( .A(_262_), .B(_263_), .C(_17__1_), .Y(_264_) );
NAND2X1 NAND2X1_56 ( .A(_264_), .B(_268_), .Y(_0__21_) );
OAI21X1 OAI21X1_50 ( .A(_265_), .B(_262_), .C(_267_), .Y(_17__2_) );
INVX1 INVX1_53 ( .A(_17__2_), .Y(_272_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_273_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_274_) );
NAND3X1 NAND3X1_23 ( .A(_272_), .B(_274_), .C(_273_), .Y(_275_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_269_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_270_) );
OAI21X1 OAI21X1_51 ( .A(_269_), .B(_270_), .C(_17__2_), .Y(_271_) );
NAND2X1 NAND2X1_58 ( .A(_271_), .B(_275_), .Y(_0__22_) );
OAI21X1 OAI21X1_52 ( .A(_272_), .B(_269_), .C(_274_), .Y(_17__3_) );
INVX1 INVX1_54 ( .A(_17__3_), .Y(_279_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_280_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_281_) );
NAND3X1 NAND3X1_24 ( .A(_279_), .B(_281_), .C(_280_), .Y(_282_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_276_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_277_) );
OAI21X1 OAI21X1_53 ( .A(_276_), .B(_277_), .C(_17__3_), .Y(_278_) );
NAND2X1 NAND2X1_60 ( .A(_278_), .B(_282_), .Y(_0__23_) );
OAI21X1 OAI21X1_54 ( .A(_279_), .B(_276_), .C(_281_), .Y(_16_) );
INVX1 INVX1_55 ( .A(cskip2_inst_cin), .Y(_286_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_287_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_288_) );
NAND3X1 NAND3X1_25 ( .A(_286_), .B(_288_), .C(_287_), .Y(_289_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_283_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_284_) );
OAI21X1 OAI21X1_55 ( .A(_283_), .B(_284_), .C(cskip2_inst_cin), .Y(_285_) );
NAND2X1 NAND2X1_62 ( .A(_285_), .B(_289_), .Y(_0__24_) );
OAI21X1 OAI21X1_56 ( .A(_286_), .B(_283_), .C(_288_), .Y(cskip2_inst_rca0_w_CARRY_1_) );
INVX1 INVX1_56 ( .A(cskip2_inst_rca0_w_CARRY_1_), .Y(_293_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_294_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_295_) );
NAND3X1 NAND3X1_26 ( .A(_293_), .B(_295_), .C(_294_), .Y(_296_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_290_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_291_) );
OAI21X1 OAI21X1_57 ( .A(_290_), .B(_291_), .C(cskip2_inst_rca0_w_CARRY_1_), .Y(_292_) );
NAND2X1 NAND2X1_64 ( .A(_292_), .B(_296_), .Y(_0__25_) );
OAI21X1 OAI21X1_58 ( .A(_293_), .B(_290_), .C(_295_), .Y(cskip2_inst_rca0_w_CARRY_2_) );
INVX1 INVX1_57 ( .A(cskip2_inst_rca0_w_CARRY_2_), .Y(_298_) );
NAND2X1 NAND2X1_65 ( .A(1'b0), .B(1'b0), .Y(_299_) );
NOR2X1 NOR2X1_69 ( .A(1'b0), .B(1'b0), .Y(_297_) );
OAI21X1 OAI21X1_59 ( .A(_298_), .B(_297_), .C(_299_), .Y(cskip2_inst_rca0_w_CARRY_3_) );
INVX1 INVX1_58 ( .A(cskip2_inst_rca0_w_CARRY_3_), .Y(_301_) );
NAND2X1 NAND2X1_66 ( .A(1'b0), .B(1'b0), .Y(_302_) );
NOR2X1 NOR2X1_70 ( .A(1'b0), .B(1'b0), .Y(_300_) );
OAI21X1 OAI21X1_60 ( .A(_301_), .B(_300_), .C(_302_), .Y(cskip2_inst_cout0) );
INVX1 INVX1_59 ( .A(i_add_term1[25]), .Y(_307_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[25]), .B(_307_), .Y(_308_) );
INVX1 INVX1_60 ( .A(i_add_term2[25]), .Y(_309_) );
NAND2X1 NAND2X1_68 ( .A(i_add_term1[25]), .B(_309_), .Y(_310_) );
INVX1 INVX1_61 ( .A(i_add_term1[24]), .Y(_303_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[24]), .B(_303_), .Y(_304_) );
INVX1 INVX1_62 ( .A(i_add_term2[24]), .Y(_305_) );
NAND2X1 NAND2X1_70 ( .A(i_add_term1[24]), .B(_305_), .Y(_306_) );
AOI22X1 AOI22X1_1 ( .A(_308_), .B(_310_), .C(_304_), .D(_306_), .Y(cskip2_inst_skip0_P) );
INVX1 INVX1_63 ( .A(cskip2_inst_cout0), .Y(_311_) );
NAND2X1 NAND2X1_71 ( .A(1'b0), .B(cskip2_inst_skip0_P), .Y(_312_) );
OAI21X1 OAI21X1_61 ( .A(cskip2_inst_skip0_P), .B(_311_), .C(_312_), .Y(w_cout_7_) );
BUFX2 BUFX2_28 ( .A(1'b0), .Y(_2__0_) );
BUFX2 BUFX2_29 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_30 ( .A(w_cout_1_), .Y(_5__0_) );
BUFX2 BUFX2_31 ( .A(_4_), .Y(_5__4_) );
BUFX2 BUFX2_32 ( .A(w_cout_2_), .Y(_8__0_) );
BUFX2 BUFX2_33 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_34 ( .A(w_cout_3_), .Y(_11__0_) );
BUFX2 BUFX2_35 ( .A(_10_), .Y(_11__4_) );
BUFX2 BUFX2_36 ( .A(w_cout_4_), .Y(_14__0_) );
BUFX2 BUFX2_37 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_38 ( .A(w_cout_5_), .Y(_17__0_) );
BUFX2 BUFX2_39 ( .A(_16_), .Y(_17__4_) );
BUFX2 BUFX2_40 ( .A(cskip2_inst_cin), .Y(cskip2_inst_rca0_w_CARRY_0_) );
BUFX2 BUFX2_41 ( .A(cskip2_inst_cout0), .Y(cskip2_inst_rca0_w_CARRY_4_) );
BUFX2 BUFX2_42 ( .A(1'b0), .Y(w_cout_0_) );
BUFX2 BUFX2_43 ( .A(cskip2_inst_cin), .Y(w_cout_6_) );
endmodule
