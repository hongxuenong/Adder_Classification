module CSkipA_58bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [57:0] i_add_term1;
input [57:0] i_add_term2;
output [57:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

INVX1 INVX1_1 ( .A(gnd), .Y(_270_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_271_) );
NAND2X1 NAND2X1_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_272_) );
NAND3X1 NAND3X1_1 ( .A(_270_), .B(_272_), .C(_271_), .Y(_273_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_267_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_268_) );
OAI21X1 OAI21X1_1 ( .A(_267_), .B(_268_), .C(gnd), .Y(_269_) );
NAND2X1 NAND2X1_2 ( .A(_269_), .B(_273_), .Y(_0__0_) );
OAI21X1 OAI21X1_2 ( .A(_270_), .B(_267_), .C(_272_), .Y(_2__1_) );
INVX1 INVX1_2 ( .A(_2__1_), .Y(_277_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_278_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_279_) );
NAND3X1 NAND3X1_2 ( .A(_277_), .B(_279_), .C(_278_), .Y(_280_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_274_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_275_) );
OAI21X1 OAI21X1_3 ( .A(_274_), .B(_275_), .C(_2__1_), .Y(_276_) );
NAND2X1 NAND2X1_4 ( .A(_276_), .B(_280_), .Y(_0__1_) );
OAI21X1 OAI21X1_4 ( .A(_277_), .B(_274_), .C(_279_), .Y(_2__2_) );
INVX1 INVX1_3 ( .A(_2__2_), .Y(_284_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_285_) );
NAND2X1 NAND2X1_5 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_286_) );
NAND3X1 NAND3X1_3 ( .A(_284_), .B(_286_), .C(_285_), .Y(_287_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_281_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_282_) );
OAI21X1 OAI21X1_5 ( .A(_281_), .B(_282_), .C(_2__2_), .Y(_283_) );
NAND2X1 NAND2X1_6 ( .A(_283_), .B(_287_), .Y(_0__2_) );
OAI21X1 OAI21X1_6 ( .A(_284_), .B(_281_), .C(_286_), .Y(_2__3_) );
INVX1 INVX1_4 ( .A(_2__3_), .Y(_291_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_292_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_293_) );
NAND3X1 NAND3X1_4 ( .A(_291_), .B(_293_), .C(_292_), .Y(_294_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_288_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_289_) );
OAI21X1 OAI21X1_7 ( .A(_288_), .B(_289_), .C(_2__3_), .Y(_290_) );
NAND2X1 NAND2X1_8 ( .A(_290_), .B(_294_), .Y(_0__3_) );
OAI21X1 OAI21X1_8 ( .A(_291_), .B(_288_), .C(_293_), .Y(_1_) );
INVX1 INVX1_5 ( .A(w_cout_1_), .Y(_298_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_299_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_300_) );
NAND3X1 NAND3X1_5 ( .A(_298_), .B(_300_), .C(_299_), .Y(_301_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_295_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_296_) );
OAI21X1 OAI21X1_9 ( .A(_295_), .B(_296_), .C(w_cout_1_), .Y(_297_) );
NAND2X1 NAND2X1_10 ( .A(_297_), .B(_301_), .Y(_0__4_) );
OAI21X1 OAI21X1_10 ( .A(_298_), .B(_295_), .C(_300_), .Y(_5__1_) );
INVX1 INVX1_6 ( .A(_5__1_), .Y(_305_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_306_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_307_) );
NAND3X1 NAND3X1_6 ( .A(_305_), .B(_307_), .C(_306_), .Y(_308_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_302_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_303_) );
OAI21X1 OAI21X1_11 ( .A(_302_), .B(_303_), .C(_5__1_), .Y(_304_) );
NAND2X1 NAND2X1_12 ( .A(_304_), .B(_308_), .Y(_0__5_) );
OAI21X1 OAI21X1_12 ( .A(_305_), .B(_302_), .C(_307_), .Y(_5__2_) );
INVX1 INVX1_7 ( .A(_5__2_), .Y(_312_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_313_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_314_) );
NAND3X1 NAND3X1_7 ( .A(_312_), .B(_314_), .C(_313_), .Y(_315_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_309_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_310_) );
OAI21X1 OAI21X1_13 ( .A(_309_), .B(_310_), .C(_5__2_), .Y(_311_) );
NAND2X1 NAND2X1_14 ( .A(_311_), .B(_315_), .Y(_0__6_) );
OAI21X1 OAI21X1_14 ( .A(_312_), .B(_309_), .C(_314_), .Y(_5__3_) );
INVX1 INVX1_8 ( .A(_5__3_), .Y(_319_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_320_) );
NAND2X1 NAND2X1_15 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_321_) );
NAND3X1 NAND3X1_8 ( .A(_319_), .B(_321_), .C(_320_), .Y(_322_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_316_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_317_) );
OAI21X1 OAI21X1_15 ( .A(_316_), .B(_317_), .C(_5__3_), .Y(_318_) );
NAND2X1 NAND2X1_16 ( .A(_318_), .B(_322_), .Y(_0__7_) );
OAI21X1 OAI21X1_16 ( .A(_319_), .B(_316_), .C(_321_), .Y(_4_) );
INVX1 INVX1_9 ( .A(w_cout_2_), .Y(_326_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_327_) );
NAND2X1 NAND2X1_17 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_328_) );
NAND3X1 NAND3X1_9 ( .A(_326_), .B(_328_), .C(_327_), .Y(_329_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_323_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_324_) );
OAI21X1 OAI21X1_17 ( .A(_323_), .B(_324_), .C(w_cout_2_), .Y(_325_) );
NAND2X1 NAND2X1_18 ( .A(_325_), .B(_329_), .Y(_0__8_) );
OAI21X1 OAI21X1_18 ( .A(_326_), .B(_323_), .C(_328_), .Y(_8__1_) );
INVX1 INVX1_10 ( .A(_8__1_), .Y(_333_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_334_) );
NAND2X1 NAND2X1_19 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_335_) );
NAND3X1 NAND3X1_10 ( .A(_333_), .B(_335_), .C(_334_), .Y(_336_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_330_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_331_) );
OAI21X1 OAI21X1_19 ( .A(_330_), .B(_331_), .C(_8__1_), .Y(_332_) );
NAND2X1 NAND2X1_20 ( .A(_332_), .B(_336_), .Y(_0__9_) );
OAI21X1 OAI21X1_20 ( .A(_333_), .B(_330_), .C(_335_), .Y(_8__2_) );
INVX1 INVX1_11 ( .A(_8__2_), .Y(_340_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_341_) );
NAND2X1 NAND2X1_21 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_342_) );
NAND3X1 NAND3X1_11 ( .A(_340_), .B(_342_), .C(_341_), .Y(_343_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_337_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_338_) );
OAI21X1 OAI21X1_21 ( .A(_337_), .B(_338_), .C(_8__2_), .Y(_339_) );
NAND2X1 NAND2X1_22 ( .A(_339_), .B(_343_), .Y(_0__10_) );
OAI21X1 OAI21X1_22 ( .A(_340_), .B(_337_), .C(_342_), .Y(_8__3_) );
INVX1 INVX1_12 ( .A(_8__3_), .Y(_347_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_348_) );
NAND2X1 NAND2X1_23 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_349_) );
NAND3X1 NAND3X1_12 ( .A(_347_), .B(_349_), .C(_348_), .Y(_350_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_344_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_345_) );
OAI21X1 OAI21X1_23 ( .A(_344_), .B(_345_), .C(_8__3_), .Y(_346_) );
NAND2X1 NAND2X1_24 ( .A(_346_), .B(_350_), .Y(_0__11_) );
OAI21X1 OAI21X1_24 ( .A(_347_), .B(_344_), .C(_349_), .Y(_7_) );
INVX1 INVX1_13 ( .A(w_cout_3_), .Y(_354_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_355_) );
NAND2X1 NAND2X1_25 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_356_) );
NAND3X1 NAND3X1_13 ( .A(_354_), .B(_356_), .C(_355_), .Y(_357_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_351_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_352_) );
OAI21X1 OAI21X1_25 ( .A(_351_), .B(_352_), .C(w_cout_3_), .Y(_353_) );
NAND2X1 NAND2X1_26 ( .A(_353_), .B(_357_), .Y(_0__12_) );
OAI21X1 OAI21X1_26 ( .A(_354_), .B(_351_), .C(_356_), .Y(_11__1_) );
INVX1 INVX1_14 ( .A(_11__1_), .Y(_361_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_362_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_363_) );
NAND3X1 NAND3X1_14 ( .A(_361_), .B(_363_), .C(_362_), .Y(_364_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_358_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_359_) );
OAI21X1 OAI21X1_27 ( .A(_358_), .B(_359_), .C(_11__1_), .Y(_360_) );
NAND2X1 NAND2X1_28 ( .A(_360_), .B(_364_), .Y(_0__13_) );
OAI21X1 OAI21X1_28 ( .A(_361_), .B(_358_), .C(_363_), .Y(_11__2_) );
INVX1 INVX1_15 ( .A(_11__2_), .Y(_368_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_369_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_370_) );
NAND3X1 NAND3X1_15 ( .A(_368_), .B(_370_), .C(_369_), .Y(_371_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_365_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_366_) );
OAI21X1 OAI21X1_29 ( .A(_365_), .B(_366_), .C(_11__2_), .Y(_367_) );
NAND2X1 NAND2X1_30 ( .A(_367_), .B(_371_), .Y(_0__14_) );
OAI21X1 OAI21X1_30 ( .A(_368_), .B(_365_), .C(_370_), .Y(_11__3_) );
INVX1 INVX1_16 ( .A(_11__3_), .Y(_375_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_376_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_377_) );
NAND3X1 NAND3X1_16 ( .A(_375_), .B(_377_), .C(_376_), .Y(_378_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_372_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_373_) );
OAI21X1 OAI21X1_31 ( .A(_372_), .B(_373_), .C(_11__3_), .Y(_374_) );
NAND2X1 NAND2X1_32 ( .A(_374_), .B(_378_), .Y(_0__15_) );
OAI21X1 OAI21X1_32 ( .A(_375_), .B(_372_), .C(_377_), .Y(_10_) );
INVX1 INVX1_17 ( .A(w_cout_4_), .Y(_382_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_383_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_384_) );
NAND3X1 NAND3X1_17 ( .A(_382_), .B(_384_), .C(_383_), .Y(_385_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_379_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_380_) );
OAI21X1 OAI21X1_33 ( .A(_379_), .B(_380_), .C(w_cout_4_), .Y(_381_) );
NAND2X1 NAND2X1_34 ( .A(_381_), .B(_385_), .Y(_0__16_) );
OAI21X1 OAI21X1_34 ( .A(_382_), .B(_379_), .C(_384_), .Y(_14__1_) );
INVX1 INVX1_18 ( .A(_14__1_), .Y(_389_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_390_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_391_) );
NAND3X1 NAND3X1_18 ( .A(_389_), .B(_391_), .C(_390_), .Y(_392_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_386_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_387_) );
OAI21X1 OAI21X1_35 ( .A(_386_), .B(_387_), .C(_14__1_), .Y(_388_) );
NAND2X1 NAND2X1_36 ( .A(_388_), .B(_392_), .Y(_0__17_) );
OAI21X1 OAI21X1_36 ( .A(_389_), .B(_386_), .C(_391_), .Y(_14__2_) );
INVX1 INVX1_19 ( .A(_14__2_), .Y(_396_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_397_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_398_) );
NAND3X1 NAND3X1_19 ( .A(_396_), .B(_398_), .C(_397_), .Y(_399_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_393_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_394_) );
OAI21X1 OAI21X1_37 ( .A(_393_), .B(_394_), .C(_14__2_), .Y(_395_) );
NAND2X1 NAND2X1_38 ( .A(_395_), .B(_399_), .Y(_0__18_) );
OAI21X1 OAI21X1_38 ( .A(_396_), .B(_393_), .C(_398_), .Y(_14__3_) );
INVX1 INVX1_20 ( .A(_14__3_), .Y(_403_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_404_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_405_) );
NAND3X1 NAND3X1_20 ( .A(_403_), .B(_405_), .C(_404_), .Y(_406_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_400_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_401_) );
OAI21X1 OAI21X1_39 ( .A(_400_), .B(_401_), .C(_14__3_), .Y(_402_) );
NAND2X1 NAND2X1_40 ( .A(_402_), .B(_406_), .Y(_0__19_) );
OAI21X1 OAI21X1_40 ( .A(_403_), .B(_400_), .C(_405_), .Y(_13_) );
INVX1 INVX1_21 ( .A(w_cout_5_), .Y(_410_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_411_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_412_) );
NAND3X1 NAND3X1_21 ( .A(_410_), .B(_412_), .C(_411_), .Y(_413_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_407_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_408_) );
OAI21X1 OAI21X1_41 ( .A(_407_), .B(_408_), .C(w_cout_5_), .Y(_409_) );
NAND2X1 NAND2X1_42 ( .A(_409_), .B(_413_), .Y(_0__20_) );
OAI21X1 OAI21X1_42 ( .A(_410_), .B(_407_), .C(_412_), .Y(_17__1_) );
INVX1 INVX1_22 ( .A(_17__1_), .Y(_417_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_418_) );
NAND2X1 NAND2X1_43 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_419_) );
NAND3X1 NAND3X1_22 ( .A(_417_), .B(_419_), .C(_418_), .Y(_420_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_414_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_415_) );
OAI21X1 OAI21X1_43 ( .A(_414_), .B(_415_), .C(_17__1_), .Y(_416_) );
NAND2X1 NAND2X1_44 ( .A(_416_), .B(_420_), .Y(_0__21_) );
OAI21X1 OAI21X1_44 ( .A(_417_), .B(_414_), .C(_419_), .Y(_17__2_) );
INVX1 INVX1_23 ( .A(_17__2_), .Y(_424_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_425_) );
NAND2X1 NAND2X1_45 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_426_) );
NAND3X1 NAND3X1_23 ( .A(_424_), .B(_426_), .C(_425_), .Y(_427_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_421_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_422_) );
OAI21X1 OAI21X1_45 ( .A(_421_), .B(_422_), .C(_17__2_), .Y(_423_) );
NAND2X1 NAND2X1_46 ( .A(_423_), .B(_427_), .Y(_0__22_) );
OAI21X1 OAI21X1_46 ( .A(_424_), .B(_421_), .C(_426_), .Y(_17__3_) );
INVX1 INVX1_24 ( .A(_17__3_), .Y(_431_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_432_) );
NAND2X1 NAND2X1_47 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_433_) );
NAND3X1 NAND3X1_24 ( .A(_431_), .B(_433_), .C(_432_), .Y(_434_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_428_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_429_) );
OAI21X1 OAI21X1_47 ( .A(_428_), .B(_429_), .C(_17__3_), .Y(_430_) );
NAND2X1 NAND2X1_48 ( .A(_430_), .B(_434_), .Y(_0__23_) );
OAI21X1 OAI21X1_48 ( .A(_431_), .B(_428_), .C(_433_), .Y(_16_) );
INVX1 INVX1_25 ( .A(w_cout_6_), .Y(_438_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_439_) );
NAND2X1 NAND2X1_49 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_440_) );
NAND3X1 NAND3X1_25 ( .A(_438_), .B(_440_), .C(_439_), .Y(_441_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_435_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_436_) );
OAI21X1 OAI21X1_49 ( .A(_435_), .B(_436_), .C(w_cout_6_), .Y(_437_) );
NAND2X1 NAND2X1_50 ( .A(_437_), .B(_441_), .Y(_0__24_) );
OAI21X1 OAI21X1_50 ( .A(_438_), .B(_435_), .C(_440_), .Y(_20__1_) );
INVX1 INVX1_26 ( .A(_20__1_), .Y(_445_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_446_) );
NAND2X1 NAND2X1_51 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_447_) );
NAND3X1 NAND3X1_26 ( .A(_445_), .B(_447_), .C(_446_), .Y(_448_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_442_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_443_) );
OAI21X1 OAI21X1_51 ( .A(_442_), .B(_443_), .C(_20__1_), .Y(_444_) );
NAND2X1 NAND2X1_52 ( .A(_444_), .B(_448_), .Y(_0__25_) );
OAI21X1 OAI21X1_52 ( .A(_445_), .B(_442_), .C(_447_), .Y(_20__2_) );
INVX1 INVX1_27 ( .A(_20__2_), .Y(_452_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_453_) );
NAND2X1 NAND2X1_53 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_454_) );
NAND3X1 NAND3X1_27 ( .A(_452_), .B(_454_), .C(_453_), .Y(_455_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_449_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_450_) );
OAI21X1 OAI21X1_53 ( .A(_449_), .B(_450_), .C(_20__2_), .Y(_451_) );
NAND2X1 NAND2X1_54 ( .A(_451_), .B(_455_), .Y(_0__26_) );
OAI21X1 OAI21X1_54 ( .A(_452_), .B(_449_), .C(_454_), .Y(_20__3_) );
INVX1 INVX1_28 ( .A(_20__3_), .Y(_459_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_460_) );
NAND2X1 NAND2X1_55 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_461_) );
NAND3X1 NAND3X1_28 ( .A(_459_), .B(_461_), .C(_460_), .Y(_462_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_456_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_457_) );
OAI21X1 OAI21X1_55 ( .A(_456_), .B(_457_), .C(_20__3_), .Y(_458_) );
NAND2X1 NAND2X1_56 ( .A(_458_), .B(_462_), .Y(_0__27_) );
OAI21X1 OAI21X1_56 ( .A(_459_), .B(_456_), .C(_461_), .Y(_19_) );
INVX1 INVX1_29 ( .A(w_cout_7_), .Y(_466_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_467_) );
NAND2X1 NAND2X1_57 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_468_) );
NAND3X1 NAND3X1_29 ( .A(_466_), .B(_468_), .C(_467_), .Y(_469_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_463_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_464_) );
OAI21X1 OAI21X1_57 ( .A(_463_), .B(_464_), .C(w_cout_7_), .Y(_465_) );
NAND2X1 NAND2X1_58 ( .A(_465_), .B(_469_), .Y(_0__28_) );
OAI21X1 OAI21X1_58 ( .A(_466_), .B(_463_), .C(_468_), .Y(_23__1_) );
INVX1 INVX1_30 ( .A(_23__1_), .Y(_473_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_474_) );
NAND2X1 NAND2X1_59 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_475_) );
NAND3X1 NAND3X1_30 ( .A(_473_), .B(_475_), .C(_474_), .Y(_476_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_470_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_471_) );
OAI21X1 OAI21X1_59 ( .A(_470_), .B(_471_), .C(_23__1_), .Y(_472_) );
NAND2X1 NAND2X1_60 ( .A(_472_), .B(_476_), .Y(_0__29_) );
OAI21X1 OAI21X1_60 ( .A(_473_), .B(_470_), .C(_475_), .Y(_23__2_) );
INVX1 INVX1_31 ( .A(_23__2_), .Y(_480_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_481_) );
NAND2X1 NAND2X1_61 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_482_) );
NAND3X1 NAND3X1_31 ( .A(_480_), .B(_482_), .C(_481_), .Y(_483_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_477_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_478_) );
OAI21X1 OAI21X1_61 ( .A(_477_), .B(_478_), .C(_23__2_), .Y(_479_) );
NAND2X1 NAND2X1_62 ( .A(_479_), .B(_483_), .Y(_0__30_) );
OAI21X1 OAI21X1_62 ( .A(_480_), .B(_477_), .C(_482_), .Y(_23__3_) );
INVX1 INVX1_32 ( .A(_23__3_), .Y(_487_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_488_) );
NAND2X1 NAND2X1_63 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_489_) );
NAND3X1 NAND3X1_32 ( .A(_487_), .B(_489_), .C(_488_), .Y(_490_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_484_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_485_) );
OAI21X1 OAI21X1_63 ( .A(_484_), .B(_485_), .C(_23__3_), .Y(_486_) );
NAND2X1 NAND2X1_64 ( .A(_486_), .B(_490_), .Y(_0__31_) );
OAI21X1 OAI21X1_64 ( .A(_487_), .B(_484_), .C(_489_), .Y(_22_) );
INVX1 INVX1_33 ( .A(w_cout_8_), .Y(_494_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_495_) );
NAND2X1 NAND2X1_65 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_496_) );
NAND3X1 NAND3X1_33 ( .A(_494_), .B(_496_), .C(_495_), .Y(_497_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_491_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_492_) );
OAI21X1 OAI21X1_65 ( .A(_491_), .B(_492_), .C(w_cout_8_), .Y(_493_) );
NAND2X1 NAND2X1_66 ( .A(_493_), .B(_497_), .Y(_0__32_) );
OAI21X1 OAI21X1_66 ( .A(_494_), .B(_491_), .C(_496_), .Y(_26__1_) );
INVX1 INVX1_34 ( .A(_26__1_), .Y(_501_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_502_) );
NAND2X1 NAND2X1_67 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_503_) );
NAND3X1 NAND3X1_34 ( .A(_501_), .B(_503_), .C(_502_), .Y(_504_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_498_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_499_) );
OAI21X1 OAI21X1_67 ( .A(_498_), .B(_499_), .C(_26__1_), .Y(_500_) );
NAND2X1 NAND2X1_68 ( .A(_500_), .B(_504_), .Y(_0__33_) );
OAI21X1 OAI21X1_68 ( .A(_501_), .B(_498_), .C(_503_), .Y(_26__2_) );
INVX1 INVX1_35 ( .A(_26__2_), .Y(_508_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_509_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_510_) );
NAND3X1 NAND3X1_35 ( .A(_508_), .B(_510_), .C(_509_), .Y(_511_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_505_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_506_) );
OAI21X1 OAI21X1_69 ( .A(_505_), .B(_506_), .C(_26__2_), .Y(_507_) );
NAND2X1 NAND2X1_70 ( .A(_507_), .B(_511_), .Y(_0__34_) );
OAI21X1 OAI21X1_70 ( .A(_508_), .B(_505_), .C(_510_), .Y(_26__3_) );
INVX1 INVX1_36 ( .A(_26__3_), .Y(_515_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_516_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_517_) );
NAND3X1 NAND3X1_36 ( .A(_515_), .B(_517_), .C(_516_), .Y(_518_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_512_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_513_) );
OAI21X1 OAI21X1_71 ( .A(_512_), .B(_513_), .C(_26__3_), .Y(_514_) );
NAND2X1 NAND2X1_72 ( .A(_514_), .B(_518_), .Y(_0__35_) );
OAI21X1 OAI21X1_72 ( .A(_515_), .B(_512_), .C(_517_), .Y(_25_) );
INVX1 INVX1_37 ( .A(w_cout_9_), .Y(_522_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_523_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_524_) );
NAND3X1 NAND3X1_37 ( .A(_522_), .B(_524_), .C(_523_), .Y(_525_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_519_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_520_) );
OAI21X1 OAI21X1_73 ( .A(_519_), .B(_520_), .C(w_cout_9_), .Y(_521_) );
NAND2X1 NAND2X1_74 ( .A(_521_), .B(_525_), .Y(_0__36_) );
OAI21X1 OAI21X1_74 ( .A(_522_), .B(_519_), .C(_524_), .Y(_29__1_) );
INVX1 INVX1_38 ( .A(_29__1_), .Y(_529_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_530_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_531_) );
NAND3X1 NAND3X1_38 ( .A(_529_), .B(_531_), .C(_530_), .Y(_532_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_526_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_527_) );
OAI21X1 OAI21X1_75 ( .A(_526_), .B(_527_), .C(_29__1_), .Y(_528_) );
NAND2X1 NAND2X1_76 ( .A(_528_), .B(_532_), .Y(_0__37_) );
OAI21X1 OAI21X1_76 ( .A(_529_), .B(_526_), .C(_531_), .Y(_29__2_) );
INVX1 INVX1_39 ( .A(_29__2_), .Y(_536_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_537_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_538_) );
NAND3X1 NAND3X1_39 ( .A(_536_), .B(_538_), .C(_537_), .Y(_539_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_533_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_534_) );
OAI21X1 OAI21X1_77 ( .A(_533_), .B(_534_), .C(_29__2_), .Y(_535_) );
NAND2X1 NAND2X1_78 ( .A(_535_), .B(_539_), .Y(_0__38_) );
OAI21X1 OAI21X1_78 ( .A(_536_), .B(_533_), .C(_538_), .Y(_29__3_) );
INVX1 INVX1_40 ( .A(_29__3_), .Y(_543_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_544_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_545_) );
NAND3X1 NAND3X1_40 ( .A(_543_), .B(_545_), .C(_544_), .Y(_546_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_540_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_541_) );
OAI21X1 OAI21X1_79 ( .A(_540_), .B(_541_), .C(_29__3_), .Y(_542_) );
NAND2X1 NAND2X1_80 ( .A(_542_), .B(_546_), .Y(_0__39_) );
OAI21X1 OAI21X1_80 ( .A(_543_), .B(_540_), .C(_545_), .Y(_28_) );
INVX1 INVX1_41 ( .A(w_cout_10_), .Y(_550_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_551_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_552_) );
NAND3X1 NAND3X1_41 ( .A(_550_), .B(_552_), .C(_551_), .Y(_553_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_547_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_548_) );
OAI21X1 OAI21X1_81 ( .A(_547_), .B(_548_), .C(w_cout_10_), .Y(_549_) );
NAND2X1 NAND2X1_82 ( .A(_549_), .B(_553_), .Y(_0__40_) );
OAI21X1 OAI21X1_82 ( .A(_550_), .B(_547_), .C(_552_), .Y(_32__1_) );
INVX1 INVX1_42 ( .A(_32__1_), .Y(_557_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_558_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_559_) );
NAND3X1 NAND3X1_42 ( .A(_557_), .B(_559_), .C(_558_), .Y(_560_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_554_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_555_) );
OAI21X1 OAI21X1_83 ( .A(_554_), .B(_555_), .C(_32__1_), .Y(_556_) );
NAND2X1 NAND2X1_84 ( .A(_556_), .B(_560_), .Y(_0__41_) );
OAI21X1 OAI21X1_84 ( .A(_557_), .B(_554_), .C(_559_), .Y(_32__2_) );
INVX1 INVX1_43 ( .A(_32__2_), .Y(_564_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_565_) );
NAND2X1 NAND2X1_85 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_566_) );
NAND3X1 NAND3X1_43 ( .A(_564_), .B(_566_), .C(_565_), .Y(_567_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_561_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_562_) );
OAI21X1 OAI21X1_85 ( .A(_561_), .B(_562_), .C(_32__2_), .Y(_563_) );
NAND2X1 NAND2X1_86 ( .A(_563_), .B(_567_), .Y(_0__42_) );
OAI21X1 OAI21X1_86 ( .A(_564_), .B(_561_), .C(_566_), .Y(_32__3_) );
INVX1 INVX1_44 ( .A(_32__3_), .Y(_571_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_572_) );
NAND2X1 NAND2X1_87 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_573_) );
NAND3X1 NAND3X1_44 ( .A(_571_), .B(_573_), .C(_572_), .Y(_574_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_568_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_569_) );
OAI21X1 OAI21X1_87 ( .A(_568_), .B(_569_), .C(_32__3_), .Y(_570_) );
NAND2X1 NAND2X1_88 ( .A(_570_), .B(_574_), .Y(_0__43_) );
OAI21X1 OAI21X1_88 ( .A(_571_), .B(_568_), .C(_573_), .Y(_31_) );
INVX1 INVX1_45 ( .A(w_cout_11_), .Y(_578_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_579_) );
NAND2X1 NAND2X1_89 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_580_) );
NAND3X1 NAND3X1_45 ( .A(_578_), .B(_580_), .C(_579_), .Y(_581_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_575_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_576_) );
OAI21X1 OAI21X1_89 ( .A(_575_), .B(_576_), .C(w_cout_11_), .Y(_577_) );
NAND2X1 NAND2X1_90 ( .A(_577_), .B(_581_), .Y(_0__44_) );
OAI21X1 OAI21X1_90 ( .A(_578_), .B(_575_), .C(_580_), .Y(_35__1_) );
INVX1 INVX1_46 ( .A(_35__1_), .Y(_585_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_586_) );
NAND2X1 NAND2X1_91 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_587_) );
NAND3X1 NAND3X1_46 ( .A(_585_), .B(_587_), .C(_586_), .Y(_588_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_582_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_583_) );
OAI21X1 OAI21X1_91 ( .A(_582_), .B(_583_), .C(_35__1_), .Y(_584_) );
NAND2X1 NAND2X1_92 ( .A(_584_), .B(_588_), .Y(_0__45_) );
OAI21X1 OAI21X1_92 ( .A(_585_), .B(_582_), .C(_587_), .Y(_35__2_) );
INVX1 INVX1_47 ( .A(_35__2_), .Y(_592_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_593_) );
NAND2X1 NAND2X1_93 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_594_) );
NAND3X1 NAND3X1_47 ( .A(_592_), .B(_594_), .C(_593_), .Y(_595_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_589_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_590_) );
OAI21X1 OAI21X1_93 ( .A(_589_), .B(_590_), .C(_35__2_), .Y(_591_) );
NAND2X1 NAND2X1_94 ( .A(_591_), .B(_595_), .Y(_0__46_) );
OAI21X1 OAI21X1_94 ( .A(_592_), .B(_589_), .C(_594_), .Y(_35__3_) );
INVX1 INVX1_48 ( .A(_35__3_), .Y(_599_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_600_) );
NAND2X1 NAND2X1_95 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_601_) );
NAND3X1 NAND3X1_48 ( .A(_599_), .B(_601_), .C(_600_), .Y(_602_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_596_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_597_) );
OAI21X1 OAI21X1_95 ( .A(_596_), .B(_597_), .C(_35__3_), .Y(_598_) );
NAND2X1 NAND2X1_96 ( .A(_598_), .B(_602_), .Y(_0__47_) );
OAI21X1 OAI21X1_96 ( .A(_599_), .B(_596_), .C(_601_), .Y(_34_) );
INVX1 INVX1_49 ( .A(w_cout_12_), .Y(_606_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_607_) );
NAND2X1 NAND2X1_97 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_608_) );
NAND3X1 NAND3X1_49 ( .A(_606_), .B(_608_), .C(_607_), .Y(_609_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_603_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_604_) );
OAI21X1 OAI21X1_97 ( .A(_603_), .B(_604_), .C(w_cout_12_), .Y(_605_) );
NAND2X1 NAND2X1_98 ( .A(_605_), .B(_609_), .Y(_0__48_) );
OAI21X1 OAI21X1_98 ( .A(_606_), .B(_603_), .C(_608_), .Y(_38__1_) );
INVX1 INVX1_50 ( .A(_38__1_), .Y(_613_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_614_) );
NAND2X1 NAND2X1_99 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_615_) );
NAND3X1 NAND3X1_50 ( .A(_613_), .B(_615_), .C(_614_), .Y(_616_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_610_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_611_) );
OAI21X1 OAI21X1_99 ( .A(_610_), .B(_611_), .C(_38__1_), .Y(_612_) );
NAND2X1 NAND2X1_100 ( .A(_612_), .B(_616_), .Y(_0__49_) );
OAI21X1 OAI21X1_100 ( .A(_613_), .B(_610_), .C(_615_), .Y(_38__2_) );
INVX1 INVX1_51 ( .A(_38__2_), .Y(_620_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_621_) );
NAND2X1 NAND2X1_101 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_622_) );
NAND3X1 NAND3X1_51 ( .A(_620_), .B(_622_), .C(_621_), .Y(_623_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_617_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_618_) );
OAI21X1 OAI21X1_101 ( .A(_617_), .B(_618_), .C(_38__2_), .Y(_619_) );
NAND2X1 NAND2X1_102 ( .A(_619_), .B(_623_), .Y(_0__50_) );
OAI21X1 OAI21X1_102 ( .A(_620_), .B(_617_), .C(_622_), .Y(_38__3_) );
INVX1 INVX1_52 ( .A(_38__3_), .Y(_627_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_628_) );
NAND2X1 NAND2X1_103 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_629_) );
NAND3X1 NAND3X1_52 ( .A(_627_), .B(_629_), .C(_628_), .Y(_630_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_624_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_625_) );
OAI21X1 OAI21X1_103 ( .A(_624_), .B(_625_), .C(_38__3_), .Y(_626_) );
NAND2X1 NAND2X1_104 ( .A(_626_), .B(_630_), .Y(_0__51_) );
OAI21X1 OAI21X1_104 ( .A(_627_), .B(_624_), .C(_629_), .Y(_37_) );
INVX1 INVX1_53 ( .A(w_cout_13_), .Y(_634_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_635_) );
NAND2X1 NAND2X1_105 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_636_) );
NAND3X1 NAND3X1_53 ( .A(_634_), .B(_636_), .C(_635_), .Y(_637_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_631_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_632_) );
OAI21X1 OAI21X1_105 ( .A(_631_), .B(_632_), .C(w_cout_13_), .Y(_633_) );
NAND2X1 NAND2X1_106 ( .A(_633_), .B(_637_), .Y(_0__52_) );
OAI21X1 OAI21X1_106 ( .A(_634_), .B(_631_), .C(_636_), .Y(_41__1_) );
INVX1 INVX1_54 ( .A(_41__1_), .Y(_641_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_642_) );
NAND2X1 NAND2X1_107 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_643_) );
NAND3X1 NAND3X1_54 ( .A(_641_), .B(_643_), .C(_642_), .Y(_644_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_638_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_639_) );
OAI21X1 OAI21X1_107 ( .A(_638_), .B(_639_), .C(_41__1_), .Y(_640_) );
NAND2X1 NAND2X1_108 ( .A(_640_), .B(_644_), .Y(_0__53_) );
OAI21X1 OAI21X1_108 ( .A(_641_), .B(_638_), .C(_643_), .Y(_41__2_) );
INVX1 INVX1_55 ( .A(_41__2_), .Y(_648_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_649_) );
NAND2X1 NAND2X1_109 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_650_) );
NAND3X1 NAND3X1_55 ( .A(_648_), .B(_650_), .C(_649_), .Y(_651_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_645_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_646_) );
OAI21X1 OAI21X1_109 ( .A(_645_), .B(_646_), .C(_41__2_), .Y(_647_) );
NAND2X1 NAND2X1_110 ( .A(_647_), .B(_651_), .Y(_0__54_) );
OAI21X1 OAI21X1_110 ( .A(_648_), .B(_645_), .C(_650_), .Y(_41__3_) );
INVX1 INVX1_56 ( .A(_41__3_), .Y(_655_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_656_) );
NAND2X1 NAND2X1_111 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_657_) );
NAND3X1 NAND3X1_56 ( .A(_655_), .B(_657_), .C(_656_), .Y(_658_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_652_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_653_) );
OAI21X1 OAI21X1_111 ( .A(_652_), .B(_653_), .C(_41__3_), .Y(_654_) );
NAND2X1 NAND2X1_112 ( .A(_654_), .B(_658_), .Y(_0__55_) );
OAI21X1 OAI21X1_112 ( .A(_655_), .B(_652_), .C(_657_), .Y(_40_) );
INVX1 INVX1_57 ( .A(cskip2_inst_cin), .Y(_662_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_663_) );
NAND2X1 NAND2X1_113 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_664_) );
NAND3X1 NAND3X1_57 ( .A(_662_), .B(_664_), .C(_663_), .Y(_665_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_659_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_660_) );
OAI21X1 OAI21X1_113 ( .A(_659_), .B(_660_), .C(cskip2_inst_cin), .Y(_661_) );
NAND2X1 NAND2X1_114 ( .A(_661_), .B(_665_), .Y(_0__56_) );
OAI21X1 OAI21X1_114 ( .A(_662_), .B(_659_), .C(_664_), .Y(cskip2_inst_rca0_w_CARRY_1_) );
INVX1 INVX1_58 ( .A(cskip2_inst_rca0_w_CARRY_1_), .Y(_669_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_670_) );
NAND2X1 NAND2X1_115 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_671_) );
NAND3X1 NAND3X1_58 ( .A(_669_), .B(_671_), .C(_670_), .Y(_672_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_666_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_667_) );
OAI21X1 OAI21X1_115 ( .A(_666_), .B(_667_), .C(cskip2_inst_rca0_w_CARRY_1_), .Y(_668_) );
NAND2X1 NAND2X1_116 ( .A(_668_), .B(_672_), .Y(_0__57_) );
OAI21X1 OAI21X1_116 ( .A(_669_), .B(_666_), .C(_671_), .Y(cskip2_inst_rca0_w_CARRY_2_) );
INVX1 INVX1_59 ( .A(cskip2_inst_rca0_w_CARRY_2_), .Y(_674_) );
NAND2X1 NAND2X1_117 ( .A(gnd), .B(gnd), .Y(_675_) );
NOR2X1 NOR2X1_59 ( .A(gnd), .B(gnd), .Y(_673_) );
OAI21X1 OAI21X1_117 ( .A(_674_), .B(_673_), .C(_675_), .Y(cskip2_inst_rca0_w_CARRY_3_) );
INVX1 INVX1_60 ( .A(cskip2_inst_rca0_w_CARRY_3_), .Y(_677_) );
NAND2X1 NAND2X1_118 ( .A(gnd), .B(gnd), .Y(_678_) );
NOR2X1 NOR2X1_60 ( .A(gnd), .B(gnd), .Y(_676_) );
OAI21X1 OAI21X1_118 ( .A(_677_), .B(_676_), .C(_678_), .Y(cskip2_inst_cout0) );
INVX1 INVX1_61 ( .A(i_add_term1[57]), .Y(_683_) );
NAND2X1 NAND2X1_119 ( .A(i_add_term2[57]), .B(_683_), .Y(_684_) );
INVX1 INVX1_62 ( .A(i_add_term2[57]), .Y(_685_) );
NAND2X1 NAND2X1_120 ( .A(i_add_term1[57]), .B(_685_), .Y(_686_) );
INVX1 INVX1_63 ( .A(i_add_term1[56]), .Y(_679_) );
NAND2X1 NAND2X1_121 ( .A(i_add_term2[56]), .B(_679_), .Y(_680_) );
INVX1 INVX1_64 ( .A(i_add_term2[56]), .Y(_681_) );
NAND2X1 NAND2X1_122 ( .A(i_add_term1[56]), .B(_681_), .Y(_682_) );
AOI22X1 AOI22X1_1 ( .A(_684_), .B(_686_), .C(_680_), .D(_682_), .Y(cskip2_inst_skip0_P) );
INVX1 INVX1_65 ( .A(cskip2_inst_cout0), .Y(_687_) );
NAND2X1 NAND2X1_123 ( .A(gnd), .B(cskip2_inst_skip0_P), .Y(_688_) );
OAI21X1 OAI21X1_119 ( .A(cskip2_inst_skip0_P), .B(_687_), .C(_688_), .Y(w_cout_15_) );
BUFX2 BUFX2_1 ( .A(w_cout_15_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_0__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_0__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_0__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_0__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .A(_0__54_), .Y(sum[54]) );
BUFX2 BUFX2_57 ( .A(_0__55_), .Y(sum[55]) );
BUFX2 BUFX2_58 ( .A(_0__56_), .Y(sum[56]) );
BUFX2 BUFX2_59 ( .A(_0__57_), .Y(sum[57]) );
INVX1 INVX1_66 ( .A(i_add_term1[0]), .Y(_43_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[0]), .B(_43_), .Y(_44_) );
INVX1 INVX1_67 ( .A(i_add_term2[0]), .Y(_45_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term1[0]), .B(_45_), .Y(_46_) );
INVX1 INVX1_68 ( .A(i_add_term1[1]), .Y(_47_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[1]), .B(_47_), .Y(_48_) );
INVX1 INVX1_69 ( .A(i_add_term2[1]), .Y(_49_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term1[1]), .B(_49_), .Y(_50_) );
OAI22X1 OAI22X1_1 ( .A(_44_), .B(_46_), .C(_48_), .D(_50_), .Y(_51_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_52_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_53_) );
NOR2X1 NOR2X1_66 ( .A(_52_), .B(_53_), .Y(_54_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_55_) );
NAND2X1 NAND2X1_124 ( .A(_54_), .B(_55_), .Y(_56_) );
NOR2X1 NOR2X1_67 ( .A(_51_), .B(_56_), .Y(_3_) );
INVX1 INVX1_70 ( .A(_1_), .Y(_57_) );
NAND2X1 NAND2X1_125 ( .A(gnd), .B(_3_), .Y(_58_) );
OAI21X1 OAI21X1_120 ( .A(_3_), .B(_57_), .C(_58_), .Y(w_cout_1_) );
INVX1 INVX1_71 ( .A(i_add_term1[4]), .Y(_59_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[4]), .B(_59_), .Y(_60_) );
INVX1 INVX1_72 ( .A(i_add_term2[4]), .Y(_61_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term1[4]), .B(_61_), .Y(_62_) );
INVX1 INVX1_73 ( .A(i_add_term1[5]), .Y(_63_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[5]), .B(_63_), .Y(_64_) );
INVX1 INVX1_74 ( .A(i_add_term2[5]), .Y(_65_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term1[5]), .B(_65_), .Y(_66_) );
OAI22X1 OAI22X1_2 ( .A(_60_), .B(_62_), .C(_64_), .D(_66_), .Y(_67_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_68_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_69_) );
NOR2X1 NOR2X1_73 ( .A(_68_), .B(_69_), .Y(_70_) );
XOR2X1 XOR2X1_2 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_71_) );
NAND2X1 NAND2X1_126 ( .A(_70_), .B(_71_), .Y(_72_) );
NOR2X1 NOR2X1_74 ( .A(_67_), .B(_72_), .Y(_6_) );
INVX1 INVX1_75 ( .A(_4_), .Y(_73_) );
NAND2X1 NAND2X1_127 ( .A(gnd), .B(_6_), .Y(_74_) );
OAI21X1 OAI21X1_121 ( .A(_6_), .B(_73_), .C(_74_), .Y(w_cout_2_) );
INVX1 INVX1_76 ( .A(i_add_term1[8]), .Y(_75_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[8]), .B(_75_), .Y(_76_) );
INVX1 INVX1_77 ( .A(i_add_term2[8]), .Y(_77_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term1[8]), .B(_77_), .Y(_78_) );
INVX1 INVX1_78 ( .A(i_add_term1[9]), .Y(_79_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[9]), .B(_79_), .Y(_80_) );
INVX1 INVX1_79 ( .A(i_add_term2[9]), .Y(_81_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term1[9]), .B(_81_), .Y(_82_) );
OAI22X1 OAI22X1_3 ( .A(_76_), .B(_78_), .C(_80_), .D(_82_), .Y(_83_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_84_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_85_) );
NOR2X1 NOR2X1_80 ( .A(_84_), .B(_85_), .Y(_86_) );
XOR2X1 XOR2X1_3 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_87_) );
NAND2X1 NAND2X1_128 ( .A(_86_), .B(_87_), .Y(_88_) );
NOR2X1 NOR2X1_81 ( .A(_83_), .B(_88_), .Y(_9_) );
INVX1 INVX1_80 ( .A(_7_), .Y(_89_) );
NAND2X1 NAND2X1_129 ( .A(gnd), .B(_9_), .Y(_90_) );
OAI21X1 OAI21X1_122 ( .A(_9_), .B(_89_), .C(_90_), .Y(w_cout_3_) );
INVX1 INVX1_81 ( .A(i_add_term1[12]), .Y(_91_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[12]), .B(_91_), .Y(_92_) );
INVX1 INVX1_82 ( .A(i_add_term2[12]), .Y(_93_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term1[12]), .B(_93_), .Y(_94_) );
INVX1 INVX1_83 ( .A(i_add_term1[13]), .Y(_95_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[13]), .B(_95_), .Y(_96_) );
INVX1 INVX1_84 ( .A(i_add_term2[13]), .Y(_97_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term1[13]), .B(_97_), .Y(_98_) );
OAI22X1 OAI22X1_4 ( .A(_92_), .B(_94_), .C(_96_), .D(_98_), .Y(_99_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_100_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_101_) );
NOR2X1 NOR2X1_87 ( .A(_100_), .B(_101_), .Y(_102_) );
XOR2X1 XOR2X1_4 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_103_) );
NAND2X1 NAND2X1_130 ( .A(_102_), .B(_103_), .Y(_104_) );
NOR2X1 NOR2X1_88 ( .A(_99_), .B(_104_), .Y(_12_) );
INVX1 INVX1_85 ( .A(_10_), .Y(_105_) );
NAND2X1 NAND2X1_131 ( .A(gnd), .B(_12_), .Y(_106_) );
OAI21X1 OAI21X1_123 ( .A(_12_), .B(_105_), .C(_106_), .Y(w_cout_4_) );
INVX1 INVX1_86 ( .A(i_add_term1[16]), .Y(_107_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[16]), .B(_107_), .Y(_108_) );
INVX1 INVX1_87 ( .A(i_add_term2[16]), .Y(_109_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term1[16]), .B(_109_), .Y(_110_) );
INVX1 INVX1_88 ( .A(i_add_term1[17]), .Y(_111_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[17]), .B(_111_), .Y(_112_) );
INVX1 INVX1_89 ( .A(i_add_term2[17]), .Y(_113_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term1[17]), .B(_113_), .Y(_114_) );
OAI22X1 OAI22X1_5 ( .A(_108_), .B(_110_), .C(_112_), .D(_114_), .Y(_115_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_116_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_117_) );
NOR2X1 NOR2X1_94 ( .A(_116_), .B(_117_), .Y(_118_) );
XOR2X1 XOR2X1_5 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_119_) );
NAND2X1 NAND2X1_132 ( .A(_118_), .B(_119_), .Y(_120_) );
NOR2X1 NOR2X1_95 ( .A(_115_), .B(_120_), .Y(_15_) );
INVX1 INVX1_90 ( .A(_13_), .Y(_121_) );
NAND2X1 NAND2X1_133 ( .A(gnd), .B(_15_), .Y(_122_) );
OAI21X1 OAI21X1_124 ( .A(_15_), .B(_121_), .C(_122_), .Y(w_cout_5_) );
INVX1 INVX1_91 ( .A(i_add_term1[20]), .Y(_123_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[20]), .B(_123_), .Y(_124_) );
INVX1 INVX1_92 ( .A(i_add_term2[20]), .Y(_125_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term1[20]), .B(_125_), .Y(_126_) );
INVX1 INVX1_93 ( .A(i_add_term1[21]), .Y(_127_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[21]), .B(_127_), .Y(_128_) );
INVX1 INVX1_94 ( .A(i_add_term2[21]), .Y(_129_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term1[21]), .B(_129_), .Y(_130_) );
OAI22X1 OAI22X1_6 ( .A(_124_), .B(_126_), .C(_128_), .D(_130_), .Y(_131_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_132_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_133_) );
NOR2X1 NOR2X1_101 ( .A(_132_), .B(_133_), .Y(_134_) );
XOR2X1 XOR2X1_6 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_135_) );
NAND2X1 NAND2X1_134 ( .A(_134_), .B(_135_), .Y(_136_) );
NOR2X1 NOR2X1_102 ( .A(_131_), .B(_136_), .Y(_18_) );
INVX1 INVX1_95 ( .A(_16_), .Y(_137_) );
NAND2X1 NAND2X1_135 ( .A(gnd), .B(_18_), .Y(_138_) );
OAI21X1 OAI21X1_125 ( .A(_18_), .B(_137_), .C(_138_), .Y(w_cout_6_) );
INVX1 INVX1_96 ( .A(i_add_term1[24]), .Y(_139_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[24]), .B(_139_), .Y(_140_) );
INVX1 INVX1_97 ( .A(i_add_term2[24]), .Y(_141_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term1[24]), .B(_141_), .Y(_142_) );
INVX1 INVX1_98 ( .A(i_add_term1[25]), .Y(_143_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[25]), .B(_143_), .Y(_144_) );
INVX1 INVX1_99 ( .A(i_add_term2[25]), .Y(_145_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term1[25]), .B(_145_), .Y(_146_) );
OAI22X1 OAI22X1_7 ( .A(_140_), .B(_142_), .C(_144_), .D(_146_), .Y(_147_) );
NOR2X1 NOR2X1_107 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_148_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_149_) );
NOR2X1 NOR2X1_108 ( .A(_148_), .B(_149_), .Y(_150_) );
XOR2X1 XOR2X1_7 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_151_) );
NAND2X1 NAND2X1_136 ( .A(_150_), .B(_151_), .Y(_152_) );
NOR2X1 NOR2X1_109 ( .A(_147_), .B(_152_), .Y(_21_) );
INVX1 INVX1_100 ( .A(_19_), .Y(_153_) );
NAND2X1 NAND2X1_137 ( .A(gnd), .B(_21_), .Y(_154_) );
OAI21X1 OAI21X1_126 ( .A(_21_), .B(_153_), .C(_154_), .Y(w_cout_7_) );
INVX1 INVX1_101 ( .A(i_add_term1[28]), .Y(_155_) );
NOR2X1 NOR2X1_110 ( .A(i_add_term2[28]), .B(_155_), .Y(_156_) );
INVX1 INVX1_102 ( .A(i_add_term2[28]), .Y(_157_) );
NOR2X1 NOR2X1_111 ( .A(i_add_term1[28]), .B(_157_), .Y(_158_) );
INVX1 INVX1_103 ( .A(i_add_term1[29]), .Y(_159_) );
NOR2X1 NOR2X1_112 ( .A(i_add_term2[29]), .B(_159_), .Y(_160_) );
INVX1 INVX1_104 ( .A(i_add_term2[29]), .Y(_161_) );
NOR2X1 NOR2X1_113 ( .A(i_add_term1[29]), .B(_161_), .Y(_162_) );
OAI22X1 OAI22X1_8 ( .A(_156_), .B(_158_), .C(_160_), .D(_162_), .Y(_163_) );
NOR2X1 NOR2X1_114 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_164_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_165_) );
NOR2X1 NOR2X1_115 ( .A(_164_), .B(_165_), .Y(_166_) );
XOR2X1 XOR2X1_8 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_167_) );
NAND2X1 NAND2X1_138 ( .A(_166_), .B(_167_), .Y(_168_) );
NOR2X1 NOR2X1_116 ( .A(_163_), .B(_168_), .Y(_24_) );
INVX1 INVX1_105 ( .A(_22_), .Y(_169_) );
NAND2X1 NAND2X1_139 ( .A(gnd), .B(_24_), .Y(_170_) );
OAI21X1 OAI21X1_127 ( .A(_24_), .B(_169_), .C(_170_), .Y(w_cout_8_) );
INVX1 INVX1_106 ( .A(i_add_term1[32]), .Y(_171_) );
NOR2X1 NOR2X1_117 ( .A(i_add_term2[32]), .B(_171_), .Y(_172_) );
INVX1 INVX1_107 ( .A(i_add_term2[32]), .Y(_173_) );
NOR2X1 NOR2X1_118 ( .A(i_add_term1[32]), .B(_173_), .Y(_174_) );
INVX1 INVX1_108 ( .A(i_add_term1[33]), .Y(_175_) );
NOR2X1 NOR2X1_119 ( .A(i_add_term2[33]), .B(_175_), .Y(_176_) );
INVX1 INVX1_109 ( .A(i_add_term2[33]), .Y(_177_) );
NOR2X1 NOR2X1_120 ( .A(i_add_term1[33]), .B(_177_), .Y(_178_) );
OAI22X1 OAI22X1_9 ( .A(_172_), .B(_174_), .C(_176_), .D(_178_), .Y(_179_) );
NOR2X1 NOR2X1_121 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_180_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_181_) );
NOR2X1 NOR2X1_122 ( .A(_180_), .B(_181_), .Y(_182_) );
XOR2X1 XOR2X1_9 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_183_) );
NAND2X1 NAND2X1_140 ( .A(_182_), .B(_183_), .Y(_184_) );
NOR2X1 NOR2X1_123 ( .A(_179_), .B(_184_), .Y(_27_) );
INVX1 INVX1_110 ( .A(_25_), .Y(_185_) );
NAND2X1 NAND2X1_141 ( .A(gnd), .B(_27_), .Y(_186_) );
OAI21X1 OAI21X1_128 ( .A(_27_), .B(_185_), .C(_186_), .Y(w_cout_9_) );
INVX1 INVX1_111 ( .A(i_add_term1[36]), .Y(_187_) );
NOR2X1 NOR2X1_124 ( .A(i_add_term2[36]), .B(_187_), .Y(_188_) );
INVX1 INVX1_112 ( .A(i_add_term2[36]), .Y(_189_) );
NOR2X1 NOR2X1_125 ( .A(i_add_term1[36]), .B(_189_), .Y(_190_) );
INVX1 INVX1_113 ( .A(i_add_term1[37]), .Y(_191_) );
NOR2X1 NOR2X1_126 ( .A(i_add_term2[37]), .B(_191_), .Y(_192_) );
INVX1 INVX1_114 ( .A(i_add_term2[37]), .Y(_193_) );
NOR2X1 NOR2X1_127 ( .A(i_add_term1[37]), .B(_193_), .Y(_194_) );
OAI22X1 OAI22X1_10 ( .A(_188_), .B(_190_), .C(_192_), .D(_194_), .Y(_195_) );
NOR2X1 NOR2X1_128 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_196_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_197_) );
NOR2X1 NOR2X1_129 ( .A(_196_), .B(_197_), .Y(_198_) );
XOR2X1 XOR2X1_10 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_199_) );
NAND2X1 NAND2X1_142 ( .A(_198_), .B(_199_), .Y(_200_) );
NOR2X1 NOR2X1_130 ( .A(_195_), .B(_200_), .Y(_30_) );
INVX1 INVX1_115 ( .A(_28_), .Y(_201_) );
NAND2X1 NAND2X1_143 ( .A(gnd), .B(_30_), .Y(_202_) );
OAI21X1 OAI21X1_129 ( .A(_30_), .B(_201_), .C(_202_), .Y(w_cout_10_) );
INVX1 INVX1_116 ( .A(i_add_term1[40]), .Y(_203_) );
NOR2X1 NOR2X1_131 ( .A(i_add_term2[40]), .B(_203_), .Y(_204_) );
INVX1 INVX1_117 ( .A(i_add_term2[40]), .Y(_205_) );
NOR2X1 NOR2X1_132 ( .A(i_add_term1[40]), .B(_205_), .Y(_206_) );
INVX1 INVX1_118 ( .A(i_add_term1[41]), .Y(_207_) );
NOR2X1 NOR2X1_133 ( .A(i_add_term2[41]), .B(_207_), .Y(_208_) );
INVX1 INVX1_119 ( .A(i_add_term2[41]), .Y(_209_) );
NOR2X1 NOR2X1_134 ( .A(i_add_term1[41]), .B(_209_), .Y(_210_) );
OAI22X1 OAI22X1_11 ( .A(_204_), .B(_206_), .C(_208_), .D(_210_), .Y(_211_) );
NOR2X1 NOR2X1_135 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_212_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_213_) );
NOR2X1 NOR2X1_136 ( .A(_212_), .B(_213_), .Y(_214_) );
XOR2X1 XOR2X1_11 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_215_) );
NAND2X1 NAND2X1_144 ( .A(_214_), .B(_215_), .Y(_216_) );
NOR2X1 NOR2X1_137 ( .A(_211_), .B(_216_), .Y(_33_) );
INVX1 INVX1_120 ( .A(_31_), .Y(_217_) );
NAND2X1 NAND2X1_145 ( .A(gnd), .B(_33_), .Y(_218_) );
OAI21X1 OAI21X1_130 ( .A(_33_), .B(_217_), .C(_218_), .Y(w_cout_11_) );
INVX1 INVX1_121 ( .A(i_add_term1[44]), .Y(_219_) );
NOR2X1 NOR2X1_138 ( .A(i_add_term2[44]), .B(_219_), .Y(_220_) );
INVX1 INVX1_122 ( .A(i_add_term2[44]), .Y(_221_) );
NOR2X1 NOR2X1_139 ( .A(i_add_term1[44]), .B(_221_), .Y(_222_) );
INVX1 INVX1_123 ( .A(i_add_term1[45]), .Y(_223_) );
NOR2X1 NOR2X1_140 ( .A(i_add_term2[45]), .B(_223_), .Y(_224_) );
INVX1 INVX1_124 ( .A(i_add_term2[45]), .Y(_225_) );
NOR2X1 NOR2X1_141 ( .A(i_add_term1[45]), .B(_225_), .Y(_226_) );
OAI22X1 OAI22X1_12 ( .A(_220_), .B(_222_), .C(_224_), .D(_226_), .Y(_227_) );
NOR2X1 NOR2X1_142 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_228_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_229_) );
NOR2X1 NOR2X1_143 ( .A(_228_), .B(_229_), .Y(_230_) );
XOR2X1 XOR2X1_12 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_231_) );
NAND2X1 NAND2X1_146 ( .A(_230_), .B(_231_), .Y(_232_) );
NOR2X1 NOR2X1_144 ( .A(_227_), .B(_232_), .Y(_36_) );
INVX1 INVX1_125 ( .A(_34_), .Y(_233_) );
NAND2X1 NAND2X1_147 ( .A(gnd), .B(_36_), .Y(_234_) );
OAI21X1 OAI21X1_131 ( .A(_36_), .B(_233_), .C(_234_), .Y(w_cout_12_) );
INVX1 INVX1_126 ( .A(i_add_term1[48]), .Y(_235_) );
NOR2X1 NOR2X1_145 ( .A(i_add_term2[48]), .B(_235_), .Y(_236_) );
INVX1 INVX1_127 ( .A(i_add_term2[48]), .Y(_237_) );
NOR2X1 NOR2X1_146 ( .A(i_add_term1[48]), .B(_237_), .Y(_238_) );
INVX1 INVX1_128 ( .A(i_add_term1[49]), .Y(_239_) );
NOR2X1 NOR2X1_147 ( .A(i_add_term2[49]), .B(_239_), .Y(_240_) );
INVX1 INVX1_129 ( .A(i_add_term2[49]), .Y(_241_) );
NOR2X1 NOR2X1_148 ( .A(i_add_term1[49]), .B(_241_), .Y(_242_) );
OAI22X1 OAI22X1_13 ( .A(_236_), .B(_238_), .C(_240_), .D(_242_), .Y(_243_) );
NOR2X1 NOR2X1_149 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_244_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_245_) );
NOR2X1 NOR2X1_150 ( .A(_244_), .B(_245_), .Y(_246_) );
XOR2X1 XOR2X1_13 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_247_) );
NAND2X1 NAND2X1_148 ( .A(_246_), .B(_247_), .Y(_248_) );
NOR2X1 NOR2X1_151 ( .A(_243_), .B(_248_), .Y(_39_) );
INVX1 INVX1_130 ( .A(_37_), .Y(_249_) );
NAND2X1 NAND2X1_149 ( .A(gnd), .B(_39_), .Y(_250_) );
OAI21X1 OAI21X1_132 ( .A(_39_), .B(_249_), .C(_250_), .Y(w_cout_13_) );
INVX1 INVX1_131 ( .A(i_add_term1[52]), .Y(_251_) );
NOR2X1 NOR2X1_152 ( .A(i_add_term2[52]), .B(_251_), .Y(_252_) );
INVX1 INVX1_132 ( .A(i_add_term2[52]), .Y(_253_) );
NOR2X1 NOR2X1_153 ( .A(i_add_term1[52]), .B(_253_), .Y(_254_) );
INVX1 INVX1_133 ( .A(i_add_term1[53]), .Y(_255_) );
NOR2X1 NOR2X1_154 ( .A(i_add_term2[53]), .B(_255_), .Y(_256_) );
INVX1 INVX1_134 ( .A(i_add_term2[53]), .Y(_257_) );
NOR2X1 NOR2X1_155 ( .A(i_add_term1[53]), .B(_257_), .Y(_258_) );
OAI22X1 OAI22X1_14 ( .A(_252_), .B(_254_), .C(_256_), .D(_258_), .Y(_259_) );
NOR2X1 NOR2X1_156 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_260_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_261_) );
NOR2X1 NOR2X1_157 ( .A(_260_), .B(_261_), .Y(_262_) );
XOR2X1 XOR2X1_14 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_263_) );
NAND2X1 NAND2X1_150 ( .A(_262_), .B(_263_), .Y(_264_) );
NOR2X1 NOR2X1_158 ( .A(_259_), .B(_264_), .Y(_42_) );
INVX1 INVX1_135 ( .A(_40_), .Y(_265_) );
NAND2X1 NAND2X1_151 ( .A(gnd), .B(_42_), .Y(_266_) );
OAI21X1 OAI21X1_133 ( .A(_42_), .B(_265_), .C(_266_), .Y(cskip2_inst_cin) );
BUFX2 BUFX2_60 ( .A(gnd), .Y(_2__0_) );
BUFX2 BUFX2_61 ( .A(_1_), .Y(_2__4_) );
BUFX2 BUFX2_62 ( .A(w_cout_1_), .Y(_5__0_) );
BUFX2 BUFX2_63 ( .A(_4_), .Y(_5__4_) );
BUFX2 BUFX2_64 ( .A(w_cout_2_), .Y(_8__0_) );
BUFX2 BUFX2_65 ( .A(_7_), .Y(_8__4_) );
BUFX2 BUFX2_66 ( .A(w_cout_3_), .Y(_11__0_) );
BUFX2 BUFX2_67 ( .A(_10_), .Y(_11__4_) );
BUFX2 BUFX2_68 ( .A(w_cout_4_), .Y(_14__0_) );
BUFX2 BUFX2_69 ( .A(_13_), .Y(_14__4_) );
BUFX2 BUFX2_70 ( .A(w_cout_5_), .Y(_17__0_) );
BUFX2 BUFX2_71 ( .A(_16_), .Y(_17__4_) );
BUFX2 BUFX2_72 ( .A(w_cout_6_), .Y(_20__0_) );
BUFX2 BUFX2_73 ( .A(_19_), .Y(_20__4_) );
BUFX2 BUFX2_74 ( .A(w_cout_7_), .Y(_23__0_) );
BUFX2 BUFX2_75 ( .A(_22_), .Y(_23__4_) );
BUFX2 BUFX2_76 ( .A(w_cout_8_), .Y(_26__0_) );
BUFX2 BUFX2_77 ( .A(_25_), .Y(_26__4_) );
BUFX2 BUFX2_78 ( .A(w_cout_9_), .Y(_29__0_) );
BUFX2 BUFX2_79 ( .A(_28_), .Y(_29__4_) );
BUFX2 BUFX2_80 ( .A(w_cout_10_), .Y(_32__0_) );
BUFX2 BUFX2_81 ( .A(_31_), .Y(_32__4_) );
BUFX2 BUFX2_82 ( .A(w_cout_11_), .Y(_35__0_) );
BUFX2 BUFX2_83 ( .A(_34_), .Y(_35__4_) );
BUFX2 BUFX2_84 ( .A(w_cout_12_), .Y(_38__0_) );
BUFX2 BUFX2_85 ( .A(_37_), .Y(_38__4_) );
BUFX2 BUFX2_86 ( .A(w_cout_13_), .Y(_41__0_) );
BUFX2 BUFX2_87 ( .A(_40_), .Y(_41__4_) );
BUFX2 BUFX2_88 ( .A(cskip2_inst_cin), .Y(cskip2_inst_rca0_w_CARRY_0_) );
BUFX2 BUFX2_89 ( .A(cskip2_inst_cout0), .Y(cskip2_inst_rca0_w_CARRY_4_) );
BUFX2 BUFX2_90 ( .A(gnd), .Y(w_cout_0_) );
BUFX2 BUFX2_91 ( .A(cskip2_inst_cin), .Y(w_cout_14_) );
endmodule
