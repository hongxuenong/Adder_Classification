module CSkipA_6bit (i_add_term1[0], i_add_term1[1], i_add_term1[2], i_add_term1[3], i_add_term1[4], i_add_term1[5], i_add_term2[0], i_add_term2[1], i_add_term2[2], i_add_term2[3], i_add_term2[4], i_add_term2[5], sum[0], sum[1], sum[2], sum[3], sum[4], sum[5], cout);

input i_add_term1[0];
input i_add_term1[1];
input i_add_term1[2];
input i_add_term1[3];
input i_add_term1[4];
input i_add_term1[5];
input i_add_term2[0];
input i_add_term2[1];
input i_add_term2[2];
input i_add_term2[3];
input i_add_term2[4];
input i_add_term2[5];
output sum[0];
output sum[1];
output sum[2];
output sum[3];
output sum[4];
output sum[5];
output cout;

NAND2X1 NAND2X1_1 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_24_) );
NAND3X1 NAND3X1_1 ( .A(_22_), .B(_24_), .C(_23_), .Y(_25_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_19_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_20_) );
OAI21X1 OAI21X1_1 ( .A(_19_), .B(_20_), .C(_3__1_), .Y(_21_) );
NAND2X1 NAND2X1_2 ( .A(_21_), .B(_25_), .Y(_1__1_) );
OAI21X1 OAI21X1_2 ( .A(_22_), .B(_19_), .C(_24_), .Y(_3__2_) );
INVX1 INVX1_1 ( .A(_3__2_), .Y(_29_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_30_) );
NAND2X1 NAND2X1_3 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_31_) );
NAND3X1 NAND3X1_2 ( .A(_29_), .B(_31_), .C(_30_), .Y(_32_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_26_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_27_) );
OAI21X1 OAI21X1_3 ( .A(_26_), .B(_27_), .C(_3__2_), .Y(_28_) );
NAND2X1 NAND2X1_4 ( .A(_28_), .B(_32_), .Y(_1__2_) );
OAI21X1 OAI21X1_4 ( .A(_29_), .B(_26_), .C(_31_), .Y(_3__3_) );
INVX1 INVX1_2 ( .A(i_add_term1[0]), .Y(_33_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[0]), .B(_33_), .Y(_34_) );
INVX1 INVX1_3 ( .A(i_add_term2[0]), .Y(_35_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term1[0]), .B(_35_), .Y(_36_) );
INVX1 INVX1_4 ( .A(i_add_term1[1]), .Y(_37_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[1]), .B(_37_), .Y(_38_) );
INVX1 INVX1_5 ( .A(i_add_term2[1]), .Y(_39_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term1[1]), .B(_39_), .Y(_40_) );
OAI22X1 OAI22X1_1 ( .A(_34_), .B(_36_), .C(_38_), .D(_40_), .Y(_41_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_42_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_43_) );
NOR2X1 NOR2X1_8 ( .A(_42_), .B(_43_), .Y(_44_) );
XOR2X1 XOR2X1_1 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_45_) );
NAND2X1 NAND2X1_5 ( .A(_44_), .B(_45_), .Y(_46_) );
NOR2X1 NOR2X1_9 ( .A(_41_), .B(_46_), .Y(_4_) );
INVX1 INVX1_6 ( .A(_2_), .Y(_47_) );
NAND2X1 NAND2X1_6 ( .A(1'b0), .B(_4_), .Y(_48_) );
OAI21X1 OAI21X1_5 ( .A(_4_), .B(_47_), .C(_48_), .Y(cskip2_inst_cin) );
INVX1 INVX1_7 ( .A(cskip2_inst_cin), .Y(_52_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_53_) );
NAND2X1 NAND2X1_7 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_54_) );
NAND3X1 NAND3X1_3 ( .A(_52_), .B(_54_), .C(_53_), .Y(_55_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_49_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_50_) );
OAI21X1 OAI21X1_6 ( .A(_49_), .B(_50_), .C(cskip2_inst_cin), .Y(_51_) );
NAND2X1 NAND2X1_8 ( .A(_51_), .B(_55_), .Y(cskip2_inst_rca0_fa0_o_sum) );
OAI21X1 OAI21X1_7 ( .A(_52_), .B(_49_), .C(_54_), .Y(cskip2_inst_rca0_c) );
INVX1 INVX1_8 ( .A(cskip2_inst_rca0_c), .Y(_59_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_60_) );
NAND2X1 NAND2X1_9 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_61_) );
NAND3X1 NAND3X1_4 ( .A(_59_), .B(_61_), .C(_60_), .Y(_62_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_56_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_57_) );
OAI21X1 OAI21X1_8 ( .A(_56_), .B(_57_), .C(cskip2_inst_rca0_c), .Y(_58_) );
NAND2X1 NAND2X1_10 ( .A(_58_), .B(_62_), .Y(cskip2_inst_rca0_fa31_o_sum) );
OAI21X1 OAI21X1_9 ( .A(_59_), .B(_56_), .C(_61_), .Y(cskip2_inst_cout0) );
INVX1 INVX1_9 ( .A(i_add_term1[5]), .Y(_67_) );
NAND2X1 NAND2X1_11 ( .A(i_add_term2[5]), .B(_67_), .Y(_68_) );
INVX1 INVX1_10 ( .A(i_add_term2[5]), .Y(_69_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term1[5]), .B(_69_), .Y(_70_) );
INVX1 INVX1_11 ( .A(i_add_term1[4]), .Y(_63_) );
NAND2X1 NAND2X1_13 ( .A(i_add_term2[4]), .B(_63_), .Y(_64_) );
INVX1 INVX1_12 ( .A(i_add_term2[4]), .Y(_65_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term1[4]), .B(_65_), .Y(_66_) );
AOI22X1 AOI22X1_1 ( .A(_68_), .B(_70_), .C(_64_), .D(_66_), .Y(cskip2_inst_skip0_P) );
INVX1 INVX1_13 ( .A(cskip2_inst_cout0), .Y(_71_) );
NAND2X1 NAND2X1_15 ( .A(1'b0), .B(cskip2_inst_skip0_P), .Y(_72_) );
OAI21X1 OAI21X1_10 ( .A(cskip2_inst_skip0_P), .B(_71_), .C(_72_), .Y(_0_) );
BUFX2 BUFX2_1 ( .A(_0_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(_1__0_), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(_1__1_), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(_1__2_), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(_1__3_), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(cskip2_inst_rca0_fa0_o_sum), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(cskip2_inst_rca0_fa31_o_sum), .Y(sum[5]) );
INVX1 INVX1_14 ( .A(1'b0), .Y(_8_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_9_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_10_) );
NAND3X1 NAND3X1_5 ( .A(_8_), .B(_10_), .C(_9_), .Y(_11_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_5_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_6_) );
OAI21X1 OAI21X1_11 ( .A(_5_), .B(_6_), .C(1'b0), .Y(_7_) );
NAND2X1 NAND2X1_17 ( .A(_7_), .B(_11_), .Y(_1__0_) );
OAI21X1 OAI21X1_12 ( .A(_8_), .B(_5_), .C(_10_), .Y(_3__1_) );
INVX1 INVX1_15 ( .A(_3__3_), .Y(_15_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_16_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_17_) );
NAND3X1 NAND3X1_6 ( .A(_15_), .B(_17_), .C(_16_), .Y(_18_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_12_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_13_) );
OAI21X1 OAI21X1_13 ( .A(_12_), .B(_13_), .C(_3__3_), .Y(_14_) );
NAND2X1 NAND2X1_19 ( .A(_14_), .B(_18_), .Y(_1__3_) );
OAI21X1 OAI21X1_14 ( .A(_15_), .B(_12_), .C(_17_), .Y(_2_) );
INVX1 INVX1_16 ( .A(_3__1_), .Y(_22_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_23_) );
BUFX2 BUFX2_8 ( .A(cskip2_inst_rca0_fa0_o_sum), .Y(_1__4_) );
BUFX2 BUFX2_9 ( .A(cskip2_inst_rca0_fa31_o_sum), .Y(_1__5_) );
endmodule
