module csa_55bit (i_add_term1, i_add_term2, sum, cout);

output cout;
input [54:0] i_add_term1;
input [54:0] i_add_term2;
output [54:0] sum;

wire vdd = 1'b1;
wire gnd = 1'b0;

NAND2X1 NAND2X1_1 ( .A(_2_), .B(rca_inst_cout), .Y(_74_) );
OAI21X1 OAI21X1_1 ( .A(rca_inst_cout), .B(_73_), .C(_74_), .Y(w_cout_1_) );
INVX1 INVX1_1 ( .A(_3__0_), .Y(_75_) );
NAND2X1 NAND2X1_2 ( .A(_4__0_), .B(rca_inst_cout), .Y(_76_) );
OAI21X1 OAI21X1_2 ( .A(rca_inst_cout), .B(_75_), .C(_76_), .Y(_0__4_) );
INVX1 INVX1_2 ( .A(_3__1_), .Y(_77_) );
NAND2X1 NAND2X1_3 ( .A(rca_inst_cout), .B(_4__1_), .Y(_78_) );
OAI21X1 OAI21X1_3 ( .A(rca_inst_cout), .B(_77_), .C(_78_), .Y(_0__5_) );
INVX1 INVX1_3 ( .A(_3__2_), .Y(_79_) );
NAND2X1 NAND2X1_4 ( .A(rca_inst_cout), .B(_4__2_), .Y(_80_) );
OAI21X1 OAI21X1_4 ( .A(rca_inst_cout), .B(_79_), .C(_80_), .Y(_0__6_) );
INVX1 INVX1_4 ( .A(_3__3_), .Y(_81_) );
NAND2X1 NAND2X1_5 ( .A(rca_inst_cout), .B(_4__3_), .Y(_82_) );
OAI21X1 OAI21X1_5 ( .A(rca_inst_cout), .B(_81_), .C(_82_), .Y(_0__7_) );
INVX1 INVX1_5 ( .A(gnd), .Y(_86_) );
OR2X2 OR2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_87_) );
NAND2X1 NAND2X1_6 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_88_) );
NAND3X1 NAND3X1_1 ( .A(_86_), .B(_88_), .C(_87_), .Y(_89_) );
NOR2X1 NOR2X1_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_83_) );
AND2X2 AND2X2_1 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_84_) );
OAI21X1 OAI21X1_6 ( .A(_83_), .B(_84_), .C(gnd), .Y(_85_) );
NAND2X1 NAND2X1_7 ( .A(_85_), .B(_89_), .Y(_3__0_) );
OAI21X1 OAI21X1_7 ( .A(_86_), .B(_83_), .C(_88_), .Y(_5__1_) );
INVX1 INVX1_6 ( .A(_5__3_), .Y(_93_) );
OR2X2 OR2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_94_) );
NAND2X1 NAND2X1_8 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_95_) );
NAND3X1 NAND3X1_2 ( .A(_93_), .B(_95_), .C(_94_), .Y(_96_) );
NOR2X1 NOR2X1_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_90_) );
AND2X2 AND2X2_2 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_91_) );
OAI21X1 OAI21X1_8 ( .A(_90_), .B(_91_), .C(_5__3_), .Y(_92_) );
NAND2X1 NAND2X1_9 ( .A(_92_), .B(_96_), .Y(_3__3_) );
OAI21X1 OAI21X1_9 ( .A(_93_), .B(_90_), .C(_95_), .Y(_1_) );
INVX1 INVX1_7 ( .A(_5__1_), .Y(_100_) );
OR2X2 OR2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_101_) );
NAND2X1 NAND2X1_10 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_102_) );
NAND3X1 NAND3X1_3 ( .A(_100_), .B(_102_), .C(_101_), .Y(_103_) );
NOR2X1 NOR2X1_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_97_) );
AND2X2 AND2X2_3 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_98_) );
OAI21X1 OAI21X1_10 ( .A(_97_), .B(_98_), .C(_5__1_), .Y(_99_) );
NAND2X1 NAND2X1_11 ( .A(_99_), .B(_103_), .Y(_3__1_) );
OAI21X1 OAI21X1_11 ( .A(_100_), .B(_97_), .C(_102_), .Y(_5__2_) );
INVX1 INVX1_8 ( .A(_5__2_), .Y(_107_) );
OR2X2 OR2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_108_) );
NAND2X1 NAND2X1_12 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_109_) );
NAND3X1 NAND3X1_4 ( .A(_107_), .B(_109_), .C(_108_), .Y(_110_) );
NOR2X1 NOR2X1_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_104_) );
AND2X2 AND2X2_4 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_105_) );
OAI21X1 OAI21X1_12 ( .A(_104_), .B(_105_), .C(_5__2_), .Y(_106_) );
NAND2X1 NAND2X1_13 ( .A(_106_), .B(_110_), .Y(_3__2_) );
OAI21X1 OAI21X1_13 ( .A(_107_), .B(_104_), .C(_109_), .Y(_5__3_) );
INVX1 INVX1_9 ( .A(vdd), .Y(_114_) );
OR2X2 OR2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_115_) );
NAND2X1 NAND2X1_14 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_116_) );
NAND3X1 NAND3X1_5 ( .A(_114_), .B(_116_), .C(_115_), .Y(_117_) );
NOR2X1 NOR2X1_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_111_) );
AND2X2 AND2X2_5 ( .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_112_) );
OAI21X1 OAI21X1_14 ( .A(_111_), .B(_112_), .C(vdd), .Y(_113_) );
NAND2X1 NAND2X1_15 ( .A(_113_), .B(_117_), .Y(_4__0_) );
OAI21X1 OAI21X1_15 ( .A(_114_), .B(_111_), .C(_116_), .Y(_6__1_) );
INVX1 INVX1_10 ( .A(_6__3_), .Y(_121_) );
OR2X2 OR2X2_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_122_) );
NAND2X1 NAND2X1_16 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_123_) );
NAND3X1 NAND3X1_6 ( .A(_121_), .B(_123_), .C(_122_), .Y(_124_) );
NOR2X1 NOR2X1_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_118_) );
AND2X2 AND2X2_6 ( .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_119_) );
OAI21X1 OAI21X1_16 ( .A(_118_), .B(_119_), .C(_6__3_), .Y(_120_) );
NAND2X1 NAND2X1_17 ( .A(_120_), .B(_124_), .Y(_4__3_) );
OAI21X1 OAI21X1_17 ( .A(_121_), .B(_118_), .C(_123_), .Y(_2_) );
INVX1 INVX1_11 ( .A(_6__1_), .Y(_128_) );
OR2X2 OR2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_129_) );
NAND2X1 NAND2X1_18 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_130_) );
NAND3X1 NAND3X1_7 ( .A(_128_), .B(_130_), .C(_129_), .Y(_131_) );
NOR2X1 NOR2X1_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_125_) );
AND2X2 AND2X2_7 ( .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_126_) );
OAI21X1 OAI21X1_18 ( .A(_125_), .B(_126_), .C(_6__1_), .Y(_127_) );
NAND2X1 NAND2X1_19 ( .A(_127_), .B(_131_), .Y(_4__1_) );
OAI21X1 OAI21X1_19 ( .A(_128_), .B(_125_), .C(_130_), .Y(_6__2_) );
INVX1 INVX1_12 ( .A(_6__2_), .Y(_135_) );
OR2X2 OR2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_136_) );
NAND2X1 NAND2X1_20 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_137_) );
NAND3X1 NAND3X1_8 ( .A(_135_), .B(_137_), .C(_136_), .Y(_138_) );
NOR2X1 NOR2X1_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_132_) );
AND2X2 AND2X2_8 ( .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_133_) );
OAI21X1 OAI21X1_20 ( .A(_132_), .B(_133_), .C(_6__2_), .Y(_134_) );
NAND2X1 NAND2X1_21 ( .A(_134_), .B(_138_), .Y(_4__2_) );
OAI21X1 OAI21X1_21 ( .A(_135_), .B(_132_), .C(_137_), .Y(_6__3_) );
INVX1 INVX1_13 ( .A(_7_), .Y(_139_) );
NAND2X1 NAND2X1_22 ( .A(_8_), .B(w_cout_1_), .Y(_140_) );
OAI21X1 OAI21X1_22 ( .A(w_cout_1_), .B(_139_), .C(_140_), .Y(w_cout_2_) );
INVX1 INVX1_14 ( .A(_9__0_), .Y(_141_) );
NAND2X1 NAND2X1_23 ( .A(_10__0_), .B(w_cout_1_), .Y(_142_) );
OAI21X1 OAI21X1_23 ( .A(w_cout_1_), .B(_141_), .C(_142_), .Y(_0__8_) );
INVX1 INVX1_15 ( .A(_9__1_), .Y(_143_) );
NAND2X1 NAND2X1_24 ( .A(w_cout_1_), .B(_10__1_), .Y(_144_) );
OAI21X1 OAI21X1_24 ( .A(w_cout_1_), .B(_143_), .C(_144_), .Y(_0__9_) );
INVX1 INVX1_16 ( .A(_9__2_), .Y(_145_) );
NAND2X1 NAND2X1_25 ( .A(w_cout_1_), .B(_10__2_), .Y(_146_) );
OAI21X1 OAI21X1_25 ( .A(w_cout_1_), .B(_145_), .C(_146_), .Y(_0__10_) );
INVX1 INVX1_17 ( .A(_9__3_), .Y(_147_) );
NAND2X1 NAND2X1_26 ( .A(w_cout_1_), .B(_10__3_), .Y(_148_) );
OAI21X1 OAI21X1_26 ( .A(w_cout_1_), .B(_147_), .C(_148_), .Y(_0__11_) );
INVX1 INVX1_18 ( .A(gnd), .Y(_152_) );
OR2X2 OR2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_153_) );
NAND2X1 NAND2X1_27 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_154_) );
NAND3X1 NAND3X1_9 ( .A(_152_), .B(_154_), .C(_153_), .Y(_155_) );
NOR2X1 NOR2X1_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_149_) );
AND2X2 AND2X2_9 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_150_) );
OAI21X1 OAI21X1_27 ( .A(_149_), .B(_150_), .C(gnd), .Y(_151_) );
NAND2X1 NAND2X1_28 ( .A(_151_), .B(_155_), .Y(_9__0_) );
OAI21X1 OAI21X1_28 ( .A(_152_), .B(_149_), .C(_154_), .Y(_11__1_) );
INVX1 INVX1_19 ( .A(_11__3_), .Y(_159_) );
OR2X2 OR2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_160_) );
NAND2X1 NAND2X1_29 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_161_) );
NAND3X1 NAND3X1_10 ( .A(_159_), .B(_161_), .C(_160_), .Y(_162_) );
NOR2X1 NOR2X1_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_156_) );
AND2X2 AND2X2_10 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_157_) );
OAI21X1 OAI21X1_29 ( .A(_156_), .B(_157_), .C(_11__3_), .Y(_158_) );
NAND2X1 NAND2X1_30 ( .A(_158_), .B(_162_), .Y(_9__3_) );
OAI21X1 OAI21X1_30 ( .A(_159_), .B(_156_), .C(_161_), .Y(_7_) );
INVX1 INVX1_20 ( .A(_11__1_), .Y(_166_) );
OR2X2 OR2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_167_) );
NAND2X1 NAND2X1_31 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_168_) );
NAND3X1 NAND3X1_11 ( .A(_166_), .B(_168_), .C(_167_), .Y(_169_) );
NOR2X1 NOR2X1_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_163_) );
AND2X2 AND2X2_11 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_164_) );
OAI21X1 OAI21X1_31 ( .A(_163_), .B(_164_), .C(_11__1_), .Y(_165_) );
NAND2X1 NAND2X1_32 ( .A(_165_), .B(_169_), .Y(_9__1_) );
OAI21X1 OAI21X1_32 ( .A(_166_), .B(_163_), .C(_168_), .Y(_11__2_) );
INVX1 INVX1_21 ( .A(_11__2_), .Y(_173_) );
OR2X2 OR2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_174_) );
NAND2X1 NAND2X1_33 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_175_) );
NAND3X1 NAND3X1_12 ( .A(_173_), .B(_175_), .C(_174_), .Y(_176_) );
NOR2X1 NOR2X1_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_170_) );
AND2X2 AND2X2_12 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_171_) );
OAI21X1 OAI21X1_33 ( .A(_170_), .B(_171_), .C(_11__2_), .Y(_172_) );
NAND2X1 NAND2X1_34 ( .A(_172_), .B(_176_), .Y(_9__2_) );
OAI21X1 OAI21X1_34 ( .A(_173_), .B(_170_), .C(_175_), .Y(_11__3_) );
INVX1 INVX1_22 ( .A(vdd), .Y(_180_) );
OR2X2 OR2X2_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_181_) );
NAND2X1 NAND2X1_35 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_182_) );
NAND3X1 NAND3X1_13 ( .A(_180_), .B(_182_), .C(_181_), .Y(_183_) );
NOR2X1 NOR2X1_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_177_) );
AND2X2 AND2X2_13 ( .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_178_) );
OAI21X1 OAI21X1_35 ( .A(_177_), .B(_178_), .C(vdd), .Y(_179_) );
NAND2X1 NAND2X1_36 ( .A(_179_), .B(_183_), .Y(_10__0_) );
OAI21X1 OAI21X1_36 ( .A(_180_), .B(_177_), .C(_182_), .Y(_12__1_) );
INVX1 INVX1_23 ( .A(_12__3_), .Y(_187_) );
OR2X2 OR2X2_14 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_188_) );
NAND2X1 NAND2X1_37 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_189_) );
NAND3X1 NAND3X1_14 ( .A(_187_), .B(_189_), .C(_188_), .Y(_190_) );
NOR2X1 NOR2X1_14 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_184_) );
AND2X2 AND2X2_14 ( .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_185_) );
OAI21X1 OAI21X1_37 ( .A(_184_), .B(_185_), .C(_12__3_), .Y(_186_) );
NAND2X1 NAND2X1_38 ( .A(_186_), .B(_190_), .Y(_10__3_) );
OAI21X1 OAI21X1_38 ( .A(_187_), .B(_184_), .C(_189_), .Y(_8_) );
INVX1 INVX1_24 ( .A(_12__1_), .Y(_194_) );
OR2X2 OR2X2_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_195_) );
NAND2X1 NAND2X1_39 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_196_) );
NAND3X1 NAND3X1_15 ( .A(_194_), .B(_196_), .C(_195_), .Y(_197_) );
NOR2X1 NOR2X1_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_191_) );
AND2X2 AND2X2_15 ( .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_192_) );
OAI21X1 OAI21X1_39 ( .A(_191_), .B(_192_), .C(_12__1_), .Y(_193_) );
NAND2X1 NAND2X1_40 ( .A(_193_), .B(_197_), .Y(_10__1_) );
OAI21X1 OAI21X1_40 ( .A(_194_), .B(_191_), .C(_196_), .Y(_12__2_) );
INVX1 INVX1_25 ( .A(_12__2_), .Y(_201_) );
OR2X2 OR2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_202_) );
NAND2X1 NAND2X1_41 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_203_) );
NAND3X1 NAND3X1_16 ( .A(_201_), .B(_203_), .C(_202_), .Y(_204_) );
NOR2X1 NOR2X1_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_198_) );
AND2X2 AND2X2_16 ( .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_199_) );
OAI21X1 OAI21X1_41 ( .A(_198_), .B(_199_), .C(_12__2_), .Y(_200_) );
NAND2X1 NAND2X1_42 ( .A(_200_), .B(_204_), .Y(_10__2_) );
OAI21X1 OAI21X1_42 ( .A(_201_), .B(_198_), .C(_203_), .Y(_12__3_) );
INVX1 INVX1_26 ( .A(_13_), .Y(_205_) );
NAND2X1 NAND2X1_43 ( .A(_14_), .B(w_cout_2_), .Y(_206_) );
OAI21X1 OAI21X1_43 ( .A(w_cout_2_), .B(_205_), .C(_206_), .Y(w_cout_3_) );
INVX1 INVX1_27 ( .A(_15__0_), .Y(_207_) );
NAND2X1 NAND2X1_44 ( .A(_16__0_), .B(w_cout_2_), .Y(_208_) );
OAI21X1 OAI21X1_44 ( .A(w_cout_2_), .B(_207_), .C(_208_), .Y(_0__12_) );
INVX1 INVX1_28 ( .A(_15__1_), .Y(_209_) );
NAND2X1 NAND2X1_45 ( .A(w_cout_2_), .B(_16__1_), .Y(_210_) );
OAI21X1 OAI21X1_45 ( .A(w_cout_2_), .B(_209_), .C(_210_), .Y(_0__13_) );
INVX1 INVX1_29 ( .A(_15__2_), .Y(_211_) );
NAND2X1 NAND2X1_46 ( .A(w_cout_2_), .B(_16__2_), .Y(_212_) );
OAI21X1 OAI21X1_46 ( .A(w_cout_2_), .B(_211_), .C(_212_), .Y(_0__14_) );
INVX1 INVX1_30 ( .A(_15__3_), .Y(_213_) );
NAND2X1 NAND2X1_47 ( .A(w_cout_2_), .B(_16__3_), .Y(_214_) );
OAI21X1 OAI21X1_47 ( .A(w_cout_2_), .B(_213_), .C(_214_), .Y(_0__15_) );
INVX1 INVX1_31 ( .A(gnd), .Y(_218_) );
OR2X2 OR2X2_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_219_) );
NAND2X1 NAND2X1_48 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_220_) );
NAND3X1 NAND3X1_17 ( .A(_218_), .B(_220_), .C(_219_), .Y(_221_) );
NOR2X1 NOR2X1_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_215_) );
AND2X2 AND2X2_17 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_216_) );
OAI21X1 OAI21X1_48 ( .A(_215_), .B(_216_), .C(gnd), .Y(_217_) );
NAND2X1 NAND2X1_49 ( .A(_217_), .B(_221_), .Y(_15__0_) );
OAI21X1 OAI21X1_49 ( .A(_218_), .B(_215_), .C(_220_), .Y(_17__1_) );
INVX1 INVX1_32 ( .A(_17__3_), .Y(_225_) );
OR2X2 OR2X2_18 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_226_) );
NAND2X1 NAND2X1_50 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_227_) );
NAND3X1 NAND3X1_18 ( .A(_225_), .B(_227_), .C(_226_), .Y(_228_) );
NOR2X1 NOR2X1_18 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_222_) );
AND2X2 AND2X2_18 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_223_) );
OAI21X1 OAI21X1_50 ( .A(_222_), .B(_223_), .C(_17__3_), .Y(_224_) );
NAND2X1 NAND2X1_51 ( .A(_224_), .B(_228_), .Y(_15__3_) );
OAI21X1 OAI21X1_51 ( .A(_225_), .B(_222_), .C(_227_), .Y(_13_) );
INVX1 INVX1_33 ( .A(_17__1_), .Y(_232_) );
OR2X2 OR2X2_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_233_) );
NAND2X1 NAND2X1_52 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_234_) );
NAND3X1 NAND3X1_19 ( .A(_232_), .B(_234_), .C(_233_), .Y(_235_) );
NOR2X1 NOR2X1_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_229_) );
AND2X2 AND2X2_19 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_230_) );
OAI21X1 OAI21X1_52 ( .A(_229_), .B(_230_), .C(_17__1_), .Y(_231_) );
NAND2X1 NAND2X1_53 ( .A(_231_), .B(_235_), .Y(_15__1_) );
OAI21X1 OAI21X1_53 ( .A(_232_), .B(_229_), .C(_234_), .Y(_17__2_) );
INVX1 INVX1_34 ( .A(_17__2_), .Y(_239_) );
OR2X2 OR2X2_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_240_) );
NAND2X1 NAND2X1_54 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_241_) );
NAND3X1 NAND3X1_20 ( .A(_239_), .B(_241_), .C(_240_), .Y(_242_) );
NOR2X1 NOR2X1_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_236_) );
AND2X2 AND2X2_20 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_237_) );
OAI21X1 OAI21X1_54 ( .A(_236_), .B(_237_), .C(_17__2_), .Y(_238_) );
NAND2X1 NAND2X1_55 ( .A(_238_), .B(_242_), .Y(_15__2_) );
OAI21X1 OAI21X1_55 ( .A(_239_), .B(_236_), .C(_241_), .Y(_17__3_) );
INVX1 INVX1_35 ( .A(vdd), .Y(_246_) );
OR2X2 OR2X2_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_247_) );
NAND2X1 NAND2X1_56 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_248_) );
NAND3X1 NAND3X1_21 ( .A(_246_), .B(_248_), .C(_247_), .Y(_249_) );
NOR2X1 NOR2X1_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_243_) );
AND2X2 AND2X2_21 ( .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_244_) );
OAI21X1 OAI21X1_56 ( .A(_243_), .B(_244_), .C(vdd), .Y(_245_) );
NAND2X1 NAND2X1_57 ( .A(_245_), .B(_249_), .Y(_16__0_) );
OAI21X1 OAI21X1_57 ( .A(_246_), .B(_243_), .C(_248_), .Y(_18__1_) );
INVX1 INVX1_36 ( .A(_18__3_), .Y(_253_) );
OR2X2 OR2X2_22 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_254_) );
NAND2X1 NAND2X1_58 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_255_) );
NAND3X1 NAND3X1_22 ( .A(_253_), .B(_255_), .C(_254_), .Y(_256_) );
NOR2X1 NOR2X1_22 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_250_) );
AND2X2 AND2X2_22 ( .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_251_) );
OAI21X1 OAI21X1_58 ( .A(_250_), .B(_251_), .C(_18__3_), .Y(_252_) );
NAND2X1 NAND2X1_59 ( .A(_252_), .B(_256_), .Y(_16__3_) );
OAI21X1 OAI21X1_59 ( .A(_253_), .B(_250_), .C(_255_), .Y(_14_) );
INVX1 INVX1_37 ( .A(_18__1_), .Y(_260_) );
OR2X2 OR2X2_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_261_) );
NAND2X1 NAND2X1_60 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_262_) );
NAND3X1 NAND3X1_23 ( .A(_260_), .B(_262_), .C(_261_), .Y(_263_) );
NOR2X1 NOR2X1_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_257_) );
AND2X2 AND2X2_23 ( .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_258_) );
OAI21X1 OAI21X1_60 ( .A(_257_), .B(_258_), .C(_18__1_), .Y(_259_) );
NAND2X1 NAND2X1_61 ( .A(_259_), .B(_263_), .Y(_16__1_) );
OAI21X1 OAI21X1_61 ( .A(_260_), .B(_257_), .C(_262_), .Y(_18__2_) );
INVX1 INVX1_38 ( .A(_18__2_), .Y(_267_) );
OR2X2 OR2X2_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_268_) );
NAND2X1 NAND2X1_62 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_269_) );
NAND3X1 NAND3X1_24 ( .A(_267_), .B(_269_), .C(_268_), .Y(_270_) );
NOR2X1 NOR2X1_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_264_) );
AND2X2 AND2X2_24 ( .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_265_) );
OAI21X1 OAI21X1_62 ( .A(_264_), .B(_265_), .C(_18__2_), .Y(_266_) );
NAND2X1 NAND2X1_63 ( .A(_266_), .B(_270_), .Y(_16__2_) );
OAI21X1 OAI21X1_63 ( .A(_267_), .B(_264_), .C(_269_), .Y(_18__3_) );
INVX1 INVX1_39 ( .A(_19_), .Y(_271_) );
NAND2X1 NAND2X1_64 ( .A(_20_), .B(w_cout_3_), .Y(_272_) );
OAI21X1 OAI21X1_64 ( .A(w_cout_3_), .B(_271_), .C(_272_), .Y(w_cout_4_) );
INVX1 INVX1_40 ( .A(_21__0_), .Y(_273_) );
NAND2X1 NAND2X1_65 ( .A(_22__0_), .B(w_cout_3_), .Y(_274_) );
OAI21X1 OAI21X1_65 ( .A(w_cout_3_), .B(_273_), .C(_274_), .Y(_0__16_) );
INVX1 INVX1_41 ( .A(_21__1_), .Y(_275_) );
NAND2X1 NAND2X1_66 ( .A(w_cout_3_), .B(_22__1_), .Y(_276_) );
OAI21X1 OAI21X1_66 ( .A(w_cout_3_), .B(_275_), .C(_276_), .Y(_0__17_) );
INVX1 INVX1_42 ( .A(_21__2_), .Y(_277_) );
NAND2X1 NAND2X1_67 ( .A(w_cout_3_), .B(_22__2_), .Y(_278_) );
OAI21X1 OAI21X1_67 ( .A(w_cout_3_), .B(_277_), .C(_278_), .Y(_0__18_) );
INVX1 INVX1_43 ( .A(_21__3_), .Y(_279_) );
NAND2X1 NAND2X1_68 ( .A(w_cout_3_), .B(_22__3_), .Y(_280_) );
OAI21X1 OAI21X1_68 ( .A(w_cout_3_), .B(_279_), .C(_280_), .Y(_0__19_) );
INVX1 INVX1_44 ( .A(gnd), .Y(_284_) );
OR2X2 OR2X2_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_285_) );
NAND2X1 NAND2X1_69 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_286_) );
NAND3X1 NAND3X1_25 ( .A(_284_), .B(_286_), .C(_285_), .Y(_287_) );
NOR2X1 NOR2X1_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_281_) );
AND2X2 AND2X2_25 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_282_) );
OAI21X1 OAI21X1_69 ( .A(_281_), .B(_282_), .C(gnd), .Y(_283_) );
NAND2X1 NAND2X1_70 ( .A(_283_), .B(_287_), .Y(_21__0_) );
OAI21X1 OAI21X1_70 ( .A(_284_), .B(_281_), .C(_286_), .Y(_23__1_) );
INVX1 INVX1_45 ( .A(_23__3_), .Y(_291_) );
OR2X2 OR2X2_26 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_292_) );
NAND2X1 NAND2X1_71 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_293_) );
NAND3X1 NAND3X1_26 ( .A(_291_), .B(_293_), .C(_292_), .Y(_294_) );
NOR2X1 NOR2X1_26 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_288_) );
AND2X2 AND2X2_26 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_289_) );
OAI21X1 OAI21X1_71 ( .A(_288_), .B(_289_), .C(_23__3_), .Y(_290_) );
NAND2X1 NAND2X1_72 ( .A(_290_), .B(_294_), .Y(_21__3_) );
OAI21X1 OAI21X1_72 ( .A(_291_), .B(_288_), .C(_293_), .Y(_19_) );
INVX1 INVX1_46 ( .A(_23__1_), .Y(_298_) );
OR2X2 OR2X2_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_299_) );
NAND2X1 NAND2X1_73 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_300_) );
NAND3X1 NAND3X1_27 ( .A(_298_), .B(_300_), .C(_299_), .Y(_301_) );
NOR2X1 NOR2X1_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_295_) );
AND2X2 AND2X2_27 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_296_) );
OAI21X1 OAI21X1_73 ( .A(_295_), .B(_296_), .C(_23__1_), .Y(_297_) );
NAND2X1 NAND2X1_74 ( .A(_297_), .B(_301_), .Y(_21__1_) );
OAI21X1 OAI21X1_74 ( .A(_298_), .B(_295_), .C(_300_), .Y(_23__2_) );
INVX1 INVX1_47 ( .A(_23__2_), .Y(_305_) );
OR2X2 OR2X2_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_306_) );
NAND2X1 NAND2X1_75 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_307_) );
NAND3X1 NAND3X1_28 ( .A(_305_), .B(_307_), .C(_306_), .Y(_308_) );
NOR2X1 NOR2X1_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_302_) );
AND2X2 AND2X2_28 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_303_) );
OAI21X1 OAI21X1_75 ( .A(_302_), .B(_303_), .C(_23__2_), .Y(_304_) );
NAND2X1 NAND2X1_76 ( .A(_304_), .B(_308_), .Y(_21__2_) );
OAI21X1 OAI21X1_76 ( .A(_305_), .B(_302_), .C(_307_), .Y(_23__3_) );
INVX1 INVX1_48 ( .A(vdd), .Y(_312_) );
OR2X2 OR2X2_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_313_) );
NAND2X1 NAND2X1_77 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_314_) );
NAND3X1 NAND3X1_29 ( .A(_312_), .B(_314_), .C(_313_), .Y(_315_) );
NOR2X1 NOR2X1_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_309_) );
AND2X2 AND2X2_29 ( .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_310_) );
OAI21X1 OAI21X1_77 ( .A(_309_), .B(_310_), .C(vdd), .Y(_311_) );
NAND2X1 NAND2X1_78 ( .A(_311_), .B(_315_), .Y(_22__0_) );
OAI21X1 OAI21X1_78 ( .A(_312_), .B(_309_), .C(_314_), .Y(_24__1_) );
INVX1 INVX1_49 ( .A(_24__3_), .Y(_319_) );
OR2X2 OR2X2_30 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_320_) );
NAND2X1 NAND2X1_79 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_321_) );
NAND3X1 NAND3X1_30 ( .A(_319_), .B(_321_), .C(_320_), .Y(_322_) );
NOR2X1 NOR2X1_30 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_316_) );
AND2X2 AND2X2_30 ( .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_317_) );
OAI21X1 OAI21X1_79 ( .A(_316_), .B(_317_), .C(_24__3_), .Y(_318_) );
NAND2X1 NAND2X1_80 ( .A(_318_), .B(_322_), .Y(_22__3_) );
OAI21X1 OAI21X1_80 ( .A(_319_), .B(_316_), .C(_321_), .Y(_20_) );
INVX1 INVX1_50 ( .A(_24__1_), .Y(_326_) );
OR2X2 OR2X2_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_327_) );
NAND2X1 NAND2X1_81 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_328_) );
NAND3X1 NAND3X1_31 ( .A(_326_), .B(_328_), .C(_327_), .Y(_329_) );
NOR2X1 NOR2X1_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_323_) );
AND2X2 AND2X2_31 ( .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_324_) );
OAI21X1 OAI21X1_81 ( .A(_323_), .B(_324_), .C(_24__1_), .Y(_325_) );
NAND2X1 NAND2X1_82 ( .A(_325_), .B(_329_), .Y(_22__1_) );
OAI21X1 OAI21X1_82 ( .A(_326_), .B(_323_), .C(_328_), .Y(_24__2_) );
INVX1 INVX1_51 ( .A(_24__2_), .Y(_333_) );
OR2X2 OR2X2_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_334_) );
NAND2X1 NAND2X1_83 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_335_) );
NAND3X1 NAND3X1_32 ( .A(_333_), .B(_335_), .C(_334_), .Y(_336_) );
NOR2X1 NOR2X1_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_330_) );
AND2X2 AND2X2_32 ( .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_331_) );
OAI21X1 OAI21X1_83 ( .A(_330_), .B(_331_), .C(_24__2_), .Y(_332_) );
NAND2X1 NAND2X1_84 ( .A(_332_), .B(_336_), .Y(_22__2_) );
OAI21X1 OAI21X1_84 ( .A(_333_), .B(_330_), .C(_335_), .Y(_24__3_) );
INVX1 INVX1_52 ( .A(_25_), .Y(_337_) );
NAND2X1 NAND2X1_85 ( .A(_26_), .B(w_cout_4_), .Y(_338_) );
OAI21X1 OAI21X1_85 ( .A(w_cout_4_), .B(_337_), .C(_338_), .Y(w_cout_5_) );
INVX1 INVX1_53 ( .A(_27__0_), .Y(_339_) );
NAND2X1 NAND2X1_86 ( .A(_28__0_), .B(w_cout_4_), .Y(_340_) );
OAI21X1 OAI21X1_86 ( .A(w_cout_4_), .B(_339_), .C(_340_), .Y(_0__20_) );
INVX1 INVX1_54 ( .A(_27__1_), .Y(_341_) );
NAND2X1 NAND2X1_87 ( .A(w_cout_4_), .B(_28__1_), .Y(_342_) );
OAI21X1 OAI21X1_87 ( .A(w_cout_4_), .B(_341_), .C(_342_), .Y(_0__21_) );
INVX1 INVX1_55 ( .A(_27__2_), .Y(_343_) );
NAND2X1 NAND2X1_88 ( .A(w_cout_4_), .B(_28__2_), .Y(_344_) );
OAI21X1 OAI21X1_88 ( .A(w_cout_4_), .B(_343_), .C(_344_), .Y(_0__22_) );
INVX1 INVX1_56 ( .A(_27__3_), .Y(_345_) );
NAND2X1 NAND2X1_89 ( .A(w_cout_4_), .B(_28__3_), .Y(_346_) );
OAI21X1 OAI21X1_89 ( .A(w_cout_4_), .B(_345_), .C(_346_), .Y(_0__23_) );
INVX1 INVX1_57 ( .A(gnd), .Y(_350_) );
OR2X2 OR2X2_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_351_) );
NAND2X1 NAND2X1_90 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_352_) );
NAND3X1 NAND3X1_33 ( .A(_350_), .B(_352_), .C(_351_), .Y(_353_) );
NOR2X1 NOR2X1_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_347_) );
AND2X2 AND2X2_33 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_348_) );
OAI21X1 OAI21X1_90 ( .A(_347_), .B(_348_), .C(gnd), .Y(_349_) );
NAND2X1 NAND2X1_91 ( .A(_349_), .B(_353_), .Y(_27__0_) );
OAI21X1 OAI21X1_91 ( .A(_350_), .B(_347_), .C(_352_), .Y(_29__1_) );
INVX1 INVX1_58 ( .A(_29__3_), .Y(_357_) );
OR2X2 OR2X2_34 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_358_) );
NAND2X1 NAND2X1_92 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_359_) );
NAND3X1 NAND3X1_34 ( .A(_357_), .B(_359_), .C(_358_), .Y(_360_) );
NOR2X1 NOR2X1_34 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_354_) );
AND2X2 AND2X2_34 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_355_) );
OAI21X1 OAI21X1_92 ( .A(_354_), .B(_355_), .C(_29__3_), .Y(_356_) );
NAND2X1 NAND2X1_93 ( .A(_356_), .B(_360_), .Y(_27__3_) );
OAI21X1 OAI21X1_93 ( .A(_357_), .B(_354_), .C(_359_), .Y(_25_) );
INVX1 INVX1_59 ( .A(_29__1_), .Y(_364_) );
OR2X2 OR2X2_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_365_) );
NAND2X1 NAND2X1_94 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_366_) );
NAND3X1 NAND3X1_35 ( .A(_364_), .B(_366_), .C(_365_), .Y(_367_) );
NOR2X1 NOR2X1_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_361_) );
AND2X2 AND2X2_35 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_362_) );
OAI21X1 OAI21X1_94 ( .A(_361_), .B(_362_), .C(_29__1_), .Y(_363_) );
NAND2X1 NAND2X1_95 ( .A(_363_), .B(_367_), .Y(_27__1_) );
OAI21X1 OAI21X1_95 ( .A(_364_), .B(_361_), .C(_366_), .Y(_29__2_) );
INVX1 INVX1_60 ( .A(_29__2_), .Y(_371_) );
OR2X2 OR2X2_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_372_) );
NAND2X1 NAND2X1_96 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_373_) );
NAND3X1 NAND3X1_36 ( .A(_371_), .B(_373_), .C(_372_), .Y(_374_) );
NOR2X1 NOR2X1_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_368_) );
AND2X2 AND2X2_36 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_369_) );
OAI21X1 OAI21X1_96 ( .A(_368_), .B(_369_), .C(_29__2_), .Y(_370_) );
NAND2X1 NAND2X1_97 ( .A(_370_), .B(_374_), .Y(_27__2_) );
OAI21X1 OAI21X1_97 ( .A(_371_), .B(_368_), .C(_373_), .Y(_29__3_) );
INVX1 INVX1_61 ( .A(vdd), .Y(_378_) );
OR2X2 OR2X2_37 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_379_) );
NAND2X1 NAND2X1_98 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_380_) );
NAND3X1 NAND3X1_37 ( .A(_378_), .B(_380_), .C(_379_), .Y(_381_) );
NOR2X1 NOR2X1_37 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_375_) );
AND2X2 AND2X2_37 ( .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_376_) );
OAI21X1 OAI21X1_98 ( .A(_375_), .B(_376_), .C(vdd), .Y(_377_) );
NAND2X1 NAND2X1_99 ( .A(_377_), .B(_381_), .Y(_28__0_) );
OAI21X1 OAI21X1_99 ( .A(_378_), .B(_375_), .C(_380_), .Y(_30__1_) );
INVX1 INVX1_62 ( .A(_30__3_), .Y(_385_) );
OR2X2 OR2X2_38 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_386_) );
NAND2X1 NAND2X1_100 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_387_) );
NAND3X1 NAND3X1_38 ( .A(_385_), .B(_387_), .C(_386_), .Y(_388_) );
NOR2X1 NOR2X1_38 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_382_) );
AND2X2 AND2X2_38 ( .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_383_) );
OAI21X1 OAI21X1_100 ( .A(_382_), .B(_383_), .C(_30__3_), .Y(_384_) );
NAND2X1 NAND2X1_101 ( .A(_384_), .B(_388_), .Y(_28__3_) );
OAI21X1 OAI21X1_101 ( .A(_385_), .B(_382_), .C(_387_), .Y(_26_) );
INVX1 INVX1_63 ( .A(_30__1_), .Y(_392_) );
OR2X2 OR2X2_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_393_) );
NAND2X1 NAND2X1_102 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_394_) );
NAND3X1 NAND3X1_39 ( .A(_392_), .B(_394_), .C(_393_), .Y(_395_) );
NOR2X1 NOR2X1_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_389_) );
AND2X2 AND2X2_39 ( .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_390_) );
OAI21X1 OAI21X1_102 ( .A(_389_), .B(_390_), .C(_30__1_), .Y(_391_) );
NAND2X1 NAND2X1_103 ( .A(_391_), .B(_395_), .Y(_28__1_) );
OAI21X1 OAI21X1_103 ( .A(_392_), .B(_389_), .C(_394_), .Y(_30__2_) );
INVX1 INVX1_64 ( .A(_30__2_), .Y(_399_) );
OR2X2 OR2X2_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_400_) );
NAND2X1 NAND2X1_104 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_401_) );
NAND3X1 NAND3X1_40 ( .A(_399_), .B(_401_), .C(_400_), .Y(_402_) );
NOR2X1 NOR2X1_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_396_) );
AND2X2 AND2X2_40 ( .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_397_) );
OAI21X1 OAI21X1_104 ( .A(_396_), .B(_397_), .C(_30__2_), .Y(_398_) );
NAND2X1 NAND2X1_105 ( .A(_398_), .B(_402_), .Y(_28__2_) );
OAI21X1 OAI21X1_105 ( .A(_399_), .B(_396_), .C(_401_), .Y(_30__3_) );
INVX1 INVX1_65 ( .A(_31_), .Y(_403_) );
NAND2X1 NAND2X1_106 ( .A(_32_), .B(w_cout_5_), .Y(_404_) );
OAI21X1 OAI21X1_106 ( .A(w_cout_5_), .B(_403_), .C(_404_), .Y(w_cout_6_) );
INVX1 INVX1_66 ( .A(_33__0_), .Y(_405_) );
NAND2X1 NAND2X1_107 ( .A(_34__0_), .B(w_cout_5_), .Y(_406_) );
OAI21X1 OAI21X1_107 ( .A(w_cout_5_), .B(_405_), .C(_406_), .Y(_0__24_) );
INVX1 INVX1_67 ( .A(_33__1_), .Y(_407_) );
NAND2X1 NAND2X1_108 ( .A(w_cout_5_), .B(_34__1_), .Y(_408_) );
OAI21X1 OAI21X1_108 ( .A(w_cout_5_), .B(_407_), .C(_408_), .Y(_0__25_) );
INVX1 INVX1_68 ( .A(_33__2_), .Y(_409_) );
NAND2X1 NAND2X1_109 ( .A(w_cout_5_), .B(_34__2_), .Y(_410_) );
OAI21X1 OAI21X1_109 ( .A(w_cout_5_), .B(_409_), .C(_410_), .Y(_0__26_) );
INVX1 INVX1_69 ( .A(_33__3_), .Y(_411_) );
NAND2X1 NAND2X1_110 ( .A(w_cout_5_), .B(_34__3_), .Y(_412_) );
OAI21X1 OAI21X1_110 ( .A(w_cout_5_), .B(_411_), .C(_412_), .Y(_0__27_) );
INVX1 INVX1_70 ( .A(gnd), .Y(_416_) );
OR2X2 OR2X2_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_417_) );
NAND2X1 NAND2X1_111 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_418_) );
NAND3X1 NAND3X1_41 ( .A(_416_), .B(_418_), .C(_417_), .Y(_419_) );
NOR2X1 NOR2X1_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_413_) );
AND2X2 AND2X2_41 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_414_) );
OAI21X1 OAI21X1_111 ( .A(_413_), .B(_414_), .C(gnd), .Y(_415_) );
NAND2X1 NAND2X1_112 ( .A(_415_), .B(_419_), .Y(_33__0_) );
OAI21X1 OAI21X1_112 ( .A(_416_), .B(_413_), .C(_418_), .Y(_35__1_) );
INVX1 INVX1_71 ( .A(_35__3_), .Y(_423_) );
OR2X2 OR2X2_42 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_424_) );
NAND2X1 NAND2X1_113 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_425_) );
NAND3X1 NAND3X1_42 ( .A(_423_), .B(_425_), .C(_424_), .Y(_426_) );
NOR2X1 NOR2X1_42 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_420_) );
AND2X2 AND2X2_42 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_421_) );
OAI21X1 OAI21X1_113 ( .A(_420_), .B(_421_), .C(_35__3_), .Y(_422_) );
NAND2X1 NAND2X1_114 ( .A(_422_), .B(_426_), .Y(_33__3_) );
OAI21X1 OAI21X1_114 ( .A(_423_), .B(_420_), .C(_425_), .Y(_31_) );
INVX1 INVX1_72 ( .A(_35__1_), .Y(_430_) );
OR2X2 OR2X2_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_431_) );
NAND2X1 NAND2X1_115 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_432_) );
NAND3X1 NAND3X1_43 ( .A(_430_), .B(_432_), .C(_431_), .Y(_433_) );
NOR2X1 NOR2X1_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_427_) );
AND2X2 AND2X2_43 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_428_) );
OAI21X1 OAI21X1_115 ( .A(_427_), .B(_428_), .C(_35__1_), .Y(_429_) );
NAND2X1 NAND2X1_116 ( .A(_429_), .B(_433_), .Y(_33__1_) );
OAI21X1 OAI21X1_116 ( .A(_430_), .B(_427_), .C(_432_), .Y(_35__2_) );
INVX1 INVX1_73 ( .A(_35__2_), .Y(_437_) );
OR2X2 OR2X2_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_438_) );
NAND2X1 NAND2X1_117 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_439_) );
NAND3X1 NAND3X1_44 ( .A(_437_), .B(_439_), .C(_438_), .Y(_440_) );
NOR2X1 NOR2X1_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_434_) );
AND2X2 AND2X2_44 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_435_) );
OAI21X1 OAI21X1_117 ( .A(_434_), .B(_435_), .C(_35__2_), .Y(_436_) );
NAND2X1 NAND2X1_118 ( .A(_436_), .B(_440_), .Y(_33__2_) );
OAI21X1 OAI21X1_118 ( .A(_437_), .B(_434_), .C(_439_), .Y(_35__3_) );
INVX1 INVX1_74 ( .A(vdd), .Y(_444_) );
OR2X2 OR2X2_45 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_445_) );
NAND2X1 NAND2X1_119 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_446_) );
NAND3X1 NAND3X1_45 ( .A(_444_), .B(_446_), .C(_445_), .Y(_447_) );
NOR2X1 NOR2X1_45 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_441_) );
AND2X2 AND2X2_45 ( .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_442_) );
OAI21X1 OAI21X1_119 ( .A(_441_), .B(_442_), .C(vdd), .Y(_443_) );
NAND2X1 NAND2X1_120 ( .A(_443_), .B(_447_), .Y(_34__0_) );
OAI21X1 OAI21X1_120 ( .A(_444_), .B(_441_), .C(_446_), .Y(_36__1_) );
INVX1 INVX1_75 ( .A(_36__3_), .Y(_451_) );
OR2X2 OR2X2_46 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_452_) );
NAND2X1 NAND2X1_121 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_453_) );
NAND3X1 NAND3X1_46 ( .A(_451_), .B(_453_), .C(_452_), .Y(_454_) );
NOR2X1 NOR2X1_46 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_448_) );
AND2X2 AND2X2_46 ( .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_449_) );
OAI21X1 OAI21X1_121 ( .A(_448_), .B(_449_), .C(_36__3_), .Y(_450_) );
NAND2X1 NAND2X1_122 ( .A(_450_), .B(_454_), .Y(_34__3_) );
OAI21X1 OAI21X1_122 ( .A(_451_), .B(_448_), .C(_453_), .Y(_32_) );
INVX1 INVX1_76 ( .A(_36__1_), .Y(_458_) );
OR2X2 OR2X2_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_459_) );
NAND2X1 NAND2X1_123 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_460_) );
NAND3X1 NAND3X1_47 ( .A(_458_), .B(_460_), .C(_459_), .Y(_461_) );
NOR2X1 NOR2X1_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_455_) );
AND2X2 AND2X2_47 ( .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_456_) );
OAI21X1 OAI21X1_123 ( .A(_455_), .B(_456_), .C(_36__1_), .Y(_457_) );
NAND2X1 NAND2X1_124 ( .A(_457_), .B(_461_), .Y(_34__1_) );
OAI21X1 OAI21X1_124 ( .A(_458_), .B(_455_), .C(_460_), .Y(_36__2_) );
INVX1 INVX1_77 ( .A(_36__2_), .Y(_465_) );
OR2X2 OR2X2_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_466_) );
NAND2X1 NAND2X1_125 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_467_) );
NAND3X1 NAND3X1_48 ( .A(_465_), .B(_467_), .C(_466_), .Y(_468_) );
NOR2X1 NOR2X1_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_462_) );
AND2X2 AND2X2_48 ( .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_463_) );
OAI21X1 OAI21X1_125 ( .A(_462_), .B(_463_), .C(_36__2_), .Y(_464_) );
NAND2X1 NAND2X1_126 ( .A(_464_), .B(_468_), .Y(_34__2_) );
OAI21X1 OAI21X1_126 ( .A(_465_), .B(_462_), .C(_467_), .Y(_36__3_) );
INVX1 INVX1_78 ( .A(_37_), .Y(_469_) );
NAND2X1 NAND2X1_127 ( .A(_38_), .B(w_cout_6_), .Y(_470_) );
OAI21X1 OAI21X1_127 ( .A(w_cout_6_), .B(_469_), .C(_470_), .Y(w_cout_7_) );
INVX1 INVX1_79 ( .A(_39__0_), .Y(_471_) );
NAND2X1 NAND2X1_128 ( .A(_40__0_), .B(w_cout_6_), .Y(_472_) );
OAI21X1 OAI21X1_128 ( .A(w_cout_6_), .B(_471_), .C(_472_), .Y(_0__28_) );
INVX1 INVX1_80 ( .A(_39__1_), .Y(_473_) );
NAND2X1 NAND2X1_129 ( .A(w_cout_6_), .B(_40__1_), .Y(_474_) );
OAI21X1 OAI21X1_129 ( .A(w_cout_6_), .B(_473_), .C(_474_), .Y(_0__29_) );
INVX1 INVX1_81 ( .A(_39__2_), .Y(_475_) );
NAND2X1 NAND2X1_130 ( .A(w_cout_6_), .B(_40__2_), .Y(_476_) );
OAI21X1 OAI21X1_130 ( .A(w_cout_6_), .B(_475_), .C(_476_), .Y(_0__30_) );
INVX1 INVX1_82 ( .A(_39__3_), .Y(_477_) );
NAND2X1 NAND2X1_131 ( .A(w_cout_6_), .B(_40__3_), .Y(_478_) );
OAI21X1 OAI21X1_131 ( .A(w_cout_6_), .B(_477_), .C(_478_), .Y(_0__31_) );
INVX1 INVX1_83 ( .A(gnd), .Y(_482_) );
OR2X2 OR2X2_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_483_) );
NAND2X1 NAND2X1_132 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_484_) );
NAND3X1 NAND3X1_49 ( .A(_482_), .B(_484_), .C(_483_), .Y(_485_) );
NOR2X1 NOR2X1_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_479_) );
AND2X2 AND2X2_49 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_480_) );
OAI21X1 OAI21X1_132 ( .A(_479_), .B(_480_), .C(gnd), .Y(_481_) );
NAND2X1 NAND2X1_133 ( .A(_481_), .B(_485_), .Y(_39__0_) );
OAI21X1 OAI21X1_133 ( .A(_482_), .B(_479_), .C(_484_), .Y(_41__1_) );
INVX1 INVX1_84 ( .A(_41__3_), .Y(_489_) );
OR2X2 OR2X2_50 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_490_) );
NAND2X1 NAND2X1_134 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_491_) );
NAND3X1 NAND3X1_50 ( .A(_489_), .B(_491_), .C(_490_), .Y(_492_) );
NOR2X1 NOR2X1_50 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_486_) );
AND2X2 AND2X2_50 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_487_) );
OAI21X1 OAI21X1_134 ( .A(_486_), .B(_487_), .C(_41__3_), .Y(_488_) );
NAND2X1 NAND2X1_135 ( .A(_488_), .B(_492_), .Y(_39__3_) );
OAI21X1 OAI21X1_135 ( .A(_489_), .B(_486_), .C(_491_), .Y(_37_) );
INVX1 INVX1_85 ( .A(_41__1_), .Y(_496_) );
OR2X2 OR2X2_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_497_) );
NAND2X1 NAND2X1_136 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_498_) );
NAND3X1 NAND3X1_51 ( .A(_496_), .B(_498_), .C(_497_), .Y(_499_) );
NOR2X1 NOR2X1_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_493_) );
AND2X2 AND2X2_51 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_494_) );
OAI21X1 OAI21X1_136 ( .A(_493_), .B(_494_), .C(_41__1_), .Y(_495_) );
NAND2X1 NAND2X1_137 ( .A(_495_), .B(_499_), .Y(_39__1_) );
OAI21X1 OAI21X1_137 ( .A(_496_), .B(_493_), .C(_498_), .Y(_41__2_) );
INVX1 INVX1_86 ( .A(_41__2_), .Y(_503_) );
OR2X2 OR2X2_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_504_) );
NAND2X1 NAND2X1_138 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_505_) );
NAND3X1 NAND3X1_52 ( .A(_503_), .B(_505_), .C(_504_), .Y(_506_) );
NOR2X1 NOR2X1_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_500_) );
AND2X2 AND2X2_52 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_501_) );
OAI21X1 OAI21X1_138 ( .A(_500_), .B(_501_), .C(_41__2_), .Y(_502_) );
NAND2X1 NAND2X1_139 ( .A(_502_), .B(_506_), .Y(_39__2_) );
OAI21X1 OAI21X1_139 ( .A(_503_), .B(_500_), .C(_505_), .Y(_41__3_) );
INVX1 INVX1_87 ( .A(vdd), .Y(_510_) );
OR2X2 OR2X2_53 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_511_) );
NAND2X1 NAND2X1_140 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_512_) );
NAND3X1 NAND3X1_53 ( .A(_510_), .B(_512_), .C(_511_), .Y(_513_) );
NOR2X1 NOR2X1_53 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_507_) );
AND2X2 AND2X2_53 ( .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_508_) );
OAI21X1 OAI21X1_140 ( .A(_507_), .B(_508_), .C(vdd), .Y(_509_) );
NAND2X1 NAND2X1_141 ( .A(_509_), .B(_513_), .Y(_40__0_) );
OAI21X1 OAI21X1_141 ( .A(_510_), .B(_507_), .C(_512_), .Y(_42__1_) );
INVX1 INVX1_88 ( .A(_42__3_), .Y(_517_) );
OR2X2 OR2X2_54 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_518_) );
NAND2X1 NAND2X1_142 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_519_) );
NAND3X1 NAND3X1_54 ( .A(_517_), .B(_519_), .C(_518_), .Y(_520_) );
NOR2X1 NOR2X1_54 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_514_) );
AND2X2 AND2X2_54 ( .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_515_) );
OAI21X1 OAI21X1_142 ( .A(_514_), .B(_515_), .C(_42__3_), .Y(_516_) );
NAND2X1 NAND2X1_143 ( .A(_516_), .B(_520_), .Y(_40__3_) );
OAI21X1 OAI21X1_143 ( .A(_517_), .B(_514_), .C(_519_), .Y(_38_) );
INVX1 INVX1_89 ( .A(_42__1_), .Y(_524_) );
OR2X2 OR2X2_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_525_) );
NAND2X1 NAND2X1_144 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_526_) );
NAND3X1 NAND3X1_55 ( .A(_524_), .B(_526_), .C(_525_), .Y(_527_) );
NOR2X1 NOR2X1_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_521_) );
AND2X2 AND2X2_55 ( .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_522_) );
OAI21X1 OAI21X1_144 ( .A(_521_), .B(_522_), .C(_42__1_), .Y(_523_) );
NAND2X1 NAND2X1_145 ( .A(_523_), .B(_527_), .Y(_40__1_) );
OAI21X1 OAI21X1_145 ( .A(_524_), .B(_521_), .C(_526_), .Y(_42__2_) );
INVX1 INVX1_90 ( .A(_42__2_), .Y(_531_) );
OR2X2 OR2X2_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_532_) );
NAND2X1 NAND2X1_146 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_533_) );
NAND3X1 NAND3X1_56 ( .A(_531_), .B(_533_), .C(_532_), .Y(_534_) );
NOR2X1 NOR2X1_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_528_) );
AND2X2 AND2X2_56 ( .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_529_) );
OAI21X1 OAI21X1_146 ( .A(_528_), .B(_529_), .C(_42__2_), .Y(_530_) );
NAND2X1 NAND2X1_147 ( .A(_530_), .B(_534_), .Y(_40__2_) );
OAI21X1 OAI21X1_147 ( .A(_531_), .B(_528_), .C(_533_), .Y(_42__3_) );
INVX1 INVX1_91 ( .A(_43_), .Y(_535_) );
NAND2X1 NAND2X1_148 ( .A(_44_), .B(w_cout_7_), .Y(_536_) );
OAI21X1 OAI21X1_148 ( .A(w_cout_7_), .B(_535_), .C(_536_), .Y(w_cout_8_) );
INVX1 INVX1_92 ( .A(_45__0_), .Y(_537_) );
NAND2X1 NAND2X1_149 ( .A(_46__0_), .B(w_cout_7_), .Y(_538_) );
OAI21X1 OAI21X1_149 ( .A(w_cout_7_), .B(_537_), .C(_538_), .Y(_0__32_) );
INVX1 INVX1_93 ( .A(_45__1_), .Y(_539_) );
NAND2X1 NAND2X1_150 ( .A(w_cout_7_), .B(_46__1_), .Y(_540_) );
OAI21X1 OAI21X1_150 ( .A(w_cout_7_), .B(_539_), .C(_540_), .Y(_0__33_) );
INVX1 INVX1_94 ( .A(_45__2_), .Y(_541_) );
NAND2X1 NAND2X1_151 ( .A(w_cout_7_), .B(_46__2_), .Y(_542_) );
OAI21X1 OAI21X1_151 ( .A(w_cout_7_), .B(_541_), .C(_542_), .Y(_0__34_) );
INVX1 INVX1_95 ( .A(_45__3_), .Y(_543_) );
NAND2X1 NAND2X1_152 ( .A(w_cout_7_), .B(_46__3_), .Y(_544_) );
OAI21X1 OAI21X1_152 ( .A(w_cout_7_), .B(_543_), .C(_544_), .Y(_0__35_) );
INVX1 INVX1_96 ( .A(gnd), .Y(_548_) );
OR2X2 OR2X2_57 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_549_) );
NAND2X1 NAND2X1_153 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_550_) );
NAND3X1 NAND3X1_57 ( .A(_548_), .B(_550_), .C(_549_), .Y(_551_) );
NOR2X1 NOR2X1_57 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_545_) );
AND2X2 AND2X2_57 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_546_) );
OAI21X1 OAI21X1_153 ( .A(_545_), .B(_546_), .C(gnd), .Y(_547_) );
NAND2X1 NAND2X1_154 ( .A(_547_), .B(_551_), .Y(_45__0_) );
OAI21X1 OAI21X1_154 ( .A(_548_), .B(_545_), .C(_550_), .Y(_47__1_) );
INVX1 INVX1_97 ( .A(_47__3_), .Y(_555_) );
OR2X2 OR2X2_58 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_556_) );
NAND2X1 NAND2X1_155 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_557_) );
NAND3X1 NAND3X1_58 ( .A(_555_), .B(_557_), .C(_556_), .Y(_558_) );
NOR2X1 NOR2X1_58 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_552_) );
AND2X2 AND2X2_58 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_553_) );
OAI21X1 OAI21X1_155 ( .A(_552_), .B(_553_), .C(_47__3_), .Y(_554_) );
NAND2X1 NAND2X1_156 ( .A(_554_), .B(_558_), .Y(_45__3_) );
OAI21X1 OAI21X1_156 ( .A(_555_), .B(_552_), .C(_557_), .Y(_43_) );
INVX1 INVX1_98 ( .A(_47__1_), .Y(_562_) );
OR2X2 OR2X2_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_563_) );
NAND2X1 NAND2X1_157 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_564_) );
NAND3X1 NAND3X1_59 ( .A(_562_), .B(_564_), .C(_563_), .Y(_565_) );
NOR2X1 NOR2X1_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_559_) );
AND2X2 AND2X2_59 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_560_) );
OAI21X1 OAI21X1_157 ( .A(_559_), .B(_560_), .C(_47__1_), .Y(_561_) );
NAND2X1 NAND2X1_158 ( .A(_561_), .B(_565_), .Y(_45__1_) );
OAI21X1 OAI21X1_158 ( .A(_562_), .B(_559_), .C(_564_), .Y(_47__2_) );
INVX1 INVX1_99 ( .A(_47__2_), .Y(_569_) );
OR2X2 OR2X2_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_570_) );
NAND2X1 NAND2X1_159 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_571_) );
NAND3X1 NAND3X1_60 ( .A(_569_), .B(_571_), .C(_570_), .Y(_572_) );
NOR2X1 NOR2X1_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_566_) );
AND2X2 AND2X2_60 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_567_) );
OAI21X1 OAI21X1_159 ( .A(_566_), .B(_567_), .C(_47__2_), .Y(_568_) );
NAND2X1 NAND2X1_160 ( .A(_568_), .B(_572_), .Y(_45__2_) );
OAI21X1 OAI21X1_160 ( .A(_569_), .B(_566_), .C(_571_), .Y(_47__3_) );
INVX1 INVX1_100 ( .A(vdd), .Y(_576_) );
OR2X2 OR2X2_61 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_577_) );
NAND2X1 NAND2X1_161 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_578_) );
NAND3X1 NAND3X1_61 ( .A(_576_), .B(_578_), .C(_577_), .Y(_579_) );
NOR2X1 NOR2X1_61 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_573_) );
AND2X2 AND2X2_61 ( .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_574_) );
OAI21X1 OAI21X1_161 ( .A(_573_), .B(_574_), .C(vdd), .Y(_575_) );
NAND2X1 NAND2X1_162 ( .A(_575_), .B(_579_), .Y(_46__0_) );
OAI21X1 OAI21X1_162 ( .A(_576_), .B(_573_), .C(_578_), .Y(_48__1_) );
INVX1 INVX1_101 ( .A(_48__3_), .Y(_583_) );
OR2X2 OR2X2_62 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_584_) );
NAND2X1 NAND2X1_163 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_585_) );
NAND3X1 NAND3X1_62 ( .A(_583_), .B(_585_), .C(_584_), .Y(_586_) );
NOR2X1 NOR2X1_62 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_580_) );
AND2X2 AND2X2_62 ( .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_581_) );
OAI21X1 OAI21X1_163 ( .A(_580_), .B(_581_), .C(_48__3_), .Y(_582_) );
NAND2X1 NAND2X1_164 ( .A(_582_), .B(_586_), .Y(_46__3_) );
OAI21X1 OAI21X1_164 ( .A(_583_), .B(_580_), .C(_585_), .Y(_44_) );
INVX1 INVX1_102 ( .A(_48__1_), .Y(_590_) );
OR2X2 OR2X2_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_591_) );
NAND2X1 NAND2X1_165 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_592_) );
NAND3X1 NAND3X1_63 ( .A(_590_), .B(_592_), .C(_591_), .Y(_593_) );
NOR2X1 NOR2X1_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_587_) );
AND2X2 AND2X2_63 ( .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_588_) );
OAI21X1 OAI21X1_165 ( .A(_587_), .B(_588_), .C(_48__1_), .Y(_589_) );
NAND2X1 NAND2X1_166 ( .A(_589_), .B(_593_), .Y(_46__1_) );
OAI21X1 OAI21X1_166 ( .A(_590_), .B(_587_), .C(_592_), .Y(_48__2_) );
INVX1 INVX1_103 ( .A(_48__2_), .Y(_597_) );
OR2X2 OR2X2_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_598_) );
NAND2X1 NAND2X1_167 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_599_) );
NAND3X1 NAND3X1_64 ( .A(_597_), .B(_599_), .C(_598_), .Y(_600_) );
NOR2X1 NOR2X1_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_594_) );
AND2X2 AND2X2_64 ( .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_595_) );
OAI21X1 OAI21X1_167 ( .A(_594_), .B(_595_), .C(_48__2_), .Y(_596_) );
NAND2X1 NAND2X1_168 ( .A(_596_), .B(_600_), .Y(_46__2_) );
OAI21X1 OAI21X1_168 ( .A(_597_), .B(_594_), .C(_599_), .Y(_48__3_) );
INVX1 INVX1_104 ( .A(_49_), .Y(_601_) );
NAND2X1 NAND2X1_169 ( .A(_50_), .B(w_cout_8_), .Y(_602_) );
OAI21X1 OAI21X1_169 ( .A(w_cout_8_), .B(_601_), .C(_602_), .Y(w_cout_9_) );
INVX1 INVX1_105 ( .A(_51__0_), .Y(_603_) );
NAND2X1 NAND2X1_170 ( .A(_52__0_), .B(w_cout_8_), .Y(_604_) );
OAI21X1 OAI21X1_170 ( .A(w_cout_8_), .B(_603_), .C(_604_), .Y(_0__36_) );
INVX1 INVX1_106 ( .A(_51__1_), .Y(_605_) );
NAND2X1 NAND2X1_171 ( .A(w_cout_8_), .B(_52__1_), .Y(_606_) );
OAI21X1 OAI21X1_171 ( .A(w_cout_8_), .B(_605_), .C(_606_), .Y(_0__37_) );
INVX1 INVX1_107 ( .A(_51__2_), .Y(_607_) );
NAND2X1 NAND2X1_172 ( .A(w_cout_8_), .B(_52__2_), .Y(_608_) );
OAI21X1 OAI21X1_172 ( .A(w_cout_8_), .B(_607_), .C(_608_), .Y(_0__38_) );
INVX1 INVX1_108 ( .A(_51__3_), .Y(_609_) );
NAND2X1 NAND2X1_173 ( .A(w_cout_8_), .B(_52__3_), .Y(_610_) );
OAI21X1 OAI21X1_173 ( .A(w_cout_8_), .B(_609_), .C(_610_), .Y(_0__39_) );
INVX1 INVX1_109 ( .A(gnd), .Y(_614_) );
OR2X2 OR2X2_65 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_615_) );
NAND2X1 NAND2X1_174 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_616_) );
NAND3X1 NAND3X1_65 ( .A(_614_), .B(_616_), .C(_615_), .Y(_617_) );
NOR2X1 NOR2X1_65 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_611_) );
AND2X2 AND2X2_65 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_612_) );
OAI21X1 OAI21X1_174 ( .A(_611_), .B(_612_), .C(gnd), .Y(_613_) );
NAND2X1 NAND2X1_175 ( .A(_613_), .B(_617_), .Y(_51__0_) );
OAI21X1 OAI21X1_175 ( .A(_614_), .B(_611_), .C(_616_), .Y(_53__1_) );
INVX1 INVX1_110 ( .A(_53__3_), .Y(_621_) );
OR2X2 OR2X2_66 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_622_) );
NAND2X1 NAND2X1_176 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_623_) );
NAND3X1 NAND3X1_66 ( .A(_621_), .B(_623_), .C(_622_), .Y(_624_) );
NOR2X1 NOR2X1_66 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_618_) );
AND2X2 AND2X2_66 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_619_) );
OAI21X1 OAI21X1_176 ( .A(_618_), .B(_619_), .C(_53__3_), .Y(_620_) );
NAND2X1 NAND2X1_177 ( .A(_620_), .B(_624_), .Y(_51__3_) );
OAI21X1 OAI21X1_177 ( .A(_621_), .B(_618_), .C(_623_), .Y(_49_) );
INVX1 INVX1_111 ( .A(_53__1_), .Y(_628_) );
OR2X2 OR2X2_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_629_) );
NAND2X1 NAND2X1_178 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_630_) );
NAND3X1 NAND3X1_67 ( .A(_628_), .B(_630_), .C(_629_), .Y(_631_) );
NOR2X1 NOR2X1_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_625_) );
AND2X2 AND2X2_67 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_626_) );
OAI21X1 OAI21X1_178 ( .A(_625_), .B(_626_), .C(_53__1_), .Y(_627_) );
NAND2X1 NAND2X1_179 ( .A(_627_), .B(_631_), .Y(_51__1_) );
OAI21X1 OAI21X1_179 ( .A(_628_), .B(_625_), .C(_630_), .Y(_53__2_) );
INVX1 INVX1_112 ( .A(_53__2_), .Y(_635_) );
OR2X2 OR2X2_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_636_) );
NAND2X1 NAND2X1_180 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_637_) );
NAND3X1 NAND3X1_68 ( .A(_635_), .B(_637_), .C(_636_), .Y(_638_) );
NOR2X1 NOR2X1_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_632_) );
AND2X2 AND2X2_68 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_633_) );
OAI21X1 OAI21X1_180 ( .A(_632_), .B(_633_), .C(_53__2_), .Y(_634_) );
NAND2X1 NAND2X1_181 ( .A(_634_), .B(_638_), .Y(_51__2_) );
OAI21X1 OAI21X1_181 ( .A(_635_), .B(_632_), .C(_637_), .Y(_53__3_) );
INVX1 INVX1_113 ( .A(vdd), .Y(_642_) );
OR2X2 OR2X2_69 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_643_) );
NAND2X1 NAND2X1_182 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_644_) );
NAND3X1 NAND3X1_69 ( .A(_642_), .B(_644_), .C(_643_), .Y(_645_) );
NOR2X1 NOR2X1_69 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_639_) );
AND2X2 AND2X2_69 ( .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_640_) );
OAI21X1 OAI21X1_182 ( .A(_639_), .B(_640_), .C(vdd), .Y(_641_) );
NAND2X1 NAND2X1_183 ( .A(_641_), .B(_645_), .Y(_52__0_) );
OAI21X1 OAI21X1_183 ( .A(_642_), .B(_639_), .C(_644_), .Y(_54__1_) );
INVX1 INVX1_114 ( .A(_54__3_), .Y(_649_) );
OR2X2 OR2X2_70 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_650_) );
NAND2X1 NAND2X1_184 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_651_) );
NAND3X1 NAND3X1_70 ( .A(_649_), .B(_651_), .C(_650_), .Y(_652_) );
NOR2X1 NOR2X1_70 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_646_) );
AND2X2 AND2X2_70 ( .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_647_) );
OAI21X1 OAI21X1_184 ( .A(_646_), .B(_647_), .C(_54__3_), .Y(_648_) );
NAND2X1 NAND2X1_185 ( .A(_648_), .B(_652_), .Y(_52__3_) );
OAI21X1 OAI21X1_185 ( .A(_649_), .B(_646_), .C(_651_), .Y(_50_) );
INVX1 INVX1_115 ( .A(_54__1_), .Y(_656_) );
OR2X2 OR2X2_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_657_) );
NAND2X1 NAND2X1_186 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_658_) );
NAND3X1 NAND3X1_71 ( .A(_656_), .B(_658_), .C(_657_), .Y(_659_) );
NOR2X1 NOR2X1_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_653_) );
AND2X2 AND2X2_71 ( .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_654_) );
OAI21X1 OAI21X1_186 ( .A(_653_), .B(_654_), .C(_54__1_), .Y(_655_) );
NAND2X1 NAND2X1_187 ( .A(_655_), .B(_659_), .Y(_52__1_) );
OAI21X1 OAI21X1_187 ( .A(_656_), .B(_653_), .C(_658_), .Y(_54__2_) );
INVX1 INVX1_116 ( .A(_54__2_), .Y(_663_) );
OR2X2 OR2X2_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_664_) );
NAND2X1 NAND2X1_188 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_665_) );
NAND3X1 NAND3X1_72 ( .A(_663_), .B(_665_), .C(_664_), .Y(_666_) );
NOR2X1 NOR2X1_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_660_) );
AND2X2 AND2X2_72 ( .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_661_) );
OAI21X1 OAI21X1_188 ( .A(_660_), .B(_661_), .C(_54__2_), .Y(_662_) );
NAND2X1 NAND2X1_189 ( .A(_662_), .B(_666_), .Y(_52__2_) );
OAI21X1 OAI21X1_189 ( .A(_663_), .B(_660_), .C(_665_), .Y(_54__3_) );
INVX1 INVX1_117 ( .A(_55_), .Y(_667_) );
NAND2X1 NAND2X1_190 ( .A(_56_), .B(w_cout_9_), .Y(_668_) );
OAI21X1 OAI21X1_190 ( .A(w_cout_9_), .B(_667_), .C(_668_), .Y(w_cout_10_) );
INVX1 INVX1_118 ( .A(_57__0_), .Y(_669_) );
NAND2X1 NAND2X1_191 ( .A(_58__0_), .B(w_cout_9_), .Y(_670_) );
OAI21X1 OAI21X1_191 ( .A(w_cout_9_), .B(_669_), .C(_670_), .Y(_0__40_) );
INVX1 INVX1_119 ( .A(_57__1_), .Y(_671_) );
NAND2X1 NAND2X1_192 ( .A(w_cout_9_), .B(_58__1_), .Y(_672_) );
OAI21X1 OAI21X1_192 ( .A(w_cout_9_), .B(_671_), .C(_672_), .Y(_0__41_) );
INVX1 INVX1_120 ( .A(_57__2_), .Y(_673_) );
NAND2X1 NAND2X1_193 ( .A(w_cout_9_), .B(_58__2_), .Y(_674_) );
OAI21X1 OAI21X1_193 ( .A(w_cout_9_), .B(_673_), .C(_674_), .Y(_0__42_) );
INVX1 INVX1_121 ( .A(_57__3_), .Y(_675_) );
NAND2X1 NAND2X1_194 ( .A(w_cout_9_), .B(_58__3_), .Y(_676_) );
OAI21X1 OAI21X1_194 ( .A(w_cout_9_), .B(_675_), .C(_676_), .Y(_0__43_) );
INVX1 INVX1_122 ( .A(gnd), .Y(_680_) );
OR2X2 OR2X2_73 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_681_) );
NAND2X1 NAND2X1_195 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_682_) );
NAND3X1 NAND3X1_73 ( .A(_680_), .B(_682_), .C(_681_), .Y(_683_) );
NOR2X1 NOR2X1_73 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_677_) );
AND2X2 AND2X2_73 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_678_) );
OAI21X1 OAI21X1_195 ( .A(_677_), .B(_678_), .C(gnd), .Y(_679_) );
NAND2X1 NAND2X1_196 ( .A(_679_), .B(_683_), .Y(_57__0_) );
OAI21X1 OAI21X1_196 ( .A(_680_), .B(_677_), .C(_682_), .Y(_59__1_) );
INVX1 INVX1_123 ( .A(_59__3_), .Y(_687_) );
OR2X2 OR2X2_74 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_688_) );
NAND2X1 NAND2X1_197 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_689_) );
NAND3X1 NAND3X1_74 ( .A(_687_), .B(_689_), .C(_688_), .Y(_690_) );
NOR2X1 NOR2X1_74 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_684_) );
AND2X2 AND2X2_74 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_685_) );
OAI21X1 OAI21X1_197 ( .A(_684_), .B(_685_), .C(_59__3_), .Y(_686_) );
NAND2X1 NAND2X1_198 ( .A(_686_), .B(_690_), .Y(_57__3_) );
OAI21X1 OAI21X1_198 ( .A(_687_), .B(_684_), .C(_689_), .Y(_55_) );
INVX1 INVX1_124 ( .A(_59__1_), .Y(_694_) );
OR2X2 OR2X2_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_695_) );
NAND2X1 NAND2X1_199 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_696_) );
NAND3X1 NAND3X1_75 ( .A(_694_), .B(_696_), .C(_695_), .Y(_697_) );
NOR2X1 NOR2X1_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_691_) );
AND2X2 AND2X2_75 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_692_) );
OAI21X1 OAI21X1_199 ( .A(_691_), .B(_692_), .C(_59__1_), .Y(_693_) );
NAND2X1 NAND2X1_200 ( .A(_693_), .B(_697_), .Y(_57__1_) );
OAI21X1 OAI21X1_200 ( .A(_694_), .B(_691_), .C(_696_), .Y(_59__2_) );
INVX1 INVX1_125 ( .A(_59__2_), .Y(_701_) );
OR2X2 OR2X2_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_702_) );
NAND2X1 NAND2X1_201 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_703_) );
NAND3X1 NAND3X1_76 ( .A(_701_), .B(_703_), .C(_702_), .Y(_704_) );
NOR2X1 NOR2X1_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_698_) );
AND2X2 AND2X2_76 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_699_) );
OAI21X1 OAI21X1_201 ( .A(_698_), .B(_699_), .C(_59__2_), .Y(_700_) );
NAND2X1 NAND2X1_202 ( .A(_700_), .B(_704_), .Y(_57__2_) );
OAI21X1 OAI21X1_202 ( .A(_701_), .B(_698_), .C(_703_), .Y(_59__3_) );
INVX1 INVX1_126 ( .A(vdd), .Y(_708_) );
OR2X2 OR2X2_77 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_709_) );
NAND2X1 NAND2X1_203 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_710_) );
NAND3X1 NAND3X1_77 ( .A(_708_), .B(_710_), .C(_709_), .Y(_711_) );
NOR2X1 NOR2X1_77 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_705_) );
AND2X2 AND2X2_77 ( .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_706_) );
OAI21X1 OAI21X1_203 ( .A(_705_), .B(_706_), .C(vdd), .Y(_707_) );
NAND2X1 NAND2X1_204 ( .A(_707_), .B(_711_), .Y(_58__0_) );
OAI21X1 OAI21X1_204 ( .A(_708_), .B(_705_), .C(_710_), .Y(_60__1_) );
INVX1 INVX1_127 ( .A(_60__3_), .Y(_715_) );
OR2X2 OR2X2_78 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_716_) );
NAND2X1 NAND2X1_205 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_717_) );
NAND3X1 NAND3X1_78 ( .A(_715_), .B(_717_), .C(_716_), .Y(_718_) );
NOR2X1 NOR2X1_78 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_712_) );
AND2X2 AND2X2_78 ( .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_713_) );
OAI21X1 OAI21X1_205 ( .A(_712_), .B(_713_), .C(_60__3_), .Y(_714_) );
NAND2X1 NAND2X1_206 ( .A(_714_), .B(_718_), .Y(_58__3_) );
OAI21X1 OAI21X1_206 ( .A(_715_), .B(_712_), .C(_717_), .Y(_56_) );
INVX1 INVX1_128 ( .A(_60__1_), .Y(_722_) );
OR2X2 OR2X2_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_723_) );
NAND2X1 NAND2X1_207 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_724_) );
NAND3X1 NAND3X1_79 ( .A(_722_), .B(_724_), .C(_723_), .Y(_725_) );
NOR2X1 NOR2X1_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_719_) );
AND2X2 AND2X2_79 ( .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_720_) );
OAI21X1 OAI21X1_207 ( .A(_719_), .B(_720_), .C(_60__1_), .Y(_721_) );
NAND2X1 NAND2X1_208 ( .A(_721_), .B(_725_), .Y(_58__1_) );
OAI21X1 OAI21X1_208 ( .A(_722_), .B(_719_), .C(_724_), .Y(_60__2_) );
INVX1 INVX1_129 ( .A(_60__2_), .Y(_729_) );
OR2X2 OR2X2_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_730_) );
NAND2X1 NAND2X1_209 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_731_) );
NAND3X1 NAND3X1_80 ( .A(_729_), .B(_731_), .C(_730_), .Y(_732_) );
NOR2X1 NOR2X1_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_726_) );
AND2X2 AND2X2_80 ( .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_727_) );
OAI21X1 OAI21X1_209 ( .A(_726_), .B(_727_), .C(_60__2_), .Y(_728_) );
NAND2X1 NAND2X1_210 ( .A(_728_), .B(_732_), .Y(_58__2_) );
OAI21X1 OAI21X1_210 ( .A(_729_), .B(_726_), .C(_731_), .Y(_60__3_) );
INVX1 INVX1_130 ( .A(_61_), .Y(_733_) );
NAND2X1 NAND2X1_211 ( .A(_62_), .B(w_cout_10_), .Y(_734_) );
OAI21X1 OAI21X1_211 ( .A(w_cout_10_), .B(_733_), .C(_734_), .Y(w_cout_11_) );
INVX1 INVX1_131 ( .A(_63__0_), .Y(_735_) );
NAND2X1 NAND2X1_212 ( .A(_64__0_), .B(w_cout_10_), .Y(_736_) );
OAI21X1 OAI21X1_212 ( .A(w_cout_10_), .B(_735_), .C(_736_), .Y(_0__44_) );
INVX1 INVX1_132 ( .A(_63__1_), .Y(_737_) );
NAND2X1 NAND2X1_213 ( .A(w_cout_10_), .B(_64__1_), .Y(_738_) );
OAI21X1 OAI21X1_213 ( .A(w_cout_10_), .B(_737_), .C(_738_), .Y(_0__45_) );
INVX1 INVX1_133 ( .A(_63__2_), .Y(_739_) );
NAND2X1 NAND2X1_214 ( .A(w_cout_10_), .B(_64__2_), .Y(_740_) );
OAI21X1 OAI21X1_214 ( .A(w_cout_10_), .B(_739_), .C(_740_), .Y(_0__46_) );
INVX1 INVX1_134 ( .A(_63__3_), .Y(_741_) );
NAND2X1 NAND2X1_215 ( .A(w_cout_10_), .B(_64__3_), .Y(_742_) );
OAI21X1 OAI21X1_215 ( .A(w_cout_10_), .B(_741_), .C(_742_), .Y(_0__47_) );
INVX1 INVX1_135 ( .A(gnd), .Y(_746_) );
OR2X2 OR2X2_81 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_747_) );
NAND2X1 NAND2X1_216 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_748_) );
NAND3X1 NAND3X1_81 ( .A(_746_), .B(_748_), .C(_747_), .Y(_749_) );
NOR2X1 NOR2X1_81 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_743_) );
AND2X2 AND2X2_81 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_744_) );
OAI21X1 OAI21X1_216 ( .A(_743_), .B(_744_), .C(gnd), .Y(_745_) );
NAND2X1 NAND2X1_217 ( .A(_745_), .B(_749_), .Y(_63__0_) );
OAI21X1 OAI21X1_217 ( .A(_746_), .B(_743_), .C(_748_), .Y(_65__1_) );
INVX1 INVX1_136 ( .A(_65__3_), .Y(_753_) );
OR2X2 OR2X2_82 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_754_) );
NAND2X1 NAND2X1_218 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_755_) );
NAND3X1 NAND3X1_82 ( .A(_753_), .B(_755_), .C(_754_), .Y(_756_) );
NOR2X1 NOR2X1_82 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_750_) );
AND2X2 AND2X2_82 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_751_) );
OAI21X1 OAI21X1_218 ( .A(_750_), .B(_751_), .C(_65__3_), .Y(_752_) );
NAND2X1 NAND2X1_219 ( .A(_752_), .B(_756_), .Y(_63__3_) );
OAI21X1 OAI21X1_219 ( .A(_753_), .B(_750_), .C(_755_), .Y(_61_) );
INVX1 INVX1_137 ( .A(_65__1_), .Y(_760_) );
OR2X2 OR2X2_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_761_) );
NAND2X1 NAND2X1_220 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_762_) );
NAND3X1 NAND3X1_83 ( .A(_760_), .B(_762_), .C(_761_), .Y(_763_) );
NOR2X1 NOR2X1_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_757_) );
AND2X2 AND2X2_83 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_758_) );
OAI21X1 OAI21X1_220 ( .A(_757_), .B(_758_), .C(_65__1_), .Y(_759_) );
NAND2X1 NAND2X1_221 ( .A(_759_), .B(_763_), .Y(_63__1_) );
OAI21X1 OAI21X1_221 ( .A(_760_), .B(_757_), .C(_762_), .Y(_65__2_) );
INVX1 INVX1_138 ( .A(_65__2_), .Y(_767_) );
OR2X2 OR2X2_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_768_) );
NAND2X1 NAND2X1_222 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_769_) );
NAND3X1 NAND3X1_84 ( .A(_767_), .B(_769_), .C(_768_), .Y(_770_) );
NOR2X1 NOR2X1_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_764_) );
AND2X2 AND2X2_84 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_765_) );
OAI21X1 OAI21X1_222 ( .A(_764_), .B(_765_), .C(_65__2_), .Y(_766_) );
NAND2X1 NAND2X1_223 ( .A(_766_), .B(_770_), .Y(_63__2_) );
OAI21X1 OAI21X1_223 ( .A(_767_), .B(_764_), .C(_769_), .Y(_65__3_) );
INVX1 INVX1_139 ( .A(vdd), .Y(_774_) );
OR2X2 OR2X2_85 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_775_) );
NAND2X1 NAND2X1_224 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_776_) );
NAND3X1 NAND3X1_85 ( .A(_774_), .B(_776_), .C(_775_), .Y(_777_) );
NOR2X1 NOR2X1_85 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_771_) );
AND2X2 AND2X2_85 ( .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_772_) );
OAI21X1 OAI21X1_224 ( .A(_771_), .B(_772_), .C(vdd), .Y(_773_) );
NAND2X1 NAND2X1_225 ( .A(_773_), .B(_777_), .Y(_64__0_) );
OAI21X1 OAI21X1_225 ( .A(_774_), .B(_771_), .C(_776_), .Y(_66__1_) );
INVX1 INVX1_140 ( .A(_66__3_), .Y(_781_) );
OR2X2 OR2X2_86 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_782_) );
NAND2X1 NAND2X1_226 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_783_) );
NAND3X1 NAND3X1_86 ( .A(_781_), .B(_783_), .C(_782_), .Y(_784_) );
NOR2X1 NOR2X1_86 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_778_) );
AND2X2 AND2X2_86 ( .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_779_) );
OAI21X1 OAI21X1_226 ( .A(_778_), .B(_779_), .C(_66__3_), .Y(_780_) );
NAND2X1 NAND2X1_227 ( .A(_780_), .B(_784_), .Y(_64__3_) );
OAI21X1 OAI21X1_227 ( .A(_781_), .B(_778_), .C(_783_), .Y(_62_) );
INVX1 INVX1_141 ( .A(_66__1_), .Y(_788_) );
OR2X2 OR2X2_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_789_) );
NAND2X1 NAND2X1_228 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_790_) );
NAND3X1 NAND3X1_87 ( .A(_788_), .B(_790_), .C(_789_), .Y(_791_) );
NOR2X1 NOR2X1_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_785_) );
AND2X2 AND2X2_87 ( .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_786_) );
OAI21X1 OAI21X1_228 ( .A(_785_), .B(_786_), .C(_66__1_), .Y(_787_) );
NAND2X1 NAND2X1_229 ( .A(_787_), .B(_791_), .Y(_64__1_) );
OAI21X1 OAI21X1_229 ( .A(_788_), .B(_785_), .C(_790_), .Y(_66__2_) );
INVX1 INVX1_142 ( .A(_66__2_), .Y(_795_) );
OR2X2 OR2X2_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_796_) );
NAND2X1 NAND2X1_230 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_797_) );
NAND3X1 NAND3X1_88 ( .A(_795_), .B(_797_), .C(_796_), .Y(_798_) );
NOR2X1 NOR2X1_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_792_) );
AND2X2 AND2X2_88 ( .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_793_) );
OAI21X1 OAI21X1_230 ( .A(_792_), .B(_793_), .C(_66__2_), .Y(_794_) );
NAND2X1 NAND2X1_231 ( .A(_794_), .B(_798_), .Y(_64__2_) );
OAI21X1 OAI21X1_231 ( .A(_795_), .B(_792_), .C(_797_), .Y(_66__3_) );
INVX1 INVX1_143 ( .A(_67_), .Y(_799_) );
NAND2X1 NAND2X1_232 ( .A(_68_), .B(w_cout_11_), .Y(_800_) );
OAI21X1 OAI21X1_232 ( .A(w_cout_11_), .B(_799_), .C(_800_), .Y(csa_inst_cin) );
INVX1 INVX1_144 ( .A(_69__0_), .Y(_801_) );
NAND2X1 NAND2X1_233 ( .A(_70__0_), .B(w_cout_11_), .Y(_802_) );
OAI21X1 OAI21X1_233 ( .A(w_cout_11_), .B(_801_), .C(_802_), .Y(_0__48_) );
INVX1 INVX1_145 ( .A(_69__1_), .Y(_803_) );
NAND2X1 NAND2X1_234 ( .A(w_cout_11_), .B(_70__1_), .Y(_804_) );
OAI21X1 OAI21X1_234 ( .A(w_cout_11_), .B(_803_), .C(_804_), .Y(_0__49_) );
INVX1 INVX1_146 ( .A(_69__2_), .Y(_805_) );
NAND2X1 NAND2X1_235 ( .A(w_cout_11_), .B(_70__2_), .Y(_806_) );
OAI21X1 OAI21X1_235 ( .A(w_cout_11_), .B(_805_), .C(_806_), .Y(_0__50_) );
INVX1 INVX1_147 ( .A(_69__3_), .Y(_807_) );
NAND2X1 NAND2X1_236 ( .A(w_cout_11_), .B(_70__3_), .Y(_808_) );
OAI21X1 OAI21X1_236 ( .A(w_cout_11_), .B(_807_), .C(_808_), .Y(_0__51_) );
INVX1 INVX1_148 ( .A(gnd), .Y(_812_) );
OR2X2 OR2X2_89 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_813_) );
NAND2X1 NAND2X1_237 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_814_) );
NAND3X1 NAND3X1_89 ( .A(_812_), .B(_814_), .C(_813_), .Y(_815_) );
NOR2X1 NOR2X1_89 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_809_) );
AND2X2 AND2X2_89 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_810_) );
OAI21X1 OAI21X1_237 ( .A(_809_), .B(_810_), .C(gnd), .Y(_811_) );
NAND2X1 NAND2X1_238 ( .A(_811_), .B(_815_), .Y(_69__0_) );
OAI21X1 OAI21X1_238 ( .A(_812_), .B(_809_), .C(_814_), .Y(_71__1_) );
INVX1 INVX1_149 ( .A(_71__3_), .Y(_819_) );
OR2X2 OR2X2_90 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_820_) );
NAND2X1 NAND2X1_239 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_821_) );
NAND3X1 NAND3X1_90 ( .A(_819_), .B(_821_), .C(_820_), .Y(_822_) );
NOR2X1 NOR2X1_90 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_816_) );
AND2X2 AND2X2_90 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_817_) );
OAI21X1 OAI21X1_239 ( .A(_816_), .B(_817_), .C(_71__3_), .Y(_818_) );
NAND2X1 NAND2X1_240 ( .A(_818_), .B(_822_), .Y(_69__3_) );
OAI21X1 OAI21X1_240 ( .A(_819_), .B(_816_), .C(_821_), .Y(_67_) );
INVX1 INVX1_150 ( .A(_71__1_), .Y(_826_) );
OR2X2 OR2X2_91 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_827_) );
NAND2X1 NAND2X1_241 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_828_) );
NAND3X1 NAND3X1_91 ( .A(_826_), .B(_828_), .C(_827_), .Y(_829_) );
NOR2X1 NOR2X1_91 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_823_) );
AND2X2 AND2X2_91 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_824_) );
OAI21X1 OAI21X1_241 ( .A(_823_), .B(_824_), .C(_71__1_), .Y(_825_) );
NAND2X1 NAND2X1_242 ( .A(_825_), .B(_829_), .Y(_69__1_) );
OAI21X1 OAI21X1_242 ( .A(_826_), .B(_823_), .C(_828_), .Y(_71__2_) );
INVX1 INVX1_151 ( .A(_71__2_), .Y(_833_) );
OR2X2 OR2X2_92 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_834_) );
NAND2X1 NAND2X1_243 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_835_) );
NAND3X1 NAND3X1_92 ( .A(_833_), .B(_835_), .C(_834_), .Y(_836_) );
NOR2X1 NOR2X1_92 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_830_) );
AND2X2 AND2X2_92 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_831_) );
OAI21X1 OAI21X1_243 ( .A(_830_), .B(_831_), .C(_71__2_), .Y(_832_) );
NAND2X1 NAND2X1_244 ( .A(_832_), .B(_836_), .Y(_69__2_) );
OAI21X1 OAI21X1_244 ( .A(_833_), .B(_830_), .C(_835_), .Y(_71__3_) );
INVX1 INVX1_152 ( .A(vdd), .Y(_840_) );
OR2X2 OR2X2_93 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_841_) );
NAND2X1 NAND2X1_245 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_842_) );
NAND3X1 NAND3X1_93 ( .A(_840_), .B(_842_), .C(_841_), .Y(_843_) );
NOR2X1 NOR2X1_93 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_837_) );
AND2X2 AND2X2_93 ( .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_838_) );
OAI21X1 OAI21X1_245 ( .A(_837_), .B(_838_), .C(vdd), .Y(_839_) );
NAND2X1 NAND2X1_246 ( .A(_839_), .B(_843_), .Y(_70__0_) );
OAI21X1 OAI21X1_246 ( .A(_840_), .B(_837_), .C(_842_), .Y(_72__1_) );
INVX1 INVX1_153 ( .A(_72__3_), .Y(_847_) );
OR2X2 OR2X2_94 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_848_) );
NAND2X1 NAND2X1_247 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_849_) );
NAND3X1 NAND3X1_94 ( .A(_847_), .B(_849_), .C(_848_), .Y(_850_) );
NOR2X1 NOR2X1_94 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_844_) );
AND2X2 AND2X2_94 ( .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_845_) );
OAI21X1 OAI21X1_247 ( .A(_844_), .B(_845_), .C(_72__3_), .Y(_846_) );
NAND2X1 NAND2X1_248 ( .A(_846_), .B(_850_), .Y(_70__3_) );
OAI21X1 OAI21X1_248 ( .A(_847_), .B(_844_), .C(_849_), .Y(_68_) );
INVX1 INVX1_154 ( .A(_72__1_), .Y(_854_) );
OR2X2 OR2X2_95 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_855_) );
NAND2X1 NAND2X1_249 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_856_) );
NAND3X1 NAND3X1_95 ( .A(_854_), .B(_856_), .C(_855_), .Y(_857_) );
NOR2X1 NOR2X1_95 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_851_) );
AND2X2 AND2X2_95 ( .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_852_) );
OAI21X1 OAI21X1_249 ( .A(_851_), .B(_852_), .C(_72__1_), .Y(_853_) );
NAND2X1 NAND2X1_250 ( .A(_853_), .B(_857_), .Y(_70__1_) );
OAI21X1 OAI21X1_250 ( .A(_854_), .B(_851_), .C(_856_), .Y(_72__2_) );
INVX1 INVX1_155 ( .A(_72__2_), .Y(_861_) );
OR2X2 OR2X2_96 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_862_) );
NAND2X1 NAND2X1_251 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_863_) );
NAND3X1 NAND3X1_96 ( .A(_861_), .B(_863_), .C(_862_), .Y(_864_) );
NOR2X1 NOR2X1_96 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_858_) );
AND2X2 AND2X2_96 ( .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_859_) );
OAI21X1 OAI21X1_251 ( .A(_858_), .B(_859_), .C(_72__2_), .Y(_860_) );
NAND2X1 NAND2X1_252 ( .A(_860_), .B(_864_), .Y(_70__2_) );
OAI21X1 OAI21X1_252 ( .A(_861_), .B(_858_), .C(_863_), .Y(_72__3_) );
INVX1 INVX1_156 ( .A(csa_inst_cout0_0), .Y(_865_) );
NAND2X1 NAND2X1_253 ( .A(csa_inst_cout0_1), .B(csa_inst_cin), .Y(_866_) );
OAI21X1 OAI21X1_253 ( .A(csa_inst_cin), .B(_865_), .C(_866_), .Y(w_cout_13_) );
INVX1 INVX1_157 ( .A(csa_inst_rca0_0_fa0_o_sum), .Y(_867_) );
NAND2X1 NAND2X1_254 ( .A(csa_inst_rca0_1_fa0_o_sum), .B(csa_inst_cin), .Y(_868_) );
OAI21X1 OAI21X1_254 ( .A(csa_inst_cin), .B(_867_), .C(_868_), .Y(_0__52_) );
INVX1 INVX1_158 ( .A(csa_inst_rca0_0_fa1_o_sum), .Y(_869_) );
NAND2X1 NAND2X1_255 ( .A(csa_inst_cin), .B(csa_inst_rca0_1_fa1_o_sum), .Y(_870_) );
OAI21X1 OAI21X1_255 ( .A(csa_inst_cin), .B(_869_), .C(_870_), .Y(_0__53_) );
INVX1 INVX1_159 ( .A(csa_inst_rca0_0_fa2_o_sum), .Y(_871_) );
NAND2X1 NAND2X1_256 ( .A(csa_inst_cin), .B(csa_inst_rca0_1_fa2_o_sum), .Y(_872_) );
OAI21X1 OAI21X1_256 ( .A(csa_inst_cin), .B(_871_), .C(_872_), .Y(_0__54_) );
INVX1 INVX1_160 ( .A(gnd), .Y(_876_) );
OR2X2 OR2X2_97 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_877_) );
NAND2X1 NAND2X1_257 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_878_) );
NAND3X1 NAND3X1_97 ( .A(_876_), .B(_878_), .C(_877_), .Y(_879_) );
NOR2X1 NOR2X1_97 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_873_) );
AND2X2 AND2X2_97 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_874_) );
OAI21X1 OAI21X1_257 ( .A(_873_), .B(_874_), .C(gnd), .Y(_875_) );
NAND2X1 NAND2X1_258 ( .A(_875_), .B(_879_), .Y(csa_inst_rca0_0_fa0_o_sum) );
OAI21X1 OAI21X1_258 ( .A(_876_), .B(_873_), .C(_878_), .Y(csa_inst_rca0_0_fa0_o_carry) );
INVX1 INVX1_161 ( .A(csa_inst_rca0_0_fa0_o_carry), .Y(_883_) );
OR2X2 OR2X2_98 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_884_) );
NAND2X1 NAND2X1_259 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_885_) );
NAND3X1 NAND3X1_98 ( .A(_883_), .B(_885_), .C(_884_), .Y(_886_) );
NOR2X1 NOR2X1_98 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_880_) );
AND2X2 AND2X2_98 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_881_) );
OAI21X1 OAI21X1_259 ( .A(_880_), .B(_881_), .C(csa_inst_rca0_0_fa0_o_carry), .Y(_882_) );
NAND2X1 NAND2X1_260 ( .A(_882_), .B(_886_), .Y(csa_inst_rca0_0_fa1_o_sum) );
OAI21X1 OAI21X1_260 ( .A(_883_), .B(_880_), .C(_885_), .Y(csa_inst_rca0_0_fa1_o_carry) );
INVX1 INVX1_162 ( .A(csa_inst_rca0_0_fa1_o_carry), .Y(_890_) );
OR2X2 OR2X2_99 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_891_) );
NAND2X1 NAND2X1_261 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_892_) );
NAND3X1 NAND3X1_99 ( .A(_890_), .B(_892_), .C(_891_), .Y(_893_) );
NOR2X1 NOR2X1_99 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_887_) );
AND2X2 AND2X2_99 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_888_) );
OAI21X1 OAI21X1_261 ( .A(_887_), .B(_888_), .C(csa_inst_rca0_0_fa1_o_carry), .Y(_889_) );
NAND2X1 NAND2X1_262 ( .A(_889_), .B(_893_), .Y(csa_inst_rca0_0_fa2_o_sum) );
OAI21X1 OAI21X1_262 ( .A(_890_), .B(_887_), .C(_892_), .Y(csa_inst_cout0_0) );
INVX1 INVX1_163 ( .A(vdd), .Y(_897_) );
OR2X2 OR2X2_100 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_898_) );
NAND2X1 NAND2X1_263 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_899_) );
NAND3X1 NAND3X1_100 ( .A(_897_), .B(_899_), .C(_898_), .Y(_900_) );
NOR2X1 NOR2X1_100 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_894_) );
AND2X2 AND2X2_100 ( .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_895_) );
OAI21X1 OAI21X1_263 ( .A(_894_), .B(_895_), .C(vdd), .Y(_896_) );
NAND2X1 NAND2X1_264 ( .A(_896_), .B(_900_), .Y(csa_inst_rca0_1_fa0_o_sum) );
OAI21X1 OAI21X1_264 ( .A(_897_), .B(_894_), .C(_899_), .Y(csa_inst_rca0_1_fa0_o_carry) );
INVX1 INVX1_164 ( .A(csa_inst_rca0_1_fa0_o_carry), .Y(_904_) );
OR2X2 OR2X2_101 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_905_) );
NAND2X1 NAND2X1_265 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_906_) );
NAND3X1 NAND3X1_101 ( .A(_904_), .B(_906_), .C(_905_), .Y(_907_) );
NOR2X1 NOR2X1_101 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_901_) );
AND2X2 AND2X2_101 ( .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_902_) );
OAI21X1 OAI21X1_265 ( .A(_901_), .B(_902_), .C(csa_inst_rca0_1_fa0_o_carry), .Y(_903_) );
NAND2X1 NAND2X1_266 ( .A(_903_), .B(_907_), .Y(csa_inst_rca0_1_fa1_o_sum) );
OAI21X1 OAI21X1_266 ( .A(_904_), .B(_901_), .C(_906_), .Y(csa_inst_rca0_1_fa1_o_carry) );
INVX1 INVX1_165 ( .A(csa_inst_rca0_1_fa1_o_carry), .Y(_911_) );
OR2X2 OR2X2_102 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_912_) );
NAND2X1 NAND2X1_267 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_913_) );
NAND3X1 NAND3X1_102 ( .A(_911_), .B(_913_), .C(_912_), .Y(_914_) );
NOR2X1 NOR2X1_102 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_908_) );
AND2X2 AND2X2_102 ( .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_909_) );
OAI21X1 OAI21X1_267 ( .A(_908_), .B(_909_), .C(csa_inst_rca0_1_fa1_o_carry), .Y(_910_) );
NAND2X1 NAND2X1_268 ( .A(_910_), .B(_914_), .Y(csa_inst_rca0_1_fa2_o_sum) );
OAI21X1 OAI21X1_268 ( .A(_911_), .B(_908_), .C(_913_), .Y(csa_inst_cout0_1) );
INVX1 INVX1_166 ( .A(gnd), .Y(_918_) );
OR2X2 OR2X2_103 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_919_) );
NAND2X1 NAND2X1_269 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_920_) );
NAND3X1 NAND3X1_103 ( .A(_918_), .B(_920_), .C(_919_), .Y(_921_) );
NOR2X1 NOR2X1_103 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_915_) );
AND2X2 AND2X2_103 ( .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_916_) );
OAI21X1 OAI21X1_269 ( .A(_915_), .B(_916_), .C(gnd), .Y(_917_) );
NAND2X1 NAND2X1_270 ( .A(_917_), .B(_921_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_270 ( .A(_918_), .B(_915_), .C(_920_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_167 ( .A(rca_inst_fa3_i_carry), .Y(_925_) );
OR2X2 OR2X2_104 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_926_) );
NAND2X1 NAND2X1_271 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_927_) );
NAND3X1 NAND3X1_104 ( .A(_925_), .B(_927_), .C(_926_), .Y(_928_) );
NOR2X1 NOR2X1_104 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_922_) );
AND2X2 AND2X2_104 ( .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_923_) );
OAI21X1 OAI21X1_271 ( .A(_922_), .B(_923_), .C(rca_inst_fa3_i_carry), .Y(_924_) );
NAND2X1 NAND2X1_272 ( .A(_924_), .B(_928_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_272 ( .A(_925_), .B(_922_), .C(_927_), .Y(rca_inst_cout) );
INVX1 INVX1_168 ( .A(rca_inst_fa0_o_carry), .Y(_932_) );
OR2X2 OR2X2_105 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_933_) );
NAND2X1 NAND2X1_273 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_934_) );
NAND3X1 NAND3X1_105 ( .A(_932_), .B(_934_), .C(_933_), .Y(_935_) );
NOR2X1 NOR2X1_105 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_929_) );
AND2X2 AND2X2_105 ( .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_930_) );
OAI21X1 OAI21X1_273 ( .A(_929_), .B(_930_), .C(rca_inst_fa0_o_carry), .Y(_931_) );
NAND2X1 NAND2X1_274 ( .A(_931_), .B(_935_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_274 ( .A(_932_), .B(_929_), .C(_934_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_169 ( .A(rca_inst_fa_1__o_carry), .Y(_939_) );
OR2X2 OR2X2_106 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_940_) );
NAND2X1 NAND2X1_275 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_941_) );
NAND3X1 NAND3X1_106 ( .A(_939_), .B(_941_), .C(_940_), .Y(_942_) );
NOR2X1 NOR2X1_106 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_936_) );
AND2X2 AND2X2_106 ( .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_937_) );
OAI21X1 OAI21X1_275 ( .A(_936_), .B(_937_), .C(rca_inst_fa_1__o_carry), .Y(_938_) );
NAND2X1 NAND2X1_276 ( .A(_938_), .B(_942_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_276 ( .A(_939_), .B(_936_), .C(_941_), .Y(rca_inst_fa3_i_carry) );
BUFX2 BUFX2_1 ( .A(w_cout_13_), .Y(cout) );
BUFX2 BUFX2_2 ( .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .A(_0__54_), .Y(sum[54]) );
INVX1 INVX1_170 ( .A(_1_), .Y(_73_) );
BUFX2 BUFX2_57 ( .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_58 ( .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_59 ( .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_60 ( .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_61 ( .A(rca_inst_cout), .Y(w_cout_0_) );
BUFX2 BUFX2_62 ( .A(csa_inst_cin), .Y(w_cout_12_) );
endmodule
