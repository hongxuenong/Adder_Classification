module csa_59bit ( gnd, vdd, i_add_term1, i_add_term2, sum, cout);

input gnd, vdd;
output cout;
input [58:0] i_add_term1;
input [58:0] i_add_term2;
output [58:0] sum;

BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(w_cout_14_), .Y(cout) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_sum), .Y(sum[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_sum), .Y(sum[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_2__o_sum), .Y(sum[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_o_sum), .Y(sum[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_0__4_), .Y(sum[4]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_0__5_), .Y(sum[5]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_0__6_), .Y(sum[6]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_0__7_), .Y(sum[7]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_0__8_), .Y(sum[8]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_0__9_), .Y(sum[9]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_0__10_), .Y(sum[10]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_0__11_), .Y(sum[11]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_0__12_), .Y(sum[12]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_0__13_), .Y(sum[13]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_0__14_), .Y(sum[14]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_0__15_), .Y(sum[15]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_0__16_), .Y(sum[16]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_0__17_), .Y(sum[17]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_0__18_), .Y(sum[18]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_0__19_), .Y(sum[19]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_0__20_), .Y(sum[20]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_0__21_), .Y(sum[21]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_0__22_), .Y(sum[22]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_0__23_), .Y(sum[23]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_0__24_), .Y(sum[24]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_0__25_), .Y(sum[25]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_0__26_), .Y(sum[26]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_0__27_), .Y(sum[27]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_0__28_), .Y(sum[28]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_0__29_), .Y(sum[29]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_0__30_), .Y(sum[30]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_0__31_), .Y(sum[31]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_0__32_), .Y(sum[32]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_0__33_), .Y(sum[33]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_0__34_), .Y(sum[34]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_0__35_), .Y(sum[35]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_0__36_), .Y(sum[36]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_0__37_), .Y(sum[37]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_0__38_), .Y(sum[38]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_0__39_), .Y(sum[39]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_0__40_), .Y(sum[40]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_0__41_), .Y(sum[41]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_0__42_), .Y(sum[42]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_0__43_), .Y(sum[43]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_0__44_), .Y(sum[44]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_0__45_), .Y(sum[45]) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_0__46_), .Y(sum[46]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_0__47_), .Y(sum[47]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_0__48_), .Y(sum[48]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_0__49_), .Y(sum[49]) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_0__50_), .Y(sum[50]) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(_0__51_), .Y(sum[51]) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(_0__52_), .Y(sum[52]) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(_0__53_), .Y(sum[53]) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_0__54_), .Y(sum[54]) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_0__55_), .Y(sum[55]) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_0__56_), .Y(sum[56]) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_0__57_), .Y(sum[57]) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(_0__58_), .Y(sum[58]) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_79_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(rca_inst_cout), .Y(_80_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_79_), .C(_80_), .Y(w_cout_1_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_3__0_), .Y(_81_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_4__0_), .B(rca_inst_cout), .Y(_82_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_81_), .C(_82_), .Y(_0__4_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_3__1_), .Y(_83_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_4__1_), .Y(_84_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_83_), .C(_84_), .Y(_0__5_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_3__2_), .Y(_85_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_4__2_), .Y(_86_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_85_), .C(_86_), .Y(_0__6_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_3__3_), .Y(_87_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_4__3_), .Y(_88_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .B(_87_), .C(_88_), .Y(_0__7_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_92_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_93_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_94_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_94_), .C(_93_), .Y(_95_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_89_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_90_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_90_), .C(gnd), .Y(_91_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_95_), .Y(_3__0_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_89_), .C(_94_), .Y(_5__1_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_5__3_), .Y(_99_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_100_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_101_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_101_), .C(_100_), .Y(_102_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_96_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_97_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_97_), .C(_5__3_), .Y(_98_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_102_), .Y(_3__3_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_96_), .C(_101_), .Y(_1_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_5__1_), .Y(_106_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_107_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_108_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_106_), .B(_108_), .C(_107_), .Y(_109_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_103_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_104_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_104_), .C(_5__1_), .Y(_105_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_109_), .Y(_3__1_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_106_), .B(_103_), .C(_108_), .Y(_5__2_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_5__2_), .Y(_113_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_114_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_115_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_115_), .C(_114_), .Y(_116_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_110_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_111_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_111_), .C(_5__2_), .Y(_112_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_116_), .Y(_3__2_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_110_), .C(_115_), .Y(_5__3_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_120_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_121_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_122_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_122_), .C(_121_), .Y(_123_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_117_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[4]), .B(i_add_term1[4]), .Y(_118_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_118_), .C(vdd), .Y(_119_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_123_), .Y(_4__0_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_117_), .C(_122_), .Y(_6__1_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_6__3_), .Y(_127_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_128_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_129_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_129_), .C(_128_), .Y(_130_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_124_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[7]), .B(i_add_term1[7]), .Y(_125_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_125_), .C(_6__3_), .Y(_126_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_130_), .Y(_4__3_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_124_), .C(_129_), .Y(_2_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_6__1_), .Y(_134_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_135_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_136_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_136_), .C(_135_), .Y(_137_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_131_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[5]), .B(i_add_term1[5]), .Y(_132_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_132_), .C(_6__1_), .Y(_133_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_137_), .Y(_4__1_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_131_), .C(_136_), .Y(_6__2_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_6__2_), .Y(_141_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_142_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_143_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_143_), .C(_142_), .Y(_144_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_138_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[6]), .B(i_add_term1[6]), .Y(_139_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_139_), .C(_6__2_), .Y(_140_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_144_), .Y(_4__2_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_138_), .C(_143_), .Y(_6__3_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_145_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(w_cout_1_), .Y(_146_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_145_), .C(_146_), .Y(w_cout_2_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_9__0_), .Y(_147_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_10__0_), .B(w_cout_1_), .Y(_148_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_147_), .C(_148_), .Y(_0__8_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_9__1_), .Y(_149_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_10__1_), .Y(_150_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_149_), .C(_150_), .Y(_0__9_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_9__2_), .Y(_151_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_10__2_), .Y(_152_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_151_), .C(_152_), .Y(_0__10_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_9__3_), .Y(_153_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_10__3_), .Y(_154_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(w_cout_1_), .B(_153_), .C(_154_), .Y(_0__11_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_158_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_159_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_160_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_160_), .C(_159_), .Y(_161_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_155_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_156_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_156_), .C(gnd), .Y(_157_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_161_), .Y(_9__0_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_155_), .C(_160_), .Y(_11__1_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_11__3_), .Y(_165_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_166_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_167_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_167_), .C(_166_), .Y(_168_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_162_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_163_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_163_), .C(_11__3_), .Y(_164_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_168_), .Y(_9__3_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_162_), .C(_167_), .Y(_7_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_11__1_), .Y(_172_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_173_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_174_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_174_), .C(_173_), .Y(_175_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_169_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_170_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_170_), .C(_11__1_), .Y(_171_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_175_), .Y(_9__1_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_169_), .C(_174_), .Y(_11__2_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_11__2_), .Y(_179_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_180_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_181_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_181_), .C(_180_), .Y(_182_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_176_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_177_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_177_), .C(_11__2_), .Y(_178_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_182_), .Y(_9__2_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_176_), .C(_181_), .Y(_11__3_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_186_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_187_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_188_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_188_), .C(_187_), .Y(_189_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_183_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[8]), .B(i_add_term1[8]), .Y(_184_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_184_), .C(vdd), .Y(_185_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_189_), .Y(_10__0_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_183_), .C(_188_), .Y(_12__1_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_12__3_), .Y(_193_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_194_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_195_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_195_), .C(_194_), .Y(_196_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_190_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[11]), .B(i_add_term1[11]), .Y(_191_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_191_), .C(_12__3_), .Y(_192_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(_196_), .Y(_10__3_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_190_), .C(_195_), .Y(_8_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_12__1_), .Y(_200_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_201_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_202_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_202_), .C(_201_), .Y(_203_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_197_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[9]), .B(i_add_term1[9]), .Y(_198_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_198_), .C(_12__1_), .Y(_199_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_203_), .Y(_10__1_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_197_), .C(_202_), .Y(_12__2_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_12__2_), .Y(_207_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_208_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_209_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_209_), .C(_208_), .Y(_210_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_204_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[10]), .B(i_add_term1[10]), .Y(_205_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_205_), .C(_12__2_), .Y(_206_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_210_), .Y(_10__2_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_204_), .C(_209_), .Y(_12__3_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_211_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(w_cout_2_), .Y(_212_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_211_), .C(_212_), .Y(w_cout_3_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_15__0_), .Y(_213_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_16__0_), .B(w_cout_2_), .Y(_214_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_213_), .C(_214_), .Y(_0__12_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_15__1_), .Y(_215_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_16__1_), .Y(_216_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_215_), .C(_216_), .Y(_0__13_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_15__2_), .Y(_217_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_16__2_), .Y(_218_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_217_), .C(_218_), .Y(_0__14_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_15__3_), .Y(_219_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_16__3_), .Y(_220_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(w_cout_2_), .B(_219_), .C(_220_), .Y(_0__15_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_224_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_225_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_226_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_226_), .C(_225_), .Y(_227_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_221_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_222_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_222_), .C(gnd), .Y(_223_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_227_), .Y(_15__0_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_221_), .C(_226_), .Y(_17__1_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_17__3_), .Y(_231_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_232_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_233_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_233_), .C(_232_), .Y(_234_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_228_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_229_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_229_), .C(_17__3_), .Y(_230_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_234_), .Y(_15__3_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_228_), .C(_233_), .Y(_13_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_17__1_), .Y(_238_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_239_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_240_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_238_), .B(_240_), .C(_239_), .Y(_241_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_235_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_236_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_236_), .C(_17__1_), .Y(_237_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_241_), .Y(_15__1_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_238_), .B(_235_), .C(_240_), .Y(_17__2_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_17__2_), .Y(_245_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_246_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_247_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_247_), .C(_246_), .Y(_248_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_242_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_243_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_243_), .C(_17__2_), .Y(_244_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_248_), .Y(_15__2_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_242_), .C(_247_), .Y(_17__3_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_252_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_253_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_254_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_254_), .C(_253_), .Y(_255_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_249_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[12]), .B(i_add_term1[12]), .Y(_250_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_250_), .C(vdd), .Y(_251_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_255_), .Y(_16__0_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_249_), .C(_254_), .Y(_18__1_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_18__3_), .Y(_259_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_260_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_261_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_261_), .C(_260_), .Y(_262_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_256_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[15]), .B(i_add_term1[15]), .Y(_257_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_257_), .C(_18__3_), .Y(_258_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_262_), .Y(_16__3_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_256_), .C(_261_), .Y(_14_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_18__1_), .Y(_266_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_267_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_268_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_268_), .C(_267_), .Y(_269_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_263_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[13]), .B(i_add_term1[13]), .Y(_264_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_264_), .C(_18__1_), .Y(_265_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_269_), .Y(_16__1_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_263_), .C(_268_), .Y(_18__2_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_18__2_), .Y(_273_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_274_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_275_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_275_), .C(_274_), .Y(_276_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_270_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[14]), .B(i_add_term1[14]), .Y(_271_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_271_), .C(_18__2_), .Y(_272_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_276_), .Y(_16__2_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_270_), .C(_275_), .Y(_18__3_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_277_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(w_cout_3_), .Y(_278_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_277_), .C(_278_), .Y(w_cout_4_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_21__0_), .Y(_279_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_22__0_), .B(w_cout_3_), .Y(_280_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_279_), .C(_280_), .Y(_0__16_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_21__1_), .Y(_281_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_22__1_), .Y(_282_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_281_), .C(_282_), .Y(_0__17_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_21__2_), .Y(_283_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_22__2_), .Y(_284_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_283_), .C(_284_), .Y(_0__18_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_21__3_), .Y(_285_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_22__3_), .Y(_286_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(w_cout_3_), .B(_285_), .C(_286_), .Y(_0__19_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_290_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_291_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_292_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_292_), .C(_291_), .Y(_293_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_287_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_288_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_287_), .B(_288_), .C(gnd), .Y(_289_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_293_), .Y(_21__0_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_287_), .C(_292_), .Y(_23__1_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_23__3_), .Y(_297_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_298_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_299_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_299_), .C(_298_), .Y(_300_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_294_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_295_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_295_), .C(_23__3_), .Y(_296_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_300_), .Y(_21__3_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_294_), .C(_299_), .Y(_19_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_23__1_), .Y(_304_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_305_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_306_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_306_), .C(_305_), .Y(_307_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_301_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_302_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_302_), .C(_23__1_), .Y(_303_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_307_), .Y(_21__1_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_301_), .C(_306_), .Y(_23__2_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_23__2_), .Y(_311_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_312_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_313_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_313_), .C(_312_), .Y(_314_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_308_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_309_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_309_), .C(_23__2_), .Y(_310_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_314_), .Y(_21__2_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_308_), .C(_313_), .Y(_23__3_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_318_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_319_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_320_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_320_), .C(_319_), .Y(_321_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_315_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[16]), .B(i_add_term1[16]), .Y(_316_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_316_), .C(vdd), .Y(_317_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_321_), .Y(_22__0_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_315_), .C(_320_), .Y(_24__1_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_24__3_), .Y(_325_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_326_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_327_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_327_), .C(_326_), .Y(_328_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_322_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[19]), .B(i_add_term1[19]), .Y(_323_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_323_), .C(_24__3_), .Y(_324_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_328_), .Y(_22__3_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_322_), .C(_327_), .Y(_20_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_24__1_), .Y(_332_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_333_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_334_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_334_), .C(_333_), .Y(_335_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_329_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[17]), .B(i_add_term1[17]), .Y(_330_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_330_), .C(_24__1_), .Y(_331_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_335_), .Y(_22__1_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_329_), .C(_334_), .Y(_24__2_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_24__2_), .Y(_339_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_340_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_341_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_341_), .C(_340_), .Y(_342_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_336_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[18]), .B(i_add_term1[18]), .Y(_337_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_337_), .C(_24__2_), .Y(_338_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_342_), .Y(_22__2_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_336_), .C(_341_), .Y(_24__3_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(_343_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(w_cout_4_), .Y(_344_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_343_), .C(_344_), .Y(w_cout_5_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_27__0_), .Y(_345_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_28__0_), .B(w_cout_4_), .Y(_346_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_345_), .C(_346_), .Y(_0__20_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_27__1_), .Y(_347_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_28__1_), .Y(_348_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_347_), .C(_348_), .Y(_0__21_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_27__2_), .Y(_349_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_28__2_), .Y(_350_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_349_), .C(_350_), .Y(_0__22_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_27__3_), .Y(_351_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_28__3_), .Y(_352_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(w_cout_4_), .B(_351_), .C(_352_), .Y(_0__23_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_356_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_357_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_358_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_358_), .C(_357_), .Y(_359_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_353_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_354_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_354_), .C(gnd), .Y(_355_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_359_), .Y(_27__0_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_353_), .C(_358_), .Y(_29__1_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_29__3_), .Y(_363_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_364_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_365_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_365_), .C(_364_), .Y(_366_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_360_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_361_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_361_), .C(_29__3_), .Y(_362_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_366_), .Y(_27__3_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_360_), .C(_365_), .Y(_25_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_29__1_), .Y(_370_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_371_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_372_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_372_), .C(_371_), .Y(_373_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_367_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_368_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_368_), .C(_29__1_), .Y(_369_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_373_), .Y(_27__1_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_367_), .C(_372_), .Y(_29__2_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_29__2_), .Y(_377_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_378_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_379_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_379_), .C(_378_), .Y(_380_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_374_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_375_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_375_), .C(_29__2_), .Y(_376_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_380_), .Y(_27__2_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_374_), .C(_379_), .Y(_29__3_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_384_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_385_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_386_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_386_), .C(_385_), .Y(_387_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_381_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[20]), .B(i_add_term1[20]), .Y(_382_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_382_), .C(vdd), .Y(_383_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_387_), .Y(_28__0_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_381_), .C(_386_), .Y(_30__1_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_30__3_), .Y(_391_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_392_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_393_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_393_), .C(_392_), .Y(_394_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_388_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[23]), .B(i_add_term1[23]), .Y(_389_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(_389_), .C(_30__3_), .Y(_390_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_394_), .Y(_28__3_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_388_), .C(_393_), .Y(_26_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_30__1_), .Y(_398_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_399_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_400_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_400_), .C(_399_), .Y(_401_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_395_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[21]), .B(i_add_term1[21]), .Y(_396_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_396_), .C(_30__1_), .Y(_397_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_401_), .Y(_28__1_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_395_), .C(_400_), .Y(_30__2_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_30__2_), .Y(_405_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_406_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_407_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_407_), .C(_406_), .Y(_408_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_402_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[22]), .B(i_add_term1[22]), .Y(_403_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_403_), .C(_30__2_), .Y(_404_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_408_), .Y(_28__2_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_402_), .C(_407_), .Y(_30__3_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_31_), .Y(_409_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(w_cout_5_), .Y(_410_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_409_), .C(_410_), .Y(w_cout_6_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_33__0_), .Y(_411_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_34__0_), .B(w_cout_5_), .Y(_412_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_411_), .C(_412_), .Y(_0__24_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_33__1_), .Y(_413_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_34__1_), .Y(_414_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_413_), .C(_414_), .Y(_0__25_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_33__2_), .Y(_415_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_34__2_), .Y(_416_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_415_), .C(_416_), .Y(_0__26_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_33__3_), .Y(_417_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_34__3_), .Y(_418_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(w_cout_5_), .B(_417_), .C(_418_), .Y(_0__27_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_422_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_423_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_424_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_422_), .B(_424_), .C(_423_), .Y(_425_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_419_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_420_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_420_), .C(gnd), .Y(_421_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_425_), .Y(_33__0_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_422_), .B(_419_), .C(_424_), .Y(_35__1_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_35__3_), .Y(_429_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_430_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_431_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(_431_), .C(_430_), .Y(_432_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_426_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_427_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_427_), .C(_35__3_), .Y(_428_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_432_), .Y(_33__3_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(_426_), .C(_431_), .Y(_31_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(_35__1_), .Y(_436_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_437_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_438_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_438_), .C(_437_), .Y(_439_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_433_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_434_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_434_), .C(_35__1_), .Y(_435_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_439_), .Y(_33__1_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_436_), .B(_433_), .C(_438_), .Y(_35__2_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_35__2_), .Y(_443_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_444_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_445_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_445_), .C(_444_), .Y(_446_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_440_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_441_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_441_), .C(_35__2_), .Y(_442_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_446_), .Y(_33__2_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_440_), .C(_445_), .Y(_35__3_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_450_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_451_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_452_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_452_), .C(_451_), .Y(_453_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_447_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[24]), .B(i_add_term1[24]), .Y(_448_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_448_), .C(vdd), .Y(_449_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_453_), .Y(_34__0_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_447_), .C(_452_), .Y(_36__1_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_36__3_), .Y(_457_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_458_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_459_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_459_), .C(_458_), .Y(_460_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_454_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[27]), .B(i_add_term1[27]), .Y(_455_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_454_), .B(_455_), .C(_36__3_), .Y(_456_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_456_), .B(_460_), .Y(_34__3_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_454_), .C(_459_), .Y(_32_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_36__1_), .Y(_464_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_465_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_466_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_466_), .C(_465_), .Y(_467_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_461_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[25]), .B(i_add_term1[25]), .Y(_462_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_462_), .C(_36__1_), .Y(_463_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_467_), .Y(_34__1_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_461_), .C(_466_), .Y(_36__2_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_36__2_), .Y(_471_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_472_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_473_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_473_), .C(_472_), .Y(_474_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_468_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[26]), .B(i_add_term1[26]), .Y(_469_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_468_), .B(_469_), .C(_36__2_), .Y(_470_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_470_), .B(_474_), .Y(_34__2_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_468_), .C(_473_), .Y(_36__3_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(_37_), .Y(_475_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(w_cout_6_), .Y(_476_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_475_), .C(_476_), .Y(w_cout_7_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_39__0_), .Y(_477_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_40__0_), .B(w_cout_6_), .Y(_478_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_477_), .C(_478_), .Y(_0__28_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_39__1_), .Y(_479_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_40__1_), .Y(_480_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_479_), .C(_480_), .Y(_0__29_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_39__2_), .Y(_481_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_40__2_), .Y(_482_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_481_), .C(_482_), .Y(_0__30_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_39__3_), .Y(_483_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_40__3_), .Y(_484_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(w_cout_6_), .B(_483_), .C(_484_), .Y(_0__31_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_488_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_489_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_490_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_490_), .C(_489_), .Y(_491_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_485_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_486_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_486_), .C(gnd), .Y(_487_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_491_), .Y(_39__0_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_485_), .C(_490_), .Y(_41__1_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_41__3_), .Y(_495_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_496_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_497_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_495_), .B(_497_), .C(_496_), .Y(_498_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_492_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_493_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_492_), .B(_493_), .C(_41__3_), .Y(_494_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_498_), .Y(_39__3_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_495_), .B(_492_), .C(_497_), .Y(_37_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_41__1_), .Y(_502_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_503_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_504_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_502_), .B(_504_), .C(_503_), .Y(_505_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_499_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_500_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_500_), .C(_41__1_), .Y(_501_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_501_), .B(_505_), .Y(_39__1_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_502_), .B(_499_), .C(_504_), .Y(_41__2_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(_41__2_), .Y(_509_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_510_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_511_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_511_), .C(_510_), .Y(_512_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_506_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_507_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_507_), .C(_41__2_), .Y(_508_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_512_), .Y(_39__2_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_506_), .C(_511_), .Y(_41__3_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_516_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_517_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_518_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_518_), .C(_517_), .Y(_519_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_513_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[28]), .B(i_add_term1[28]), .Y(_514_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_514_), .C(vdd), .Y(_515_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_515_), .B(_519_), .Y(_40__0_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_513_), .C(_518_), .Y(_42__1_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(_42__3_), .Y(_523_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_524_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_525_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_525_), .C(_524_), .Y(_526_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_520_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[31]), .B(i_add_term1[31]), .Y(_521_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_521_), .C(_42__3_), .Y(_522_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_522_), .B(_526_), .Y(_40__3_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_520_), .C(_525_), .Y(_38_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_42__1_), .Y(_530_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_531_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_532_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_532_), .C(_531_), .Y(_533_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_527_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[29]), .B(i_add_term1[29]), .Y(_528_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_528_), .C(_42__1_), .Y(_529_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_533_), .Y(_40__1_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_527_), .C(_532_), .Y(_42__2_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(_42__2_), .Y(_537_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_538_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_539_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_539_), .C(_538_), .Y(_540_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_534_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[30]), .B(i_add_term1[30]), .Y(_535_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_535_), .C(_42__2_), .Y(_536_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_536_), .B(_540_), .Y(_40__2_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_534_), .C(_539_), .Y(_42__3_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(_541_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(w_cout_7_), .Y(_542_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_541_), .C(_542_), .Y(w_cout_8_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(_45__0_), .Y(_543_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_46__0_), .B(w_cout_7_), .Y(_544_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_543_), .C(_544_), .Y(_0__32_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_45__1_), .Y(_545_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_46__1_), .Y(_546_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_545_), .C(_546_), .Y(_0__33_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_45__2_), .Y(_547_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_46__2_), .Y(_548_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_547_), .C(_548_), .Y(_0__34_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(_45__3_), .Y(_549_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_46__3_), .Y(_550_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(w_cout_7_), .B(_549_), .C(_550_), .Y(_0__35_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_554_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_555_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_556_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_556_), .C(_555_), .Y(_557_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_551_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_552_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_551_), .B(_552_), .C(gnd), .Y(_553_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_553_), .B(_557_), .Y(_45__0_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_551_), .C(_556_), .Y(_47__1_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(_47__3_), .Y(_561_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_562_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_563_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_563_), .C(_562_), .Y(_564_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_558_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_559_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_559_), .C(_47__3_), .Y(_560_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_560_), .B(_564_), .Y(_45__3_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_558_), .C(_563_), .Y(_43_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(_47__1_), .Y(_568_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_569_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_570_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_570_), .C(_569_), .Y(_571_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_565_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_566_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_566_), .C(_47__1_), .Y(_567_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_567_), .B(_571_), .Y(_45__1_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_565_), .C(_570_), .Y(_47__2_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(_47__2_), .Y(_575_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_576_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_577_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_577_), .C(_576_), .Y(_578_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_572_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_573_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_572_), .B(_573_), .C(_47__2_), .Y(_574_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_574_), .B(_578_), .Y(_45__2_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_572_), .C(_577_), .Y(_47__3_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_582_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_583_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_584_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_584_), .C(_583_), .Y(_585_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_579_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[32]), .B(i_add_term1[32]), .Y(_580_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_579_), .B(_580_), .C(vdd), .Y(_581_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_581_), .B(_585_), .Y(_46__0_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_579_), .C(_584_), .Y(_48__1_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(_48__3_), .Y(_589_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_590_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_591_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_589_), .B(_591_), .C(_590_), .Y(_592_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_586_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[35]), .B(i_add_term1[35]), .Y(_587_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_586_), .B(_587_), .C(_48__3_), .Y(_588_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_588_), .B(_592_), .Y(_46__3_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_589_), .B(_586_), .C(_591_), .Y(_44_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_48__1_), .Y(_596_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_597_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_598_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_598_), .C(_597_), .Y(_599_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_593_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[33]), .B(i_add_term1[33]), .Y(_594_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_594_), .C(_48__1_), .Y(_595_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_595_), .B(_599_), .Y(_46__1_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_593_), .C(_598_), .Y(_48__2_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(_48__2_), .Y(_603_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_604_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_605_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_603_), .B(_605_), .C(_604_), .Y(_606_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_600_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[34]), .B(i_add_term1[34]), .Y(_601_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_601_), .C(_48__2_), .Y(_602_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_602_), .B(_606_), .Y(_46__2_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_603_), .B(_600_), .C(_605_), .Y(_48__3_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_49_), .Y(_607_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(w_cout_8_), .Y(_608_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_607_), .C(_608_), .Y(w_cout_9_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_51__0_), .Y(_609_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_52__0_), .B(w_cout_8_), .Y(_610_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_609_), .C(_610_), .Y(_0__36_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_51__1_), .Y(_611_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_52__1_), .Y(_612_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_611_), .C(_612_), .Y(_0__37_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_51__2_), .Y(_613_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_52__2_), .Y(_614_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_613_), .C(_614_), .Y(_0__38_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_51__3_), .Y(_615_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_52__3_), .Y(_616_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(w_cout_8_), .B(_615_), .C(_616_), .Y(_0__39_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_620_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_621_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_622_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_622_), .C(_621_), .Y(_623_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_617_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_618_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_617_), .B(_618_), .C(gnd), .Y(_619_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_623_), .Y(_51__0_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_620_), .B(_617_), .C(_622_), .Y(_53__1_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_53__3_), .Y(_627_) );
OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_628_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_629_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(_629_), .C(_628_), .Y(_630_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_624_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_625_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_624_), .B(_625_), .C(_53__3_), .Y(_626_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_630_), .Y(_51__3_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(_624_), .C(_629_), .Y(_49_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(_53__1_), .Y(_634_) );
OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_635_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_636_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_634_), .B(_636_), .C(_635_), .Y(_637_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_631_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_632_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_631_), .B(_632_), .C(_53__1_), .Y(_633_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_637_), .Y(_51__1_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_634_), .B(_631_), .C(_636_), .Y(_53__2_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(_53__2_), .Y(_641_) );
OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_642_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_643_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_641_), .B(_643_), .C(_642_), .Y(_644_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_638_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_639_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_639_), .C(_53__2_), .Y(_640_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(_644_), .Y(_51__2_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_641_), .B(_638_), .C(_643_), .Y(_53__3_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_648_) );
OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_649_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_650_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_650_), .C(_649_), .Y(_651_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_645_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[36]), .B(i_add_term1[36]), .Y(_646_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_645_), .B(_646_), .C(vdd), .Y(_647_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_647_), .B(_651_), .Y(_52__0_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_648_), .B(_645_), .C(_650_), .Y(_54__1_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(_54__3_), .Y(_655_) );
OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_656_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_657_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_657_), .C(_656_), .Y(_658_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_652_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[39]), .B(i_add_term1[39]), .Y(_653_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_653_), .C(_54__3_), .Y(_654_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_654_), .B(_658_), .Y(_52__3_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_652_), .C(_657_), .Y(_50_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(_54__1_), .Y(_662_) );
OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_663_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_664_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_664_), .C(_663_), .Y(_665_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_659_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[37]), .B(i_add_term1[37]), .Y(_660_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_659_), .B(_660_), .C(_54__1_), .Y(_661_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_661_), .B(_665_), .Y(_52__1_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_659_), .C(_664_), .Y(_54__2_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(_54__2_), .Y(_669_) );
OR2X2 OR2X2_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_670_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_671_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_669_), .B(_671_), .C(_670_), .Y(_672_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_666_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[38]), .B(i_add_term1[38]), .Y(_667_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_666_), .B(_667_), .C(_54__2_), .Y(_668_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_672_), .Y(_52__2_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_669_), .B(_666_), .C(_671_), .Y(_54__3_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(_55_), .Y(_673_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(w_cout_9_), .Y(_674_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_673_), .C(_674_), .Y(w_cout_10_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(_57__0_), .Y(_675_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_58__0_), .B(w_cout_9_), .Y(_676_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_675_), .C(_676_), .Y(_0__40_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(_57__1_), .Y(_677_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_58__1_), .Y(_678_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_677_), .C(_678_), .Y(_0__41_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(_57__2_), .Y(_679_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_58__2_), .Y(_680_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_679_), .C(_680_), .Y(_0__42_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(_57__3_), .Y(_681_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_58__3_), .Y(_682_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(w_cout_9_), .B(_681_), .C(_682_), .Y(_0__43_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_686_) );
OR2X2 OR2X2_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_687_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_688_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_686_), .B(_688_), .C(_687_), .Y(_689_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_683_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_684_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_683_), .B(_684_), .C(gnd), .Y(_685_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_689_), .Y(_57__0_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_686_), .B(_683_), .C(_688_), .Y(_59__1_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(_59__3_), .Y(_693_) );
OR2X2 OR2X2_74 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_694_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_695_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_695_), .C(_694_), .Y(_696_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_690_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_691_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_690_), .B(_691_), .C(_59__3_), .Y(_692_) );
NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_692_), .B(_696_), .Y(_57__3_) );
OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_690_), .C(_695_), .Y(_55_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(_59__1_), .Y(_700_) );
OR2X2 OR2X2_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_701_) );
NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_702_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_700_), .B(_702_), .C(_701_), .Y(_703_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_697_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_698_) );
OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_697_), .B(_698_), .C(_59__1_), .Y(_699_) );
NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_703_), .Y(_57__1_) );
OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_700_), .B(_697_), .C(_702_), .Y(_59__2_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(_59__2_), .Y(_707_) );
OR2X2 OR2X2_76 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_708_) );
NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_709_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_707_), .B(_709_), .C(_708_), .Y(_710_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_704_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_705_) );
OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_705_), .C(_59__2_), .Y(_706_) );
NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_710_), .Y(_57__2_) );
OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_707_), .B(_704_), .C(_709_), .Y(_59__3_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_714_) );
OR2X2 OR2X2_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_715_) );
NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_716_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_714_), .B(_716_), .C(_715_), .Y(_717_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_711_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[40]), .B(i_add_term1[40]), .Y(_712_) );
OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_712_), .C(vdd), .Y(_713_) );
NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_717_), .Y(_58__0_) );
OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_714_), .B(_711_), .C(_716_), .Y(_60__1_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(_60__3_), .Y(_721_) );
OR2X2 OR2X2_78 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_722_) );
NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_723_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_721_), .B(_723_), .C(_722_), .Y(_724_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_718_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[43]), .B(i_add_term1[43]), .Y(_719_) );
OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_718_), .B(_719_), .C(_60__3_), .Y(_720_) );
NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_720_), .B(_724_), .Y(_58__3_) );
OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_721_), .B(_718_), .C(_723_), .Y(_56_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(_60__1_), .Y(_728_) );
OR2X2 OR2X2_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_729_) );
NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_730_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_728_), .B(_730_), .C(_729_), .Y(_731_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_725_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[41]), .B(i_add_term1[41]), .Y(_726_) );
OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(_726_), .C(_60__1_), .Y(_727_) );
NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_727_), .B(_731_), .Y(_58__1_) );
OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_728_), .B(_725_), .C(_730_), .Y(_60__2_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(_60__2_), .Y(_735_) );
OR2X2 OR2X2_80 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_736_) );
NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_737_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_735_), .B(_737_), .C(_736_), .Y(_738_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_732_) );
AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[42]), .B(i_add_term1[42]), .Y(_733_) );
OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_733_), .C(_60__2_), .Y(_734_) );
NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_734_), .B(_738_), .Y(_58__2_) );
OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_735_), .B(_732_), .C(_737_), .Y(_60__3_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(_61_), .Y(_739_) );
NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(w_cout_10_), .Y(_740_) );
OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_739_), .C(_740_), .Y(w_cout_11_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(_63__0_), .Y(_741_) );
NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_64__0_), .B(w_cout_10_), .Y(_742_) );
OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_741_), .C(_742_), .Y(_0__44_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(_63__1_), .Y(_743_) );
NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_64__1_), .Y(_744_) );
OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_743_), .C(_744_), .Y(_0__45_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(_63__2_), .Y(_745_) );
NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_64__2_), .Y(_746_) );
OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_745_), .C(_746_), .Y(_0__46_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(_63__3_), .Y(_747_) );
NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_64__3_), .Y(_748_) );
OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(w_cout_10_), .B(_747_), .C(_748_), .Y(_0__47_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_752_) );
OR2X2 OR2X2_81 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_753_) );
NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_754_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(_754_), .C(_753_), .Y(_755_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_749_) );
AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_750_) );
OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(_750_), .C(gnd), .Y(_751_) );
NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_751_), .B(_755_), .Y(_63__0_) );
OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(_749_), .C(_754_), .Y(_65__1_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(_65__3_), .Y(_759_) );
OR2X2 OR2X2_82 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_760_) );
NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_761_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_759_), .B(_761_), .C(_760_), .Y(_762_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_756_) );
AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_757_) );
OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_756_), .B(_757_), .C(_65__3_), .Y(_758_) );
NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_758_), .B(_762_), .Y(_63__3_) );
OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_759_), .B(_756_), .C(_761_), .Y(_61_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(_65__1_), .Y(_766_) );
OR2X2 OR2X2_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_767_) );
NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_768_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_766_), .B(_768_), .C(_767_), .Y(_769_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_763_) );
AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_764_) );
OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_763_), .B(_764_), .C(_65__1_), .Y(_765_) );
NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_765_), .B(_769_), .Y(_63__1_) );
OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_766_), .B(_763_), .C(_768_), .Y(_65__2_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(_65__2_), .Y(_773_) );
OR2X2 OR2X2_84 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_774_) );
NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_775_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_775_), .C(_774_), .Y(_776_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_770_) );
AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_771_) );
OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_770_), .B(_771_), .C(_65__2_), .Y(_772_) );
NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_772_), .B(_776_), .Y(_63__2_) );
OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_770_), .C(_775_), .Y(_65__3_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_780_) );
OR2X2 OR2X2_85 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_781_) );
NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_782_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_780_), .B(_782_), .C(_781_), .Y(_783_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_777_) );
AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[44]), .B(i_add_term1[44]), .Y(_778_) );
OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_777_), .B(_778_), .C(vdd), .Y(_779_) );
NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_779_), .B(_783_), .Y(_64__0_) );
OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_780_), .B(_777_), .C(_782_), .Y(_66__1_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(_66__3_), .Y(_787_) );
OR2X2 OR2X2_86 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_788_) );
NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_789_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_789_), .C(_788_), .Y(_790_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_784_) );
AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[47]), .B(i_add_term1[47]), .Y(_785_) );
OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_784_), .B(_785_), .C(_66__3_), .Y(_786_) );
NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(_790_), .Y(_64__3_) );
OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_784_), .C(_789_), .Y(_62_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(_66__1_), .Y(_794_) );
OR2X2 OR2X2_87 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_795_) );
NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_796_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_796_), .C(_795_), .Y(_797_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_791_) );
AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[45]), .B(i_add_term1[45]), .Y(_792_) );
OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_791_), .B(_792_), .C(_66__1_), .Y(_793_) );
NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(_797_), .Y(_64__1_) );
OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_791_), .C(_796_), .Y(_66__2_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(_66__2_), .Y(_801_) );
OR2X2 OR2X2_88 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_802_) );
NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_803_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_801_), .B(_803_), .C(_802_), .Y(_804_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_798_) );
AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[46]), .B(i_add_term1[46]), .Y(_799_) );
OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_798_), .B(_799_), .C(_66__2_), .Y(_800_) );
NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_800_), .B(_804_), .Y(_64__2_) );
OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_801_), .B(_798_), .C(_803_), .Y(_66__3_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(_67_), .Y(_805_) );
NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(w_cout_11_), .Y(_806_) );
OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_805_), .C(_806_), .Y(w_cout_12_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(_69__0_), .Y(_807_) );
NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_70__0_), .B(w_cout_11_), .Y(_808_) );
OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_807_), .C(_808_), .Y(_0__48_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(_69__1_), .Y(_809_) );
NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_70__1_), .Y(_810_) );
OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_809_), .C(_810_), .Y(_0__49_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(_69__2_), .Y(_811_) );
NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_70__2_), .Y(_812_) );
OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_811_), .C(_812_), .Y(_0__50_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(_69__3_), .Y(_813_) );
NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_70__3_), .Y(_814_) );
OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(w_cout_11_), .B(_813_), .C(_814_), .Y(_0__51_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_818_) );
OR2X2 OR2X2_89 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_819_) );
NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_820_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_820_), .C(_819_), .Y(_821_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_815_) );
AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_816_) );
OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_815_), .B(_816_), .C(gnd), .Y(_817_) );
NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_817_), .B(_821_), .Y(_69__0_) );
OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_815_), .C(_820_), .Y(_71__1_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(_71__3_), .Y(_825_) );
OR2X2 OR2X2_90 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_826_) );
NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_827_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_825_), .B(_827_), .C(_826_), .Y(_828_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_822_) );
AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_823_) );
OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_822_), .B(_823_), .C(_71__3_), .Y(_824_) );
NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_824_), .B(_828_), .Y(_69__3_) );
OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_825_), .B(_822_), .C(_827_), .Y(_67_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(_71__1_), .Y(_832_) );
OR2X2 OR2X2_91 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_833_) );
NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_834_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_832_), .B(_834_), .C(_833_), .Y(_835_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_829_) );
AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_830_) );
OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_829_), .B(_830_), .C(_71__1_), .Y(_831_) );
NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_831_), .B(_835_), .Y(_69__1_) );
OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_832_), .B(_829_), .C(_834_), .Y(_71__2_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(_71__2_), .Y(_839_) );
OR2X2 OR2X2_92 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_840_) );
NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_841_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(_841_), .C(_840_), .Y(_842_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_836_) );
AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_837_) );
OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_836_), .B(_837_), .C(_71__2_), .Y(_838_) );
NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_838_), .B(_842_), .Y(_69__2_) );
OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(_836_), .C(_841_), .Y(_71__3_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_846_) );
OR2X2 OR2X2_93 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_847_) );
NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_848_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_848_), .C(_847_), .Y(_849_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_843_) );
AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[48]), .B(i_add_term1[48]), .Y(_844_) );
OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_844_), .C(vdd), .Y(_845_) );
NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_845_), .B(_849_), .Y(_70__0_) );
OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_843_), .C(_848_), .Y(_72__1_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(_72__3_), .Y(_853_) );
OR2X2 OR2X2_94 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_854_) );
NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_855_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_853_), .B(_855_), .C(_854_), .Y(_856_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_850_) );
AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[51]), .B(i_add_term1[51]), .Y(_851_) );
OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_850_), .B(_851_), .C(_72__3_), .Y(_852_) );
NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_852_), .B(_856_), .Y(_70__3_) );
OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_853_), .B(_850_), .C(_855_), .Y(_68_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(_72__1_), .Y(_860_) );
OR2X2 OR2X2_95 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_861_) );
NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_862_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_860_), .B(_862_), .C(_861_), .Y(_863_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_857_) );
AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[49]), .B(i_add_term1[49]), .Y(_858_) );
OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_857_), .B(_858_), .C(_72__1_), .Y(_859_) );
NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_859_), .B(_863_), .Y(_70__1_) );
OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_860_), .B(_857_), .C(_862_), .Y(_72__2_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(_72__2_), .Y(_867_) );
OR2X2 OR2X2_96 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_868_) );
NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_869_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_867_), .B(_869_), .C(_868_), .Y(_870_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_864_) );
AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[50]), .B(i_add_term1[50]), .Y(_865_) );
OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_864_), .B(_865_), .C(_72__2_), .Y(_866_) );
NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_866_), .B(_870_), .Y(_70__2_) );
OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_867_), .B(_864_), .C(_869_), .Y(_72__3_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(_73_), .Y(_871_) );
NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(w_cout_12_), .Y(_872_) );
OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_871_), .C(_872_), .Y(csa_inst_cin) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(_75__0_), .Y(_873_) );
NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_76__0_), .B(w_cout_12_), .Y(_874_) );
OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_873_), .C(_874_), .Y(_0__52_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(_75__1_), .Y(_875_) );
NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_76__1_), .Y(_876_) );
OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_875_), .C(_876_), .Y(_0__53_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(_75__2_), .Y(_877_) );
NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_76__2_), .Y(_878_) );
OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_877_), .C(_878_), .Y(_0__54_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(_75__3_), .Y(_879_) );
NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_76__3_), .Y(_880_) );
OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(w_cout_12_), .B(_879_), .C(_880_), .Y(_0__55_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_884_) );
OR2X2 OR2X2_97 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_885_) );
NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_886_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_884_), .B(_886_), .C(_885_), .Y(_887_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_881_) );
AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_882_) );
OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_882_), .C(gnd), .Y(_883_) );
NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_883_), .B(_887_), .Y(_75__0_) );
OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_884_), .B(_881_), .C(_886_), .Y(_77__1_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(_77__3_), .Y(_891_) );
OR2X2 OR2X2_98 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_892_) );
NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_893_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_891_), .B(_893_), .C(_892_), .Y(_894_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_888_) );
AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_889_) );
OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_888_), .B(_889_), .C(_77__3_), .Y(_890_) );
NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_890_), .B(_894_), .Y(_75__3_) );
OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_891_), .B(_888_), .C(_893_), .Y(_73_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(_77__1_), .Y(_898_) );
OR2X2 OR2X2_99 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_899_) );
NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_900_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_898_), .B(_900_), .C(_899_), .Y(_901_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_895_) );
AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_896_) );
OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_895_), .B(_896_), .C(_77__1_), .Y(_897_) );
NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_897_), .B(_901_), .Y(_75__1_) );
OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_898_), .B(_895_), .C(_900_), .Y(_77__2_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(_77__2_), .Y(_905_) );
OR2X2 OR2X2_100 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_906_) );
NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_907_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_905_), .B(_907_), .C(_906_), .Y(_908_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_902_) );
AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_903_) );
OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_902_), .B(_903_), .C(_77__2_), .Y(_904_) );
NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_904_), .B(_908_), .Y(_75__2_) );
OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_905_), .B(_902_), .C(_907_), .Y(_77__3_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_912_) );
OR2X2 OR2X2_101 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_913_) );
NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_914_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_912_), .B(_914_), .C(_913_), .Y(_915_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_909_) );
AND2X2 AND2X2_101 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[52]), .B(i_add_term1[52]), .Y(_910_) );
OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_910_), .C(vdd), .Y(_911_) );
NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_911_), .B(_915_), .Y(_76__0_) );
OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_912_), .B(_909_), .C(_914_), .Y(_78__1_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(_78__3_), .Y(_919_) );
OR2X2 OR2X2_102 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_920_) );
NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_921_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_919_), .B(_921_), .C(_920_), .Y(_922_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_916_) );
AND2X2 AND2X2_102 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[55]), .B(i_add_term1[55]), .Y(_917_) );
OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_916_), .B(_917_), .C(_78__3_), .Y(_918_) );
NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_918_), .B(_922_), .Y(_76__3_) );
OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_919_), .B(_916_), .C(_921_), .Y(_74_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(_78__1_), .Y(_926_) );
OR2X2 OR2X2_103 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_927_) );
NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_928_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_926_), .B(_928_), .C(_927_), .Y(_929_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_923_) );
AND2X2 AND2X2_103 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[53]), .B(i_add_term1[53]), .Y(_924_) );
OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_924_), .C(_78__1_), .Y(_925_) );
NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_925_), .B(_929_), .Y(_76__1_) );
OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_926_), .B(_923_), .C(_928_), .Y(_78__2_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(_78__2_), .Y(_933_) );
OR2X2 OR2X2_104 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_934_) );
NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_935_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_935_), .C(_934_), .Y(_936_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_930_) );
AND2X2 AND2X2_104 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[54]), .B(i_add_term1[54]), .Y(_931_) );
OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_931_), .C(_78__2_), .Y(_932_) );
NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_936_), .Y(_76__2_) );
OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_930_), .C(_935_), .Y(_78__3_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cout0_0), .Y(_937_) );
NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cout0_1), .B(csa_inst_cin), .Y(_938_) );
OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .B(_937_), .C(_938_), .Y(w_cout_14_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_0_fa0_o_sum), .Y(_939_) );
NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_1_fa0_o_sum), .B(csa_inst_cin), .Y(_940_) );
OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .B(_939_), .C(_940_), .Y(_0__56_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_0_fa1_o_sum), .Y(_941_) );
NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .B(csa_inst_rca0_1_fa1_o_sum), .Y(_942_) );
OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .B(_941_), .C(_942_), .Y(_0__57_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_0_fa2_o_sum), .Y(_943_) );
NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .B(csa_inst_rca0_1_fa2_o_sum), .Y(_944_) );
OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .B(_943_), .C(_944_), .Y(_0__58_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_948_) );
OR2X2 OR2X2_105 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_949_) );
NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_950_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_948_), .B(_950_), .C(_949_), .Y(_951_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_945_) );
AND2X2 AND2X2_105 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_946_) );
OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_945_), .B(_946_), .C(gnd), .Y(_947_) );
NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_947_), .B(_951_), .Y(csa_inst_rca0_0_fa0_o_sum) );
OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_948_), .B(_945_), .C(_950_), .Y(csa_inst_rca0_0_fa0_o_carry) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_0_fa0_o_carry), .Y(_955_) );
OR2X2 OR2X2_106 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_956_) );
NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_957_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_955_), .B(_957_), .C(_956_), .Y(_958_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_952_) );
AND2X2 AND2X2_106 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_953_) );
OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_952_), .B(_953_), .C(csa_inst_rca0_0_fa0_o_carry), .Y(_954_) );
NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_954_), .B(_958_), .Y(csa_inst_rca0_0_fa1_o_sum) );
OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_955_), .B(_952_), .C(_957_), .Y(csa_inst_rca0_0_fa1_o_carry) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_0_fa1_o_carry), .Y(_962_) );
OR2X2 OR2X2_107 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_963_) );
NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_964_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_964_), .C(_963_), .Y(_965_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_959_) );
AND2X2 AND2X2_107 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_960_) );
OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_959_), .B(_960_), .C(csa_inst_rca0_0_fa1_o_carry), .Y(_961_) );
NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_961_), .B(_965_), .Y(csa_inst_rca0_0_fa2_o_sum) );
OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_959_), .C(_964_), .Y(csa_inst_cout0_0) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(vdd), .Y(_969_) );
OR2X2 OR2X2_108 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_970_) );
NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_971_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_969_), .B(_971_), .C(_970_), .Y(_972_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_966_) );
AND2X2 AND2X2_108 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[56]), .B(i_add_term1[56]), .Y(_967_) );
OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_966_), .B(_967_), .C(vdd), .Y(_968_) );
NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_968_), .B(_972_), .Y(csa_inst_rca0_1_fa0_o_sum) );
OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_969_), .B(_966_), .C(_971_), .Y(csa_inst_rca0_1_fa0_o_carry) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_1_fa0_o_carry), .Y(_976_) );
OR2X2 OR2X2_109 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_977_) );
NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_978_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(_978_), .C(_977_), .Y(_979_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_973_) );
AND2X2 AND2X2_109 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[57]), .B(i_add_term1[57]), .Y(_974_) );
OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_973_), .B(_974_), .C(csa_inst_rca0_1_fa0_o_carry), .Y(_975_) );
NAND2X1 NAND2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_975_), .B(_979_), .Y(csa_inst_rca0_1_fa1_o_sum) );
OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(_973_), .C(_978_), .Y(csa_inst_rca0_1_fa1_o_carry) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_rca0_1_fa1_o_carry), .Y(_983_) );
OR2X2 OR2X2_110 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_984_) );
NAND2X1 NAND2X1_288 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_985_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_985_), .C(_984_), .Y(_986_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_980_) );
AND2X2 AND2X2_110 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[58]), .B(i_add_term1[58]), .Y(_981_) );
OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_980_), .B(_981_), .C(csa_inst_rca0_1_fa1_o_carry), .Y(_982_) );
NAND2X1 NAND2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_982_), .B(_986_), .Y(csa_inst_rca0_1_fa2_o_sum) );
OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_980_), .C(_985_), .Y(csa_inst_cout0_1) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_990_) );
OR2X2 OR2X2_111 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_991_) );
NAND2X1 NAND2X1_290 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_992_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_992_), .C(_991_), .Y(_993_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_987_) );
AND2X2 AND2X2_111 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[0]), .B(i_add_term1[0]), .Y(_988_) );
OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_987_), .B(_988_), .C(gnd), .Y(_989_) );
NAND2X1 NAND2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_989_), .B(_993_), .Y(rca_inst_fa0_o_sum) );
OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_987_), .C(_992_), .Y(rca_inst_fa0_o_carry) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_i_carry), .Y(_997_) );
OR2X2 OR2X2_112 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_998_) );
NAND2X1 NAND2X1_292 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_999_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_997_), .B(_999_), .C(_998_), .Y(_1000_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_994_) );
AND2X2 AND2X2_112 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[3]), .B(i_add_term1[3]), .Y(_995_) );
OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_994_), .B(_995_), .C(rca_inst_fa3_i_carry), .Y(_996_) );
NAND2X1 NAND2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_996_), .B(_1000_), .Y(rca_inst_fa3_o_sum) );
OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_997_), .B(_994_), .C(_999_), .Y(rca_inst_cout) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_carry), .Y(_1004_) );
OR2X2 OR2X2_113 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1005_) );
NAND2X1 NAND2X1_294 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1006_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .B(_1006_), .C(_1005_), .Y(_1007_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1001_) );
AND2X2 AND2X2_113 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[1]), .B(i_add_term1[1]), .Y(_1002_) );
OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .B(_1002_), .C(rca_inst_fa0_o_carry), .Y(_1003_) );
NAND2X1 NAND2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_1003_), .B(_1007_), .Y(rca_inst_fa_1__o_sum) );
OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .B(_1001_), .C(_1006_), .Y(rca_inst_fa_1__o_carry) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_carry), .Y(_1011_) );
OR2X2 OR2X2_114 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1012_) );
NAND2X1 NAND2X1_296 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1013_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .B(_1013_), .C(_1012_), .Y(_1014_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1008_) );
AND2X2 AND2X2_114 ( .gnd(gnd), .vdd(vdd), .A(i_add_term2[2]), .B(i_add_term1[2]), .Y(_1009_) );
OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1008_), .B(_1009_), .C(rca_inst_fa_1__o_carry), .Y(_1010_) );
NAND2X1 NAND2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_1010_), .B(_1014_), .Y(rca_inst_fa_2__o_sum) );
OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .B(_1008_), .C(_1013_), .Y(rca_inst_fa3_i_carry) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa0_o_sum), .Y(_0__0_) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_1__o_sum), .Y(_0__1_) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa_2__o_sum), .Y(_0__2_) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_fa3_o_sum), .Y(_0__3_) );
BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(rca_inst_cout), .Y(w_cout_0_) );
BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(csa_inst_cin), .Y(w_cout_13_) );
endmodule
