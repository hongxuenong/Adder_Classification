module cla_19bit (i_add1[0], i_add1[1], i_add1[2], i_add1[3], i_add1[4], i_add1[5], i_add1[6], i_add1[7], i_add1[8], i_add1[9], i_add1[10], i_add1[11], i_add1[12], i_add1[13], i_add1[14], i_add1[15], i_add1[16], i_add1[17], i_add1[18], i_add2[0], i_add2[1], i_add2[2], i_add2[3], i_add2[4], i_add2[5], i_add2[6], i_add2[7], i_add2[8], i_add2[9], i_add2[10], i_add2[11], i_add2[12], i_add2[13], i_add2[14], i_add2[15], i_add2[16], i_add2[17], i_add2[18], o_result[0], o_result[1], o_result[2], o_result[3], o_result[4], o_result[5], o_result[6], o_result[7], o_result[8], o_result[9], o_result[10], o_result[11], o_result[12], o_result[13], o_result[14], o_result[15], o_result[16], o_result[17], o_result[18], o_result[19]);

input i_add1[0];
input i_add1[1];
input i_add1[2];
input i_add1[3];
input i_add1[4];
input i_add1[5];
input i_add1[6];
input i_add1[7];
input i_add1[8];
input i_add1[9];
input i_add1[10];
input i_add1[11];
input i_add1[12];
input i_add1[13];
input i_add1[14];
input i_add1[15];
input i_add1[16];
input i_add1[17];
input i_add1[18];
input i_add2[0];
input i_add2[1];
input i_add2[2];
input i_add2[3];
input i_add2[4];
input i_add2[5];
input i_add2[6];
input i_add2[7];
input i_add2[8];
input i_add2[9];
input i_add2[10];
input i_add2[11];
input i_add2[12];
input i_add2[13];
input i_add2[14];
input i_add2[15];
input i_add2[16];
input i_add2[17];
input i_add2[18];
output o_result[0];
output o_result[1];
output o_result[2];
output o_result[3];
output o_result[4];
output o_result[5];
output o_result[6];
output o_result[7];
output o_result[8];
output o_result[9];
output o_result[10];
output o_result[11];
output o_result[12];
output o_result[13];
output o_result[14];
output o_result[15];
output o_result[16];
output o_result[17];
output o_result[18];
output o_result[19];

NAND2X1 NAND2X1_1 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_57_) );
INVX1 INVX1_1 ( .A(_57_), .Y(w_C_1_) );
NAND2X1 NAND2X1_2 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_58_) );
NAND2X1 NAND2X1_3 ( .A(_57_), .B(_58_), .Y(_59_) );
OAI21X1 OAI21X1_1 ( .A(i_add2[1]), .B(i_add1[1]), .C(_59_), .Y(_60_) );
INVX1 INVX1_2 ( .A(_60_), .Y(w_C_2_) );
NAND2X1 NAND2X1_4 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_61_) );
OR2X2 OR2X2_1 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_62_) );
OR2X2 OR2X2_2 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_63_) );
NAND3X1 NAND3X1_1 ( .A(_62_), .B(_63_), .C(_59_), .Y(_64_) );
NAND2X1 NAND2X1_5 ( .A(_61_), .B(_64_), .Y(w_C_3_) );
INVX1 INVX1_3 ( .A(i_add2[3]), .Y(_65_) );
INVX1 INVX1_4 ( .A(i_add1[3]), .Y(_66_) );
NAND2X1 NAND2X1_6 ( .A(_65_), .B(_66_), .Y(_67_) );
NAND2X1 NAND2X1_7 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_68_) );
NAND3X1 NAND3X1_2 ( .A(_61_), .B(_68_), .C(_64_), .Y(_69_) );
AND2X2 AND2X2_1 ( .A(_69_), .B(_67_), .Y(w_C_4_) );
NAND2X1 NAND2X1_8 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_70_) );
OR2X2 OR2X2_3 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_71_) );
NAND3X1 NAND3X1_3 ( .A(_67_), .B(_71_), .C(_69_), .Y(_72_) );
NAND2X1 NAND2X1_9 ( .A(_70_), .B(_72_), .Y(w_C_5_) );
NAND2X1 NAND2X1_10 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_73_) );
NAND3X1 NAND3X1_4 ( .A(_70_), .B(_73_), .C(_72_), .Y(_74_) );
OAI21X1 OAI21X1_2 ( .A(i_add2[5]), .B(i_add1[5]), .C(_74_), .Y(_75_) );
INVX1 INVX1_5 ( .A(_75_), .Y(w_C_6_) );
INVX1 INVX1_6 ( .A(i_add2[6]), .Y(_76_) );
INVX1 INVX1_7 ( .A(i_add1[6]), .Y(_77_) );
NOR2X1 NOR2X1_1 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_78_) );
INVX1 INVX1_8 ( .A(_78_), .Y(_79_) );
NOR2X1 NOR2X1_2 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_80_) );
INVX1 INVX1_9 ( .A(_80_), .Y(_81_) );
NAND3X1 NAND3X1_5 ( .A(_79_), .B(_81_), .C(_74_), .Y(_82_) );
OAI21X1 OAI21X1_3 ( .A(_76_), .B(_77_), .C(_82_), .Y(w_C_7_) );
NOR2X1 NOR2X1_3 ( .A(_76_), .B(_77_), .Y(_83_) );
INVX1 INVX1_10 ( .A(_83_), .Y(_84_) );
AND2X2 AND2X2_2 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_85_) );
INVX1 INVX1_11 ( .A(_85_), .Y(_86_) );
NAND3X1 NAND3X1_6 ( .A(_84_), .B(_86_), .C(_82_), .Y(_87_) );
OAI21X1 OAI21X1_4 ( .A(i_add2[7]), .B(i_add1[7]), .C(_87_), .Y(_88_) );
INVX1 INVX1_12 ( .A(_88_), .Y(w_C_8_) );
INVX1 INVX1_13 ( .A(i_add2[8]), .Y(_89_) );
INVX1 INVX1_14 ( .A(i_add1[8]), .Y(_90_) );
NOR2X1 NOR2X1_4 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_0_) );
INVX1 INVX1_15 ( .A(_0_), .Y(_1_) );
NOR2X1 NOR2X1_5 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_2_) );
INVX1 INVX1_16 ( .A(_2_), .Y(_3_) );
NAND3X1 NAND3X1_7 ( .A(_1_), .B(_3_), .C(_87_), .Y(_4_) );
OAI21X1 OAI21X1_5 ( .A(_89_), .B(_90_), .C(_4_), .Y(w_C_9_) );
NOR2X1 NOR2X1_6 ( .A(_89_), .B(_90_), .Y(_5_) );
INVX1 INVX1_17 ( .A(_5_), .Y(_6_) );
AND2X2 AND2X2_3 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_7_) );
INVX1 INVX1_18 ( .A(_7_), .Y(_8_) );
NAND3X1 NAND3X1_8 ( .A(_6_), .B(_8_), .C(_4_), .Y(_9_) );
OAI21X1 OAI21X1_6 ( .A(i_add2[9]), .B(i_add1[9]), .C(_9_), .Y(_10_) );
INVX1 INVX1_19 ( .A(_10_), .Y(w_C_10_) );
INVX1 INVX1_20 ( .A(i_add2[10]), .Y(_11_) );
INVX1 INVX1_21 ( .A(i_add1[10]), .Y(_12_) );
NOR2X1 NOR2X1_7 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_13_) );
INVX1 INVX1_22 ( .A(_13_), .Y(_14_) );
NOR2X1 NOR2X1_8 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_15_) );
INVX1 INVX1_23 ( .A(_15_), .Y(_16_) );
NAND3X1 NAND3X1_9 ( .A(_14_), .B(_16_), .C(_9_), .Y(_17_) );
OAI21X1 OAI21X1_7 ( .A(_11_), .B(_12_), .C(_17_), .Y(w_C_11_) );
NOR2X1 NOR2X1_9 ( .A(_11_), .B(_12_), .Y(_18_) );
INVX1 INVX1_24 ( .A(_18_), .Y(_19_) );
AND2X2 AND2X2_4 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_20_) );
INVX1 INVX1_25 ( .A(_20_), .Y(_21_) );
NAND3X1 NAND3X1_10 ( .A(_19_), .B(_21_), .C(_17_), .Y(_22_) );
OAI21X1 OAI21X1_8 ( .A(i_add2[11]), .B(i_add1[11]), .C(_22_), .Y(_23_) );
INVX1 INVX1_26 ( .A(_23_), .Y(w_C_12_) );
INVX1 INVX1_27 ( .A(i_add2[12]), .Y(_24_) );
INVX1 INVX1_28 ( .A(i_add1[12]), .Y(_25_) );
NOR2X1 NOR2X1_10 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_26_) );
INVX1 INVX1_29 ( .A(_26_), .Y(_27_) );
NOR2X1 NOR2X1_11 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_28_) );
INVX1 INVX1_30 ( .A(_28_), .Y(_29_) );
NAND3X1 NAND3X1_11 ( .A(_27_), .B(_29_), .C(_22_), .Y(_30_) );
OAI21X1 OAI21X1_9 ( .A(_24_), .B(_25_), .C(_30_), .Y(w_C_13_) );
NOR2X1 NOR2X1_12 ( .A(_24_), .B(_25_), .Y(_31_) );
INVX1 INVX1_31 ( .A(_31_), .Y(_32_) );
AND2X2 AND2X2_5 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_33_) );
INVX1 INVX1_32 ( .A(_33_), .Y(_34_) );
NAND3X1 NAND3X1_12 ( .A(_32_), .B(_34_), .C(_30_), .Y(_35_) );
OAI21X1 OAI21X1_10 ( .A(i_add2[13]), .B(i_add1[13]), .C(_35_), .Y(_36_) );
INVX1 INVX1_33 ( .A(_36_), .Y(w_C_14_) );
NAND2X1 NAND2X1_11 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_37_) );
NOR2X1 NOR2X1_13 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_38_) );
OAI21X1 OAI21X1_11 ( .A(_38_), .B(_36_), .C(_37_), .Y(w_C_15_) );
OR2X2 OR2X2_4 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_39_) );
NOR2X1 NOR2X1_14 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_40_) );
INVX1 INVX1_34 ( .A(_40_), .Y(_41_) );
INVX1 INVX1_35 ( .A(_38_), .Y(_42_) );
NAND3X1 NAND3X1_13 ( .A(_41_), .B(_42_), .C(_35_), .Y(_43_) );
NAND2X1 NAND2X1_12 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_44_) );
NAND3X1 NAND3X1_14 ( .A(_37_), .B(_44_), .C(_43_), .Y(_45_) );
AND2X2 AND2X2_6 ( .A(_45_), .B(_39_), .Y(w_C_16_) );
INVX1 INVX1_36 ( .A(i_add2[16]), .Y(_46_) );
INVX1 INVX1_37 ( .A(i_add1[16]), .Y(_47_) );
NAND2X1 NAND2X1_13 ( .A(_46_), .B(_47_), .Y(_48_) );
NAND3X1 NAND3X1_15 ( .A(_39_), .B(_48_), .C(_45_), .Y(_49_) );
OAI21X1 OAI21X1_12 ( .A(_46_), .B(_47_), .C(_49_), .Y(w_C_17_) );
OR2X2 OR2X2_5 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_50_) );
NAND2X1 NAND2X1_14 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_51_) );
NAND2X1 NAND2X1_15 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_52_) );
NAND3X1 NAND3X1_16 ( .A(_51_), .B(_52_), .C(_49_), .Y(_53_) );
AND2X2 AND2X2_7 ( .A(_53_), .B(_50_), .Y(w_C_18_) );
NAND2X1 NAND2X1_16 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_54_) );
OR2X2 OR2X2_6 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_55_) );
NAND3X1 NAND3X1_17 ( .A(_50_), .B(_55_), .C(_53_), .Y(_56_) );
NAND2X1 NAND2X1_17 ( .A(_54_), .B(_56_), .Y(w_C_19_) );
BUFX2 BUFX2_1 ( .A(_91__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .A(_91__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .A(_91__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .A(_91__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .A(_91__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .A(_91__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .A(_91__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .A(_91__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .A(_91__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .A(_91__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .A(_91__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .A(_91__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .A(_91__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .A(_91__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .A(_91__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .A(_91__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .A(_91__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .A(_91__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .A(_91__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .A(w_C_19_), .Y(o_result[19]) );
INVX1 INVX1_38 ( .A(w_C_4_), .Y(_95_) );
OR2X2 OR2X2_7 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_96_) );
NAND2X1 NAND2X1_18 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_97_) );
NAND3X1 NAND3X1_18 ( .A(_95_), .B(_97_), .C(_96_), .Y(_98_) );
NOR2X1 NOR2X1_15 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_92_) );
AND2X2 AND2X2_8 ( .A(i_add2[4]), .B(i_add1[4]), .Y(_93_) );
OAI21X1 OAI21X1_13 ( .A(_92_), .B(_93_), .C(w_C_4_), .Y(_94_) );
NAND2X1 NAND2X1_19 ( .A(_94_), .B(_98_), .Y(_91__4_) );
INVX1 INVX1_39 ( .A(w_C_5_), .Y(_102_) );
OR2X2 OR2X2_8 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_103_) );
NAND2X1 NAND2X1_20 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_104_) );
NAND3X1 NAND3X1_19 ( .A(_102_), .B(_104_), .C(_103_), .Y(_105_) );
NOR2X1 NOR2X1_16 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_99_) );
AND2X2 AND2X2_9 ( .A(i_add2[5]), .B(i_add1[5]), .Y(_100_) );
OAI21X1 OAI21X1_14 ( .A(_99_), .B(_100_), .C(w_C_5_), .Y(_101_) );
NAND2X1 NAND2X1_21 ( .A(_101_), .B(_105_), .Y(_91__5_) );
INVX1 INVX1_40 ( .A(w_C_6_), .Y(_109_) );
OR2X2 OR2X2_9 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_110_) );
NAND2X1 NAND2X1_22 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_111_) );
NAND3X1 NAND3X1_20 ( .A(_109_), .B(_111_), .C(_110_), .Y(_112_) );
NOR2X1 NOR2X1_17 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_106_) );
AND2X2 AND2X2_10 ( .A(i_add2[6]), .B(i_add1[6]), .Y(_107_) );
OAI21X1 OAI21X1_15 ( .A(_106_), .B(_107_), .C(w_C_6_), .Y(_108_) );
NAND2X1 NAND2X1_23 ( .A(_108_), .B(_112_), .Y(_91__6_) );
INVX1 INVX1_41 ( .A(w_C_7_), .Y(_116_) );
OR2X2 OR2X2_10 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_117_) );
NAND2X1 NAND2X1_24 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_118_) );
NAND3X1 NAND3X1_21 ( .A(_116_), .B(_118_), .C(_117_), .Y(_119_) );
NOR2X1 NOR2X1_18 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_113_) );
AND2X2 AND2X2_11 ( .A(i_add2[7]), .B(i_add1[7]), .Y(_114_) );
OAI21X1 OAI21X1_16 ( .A(_113_), .B(_114_), .C(w_C_7_), .Y(_115_) );
NAND2X1 NAND2X1_25 ( .A(_115_), .B(_119_), .Y(_91__7_) );
INVX1 INVX1_42 ( .A(w_C_8_), .Y(_123_) );
OR2X2 OR2X2_11 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_124_) );
NAND2X1 NAND2X1_26 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_125_) );
NAND3X1 NAND3X1_22 ( .A(_123_), .B(_125_), .C(_124_), .Y(_126_) );
NOR2X1 NOR2X1_19 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_120_) );
AND2X2 AND2X2_12 ( .A(i_add2[8]), .B(i_add1[8]), .Y(_121_) );
OAI21X1 OAI21X1_17 ( .A(_120_), .B(_121_), .C(w_C_8_), .Y(_122_) );
NAND2X1 NAND2X1_27 ( .A(_122_), .B(_126_), .Y(_91__8_) );
INVX1 INVX1_43 ( .A(w_C_9_), .Y(_130_) );
OR2X2 OR2X2_12 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_131_) );
NAND2X1 NAND2X1_28 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_132_) );
NAND3X1 NAND3X1_23 ( .A(_130_), .B(_132_), .C(_131_), .Y(_133_) );
NOR2X1 NOR2X1_20 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_127_) );
AND2X2 AND2X2_13 ( .A(i_add2[9]), .B(i_add1[9]), .Y(_128_) );
OAI21X1 OAI21X1_18 ( .A(_127_), .B(_128_), .C(w_C_9_), .Y(_129_) );
NAND2X1 NAND2X1_29 ( .A(_129_), .B(_133_), .Y(_91__9_) );
INVX1 INVX1_44 ( .A(w_C_10_), .Y(_137_) );
OR2X2 OR2X2_13 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_138_) );
NAND2X1 NAND2X1_30 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_139_) );
NAND3X1 NAND3X1_24 ( .A(_137_), .B(_139_), .C(_138_), .Y(_140_) );
NOR2X1 NOR2X1_21 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_134_) );
AND2X2 AND2X2_14 ( .A(i_add2[10]), .B(i_add1[10]), .Y(_135_) );
OAI21X1 OAI21X1_19 ( .A(_134_), .B(_135_), .C(w_C_10_), .Y(_136_) );
NAND2X1 NAND2X1_31 ( .A(_136_), .B(_140_), .Y(_91__10_) );
INVX1 INVX1_45 ( .A(w_C_11_), .Y(_144_) );
OR2X2 OR2X2_14 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_145_) );
NAND2X1 NAND2X1_32 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_146_) );
NAND3X1 NAND3X1_25 ( .A(_144_), .B(_146_), .C(_145_), .Y(_147_) );
NOR2X1 NOR2X1_22 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_141_) );
AND2X2 AND2X2_15 ( .A(i_add2[11]), .B(i_add1[11]), .Y(_142_) );
OAI21X1 OAI21X1_20 ( .A(_141_), .B(_142_), .C(w_C_11_), .Y(_143_) );
NAND2X1 NAND2X1_33 ( .A(_143_), .B(_147_), .Y(_91__11_) );
INVX1 INVX1_46 ( .A(w_C_12_), .Y(_151_) );
OR2X2 OR2X2_15 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_152_) );
NAND2X1 NAND2X1_34 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_153_) );
NAND3X1 NAND3X1_26 ( .A(_151_), .B(_153_), .C(_152_), .Y(_154_) );
NOR2X1 NOR2X1_23 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_148_) );
AND2X2 AND2X2_16 ( .A(i_add2[12]), .B(i_add1[12]), .Y(_149_) );
OAI21X1 OAI21X1_21 ( .A(_148_), .B(_149_), .C(w_C_12_), .Y(_150_) );
NAND2X1 NAND2X1_35 ( .A(_150_), .B(_154_), .Y(_91__12_) );
INVX1 INVX1_47 ( .A(w_C_13_), .Y(_158_) );
OR2X2 OR2X2_16 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_159_) );
NAND2X1 NAND2X1_36 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_160_) );
NAND3X1 NAND3X1_27 ( .A(_158_), .B(_160_), .C(_159_), .Y(_161_) );
NOR2X1 NOR2X1_24 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_155_) );
AND2X2 AND2X2_17 ( .A(i_add2[13]), .B(i_add1[13]), .Y(_156_) );
OAI21X1 OAI21X1_22 ( .A(_155_), .B(_156_), .C(w_C_13_), .Y(_157_) );
NAND2X1 NAND2X1_37 ( .A(_157_), .B(_161_), .Y(_91__13_) );
INVX1 INVX1_48 ( .A(w_C_14_), .Y(_165_) );
OR2X2 OR2X2_17 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_166_) );
NAND2X1 NAND2X1_38 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_167_) );
NAND3X1 NAND3X1_28 ( .A(_165_), .B(_167_), .C(_166_), .Y(_168_) );
NOR2X1 NOR2X1_25 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_162_) );
AND2X2 AND2X2_18 ( .A(i_add2[14]), .B(i_add1[14]), .Y(_163_) );
OAI21X1 OAI21X1_23 ( .A(_162_), .B(_163_), .C(w_C_14_), .Y(_164_) );
NAND2X1 NAND2X1_39 ( .A(_164_), .B(_168_), .Y(_91__14_) );
INVX1 INVX1_49 ( .A(w_C_15_), .Y(_172_) );
OR2X2 OR2X2_18 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_173_) );
NAND2X1 NAND2X1_40 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_174_) );
NAND3X1 NAND3X1_29 ( .A(_172_), .B(_174_), .C(_173_), .Y(_175_) );
NOR2X1 NOR2X1_26 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_169_) );
AND2X2 AND2X2_19 ( .A(i_add2[15]), .B(i_add1[15]), .Y(_170_) );
OAI21X1 OAI21X1_24 ( .A(_169_), .B(_170_), .C(w_C_15_), .Y(_171_) );
NAND2X1 NAND2X1_41 ( .A(_171_), .B(_175_), .Y(_91__15_) );
INVX1 INVX1_50 ( .A(w_C_16_), .Y(_179_) );
OR2X2 OR2X2_19 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_180_) );
NAND2X1 NAND2X1_42 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_181_) );
NAND3X1 NAND3X1_30 ( .A(_179_), .B(_181_), .C(_180_), .Y(_182_) );
NOR2X1 NOR2X1_27 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_176_) );
AND2X2 AND2X2_20 ( .A(i_add2[16]), .B(i_add1[16]), .Y(_177_) );
OAI21X1 OAI21X1_25 ( .A(_176_), .B(_177_), .C(w_C_16_), .Y(_178_) );
NAND2X1 NAND2X1_43 ( .A(_178_), .B(_182_), .Y(_91__16_) );
INVX1 INVX1_51 ( .A(w_C_17_), .Y(_186_) );
OR2X2 OR2X2_20 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_187_) );
NAND2X1 NAND2X1_44 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_188_) );
NAND3X1 NAND3X1_31 ( .A(_186_), .B(_188_), .C(_187_), .Y(_189_) );
NOR2X1 NOR2X1_28 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_183_) );
AND2X2 AND2X2_21 ( .A(i_add2[17]), .B(i_add1[17]), .Y(_184_) );
OAI21X1 OAI21X1_26 ( .A(_183_), .B(_184_), .C(w_C_17_), .Y(_185_) );
NAND2X1 NAND2X1_45 ( .A(_185_), .B(_189_), .Y(_91__17_) );
INVX1 INVX1_52 ( .A(w_C_18_), .Y(_193_) );
OR2X2 OR2X2_21 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_194_) );
NAND2X1 NAND2X1_46 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_195_) );
NAND3X1 NAND3X1_32 ( .A(_193_), .B(_195_), .C(_194_), .Y(_196_) );
NOR2X1 NOR2X1_29 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_190_) );
AND2X2 AND2X2_22 ( .A(i_add2[18]), .B(i_add1[18]), .Y(_191_) );
OAI21X1 OAI21X1_27 ( .A(_190_), .B(_191_), .C(w_C_18_), .Y(_192_) );
NAND2X1 NAND2X1_47 ( .A(_192_), .B(_196_), .Y(_91__18_) );
INVX1 INVX1_53 ( .A(1'b0), .Y(_200_) );
OR2X2 OR2X2_22 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_201_) );
NAND2X1 NAND2X1_48 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_202_) );
NAND3X1 NAND3X1_33 ( .A(_200_), .B(_202_), .C(_201_), .Y(_203_) );
NOR2X1 NOR2X1_30 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_197_) );
AND2X2 AND2X2_23 ( .A(i_add2[0]), .B(i_add1[0]), .Y(_198_) );
OAI21X1 OAI21X1_28 ( .A(_197_), .B(_198_), .C(1'b0), .Y(_199_) );
NAND2X1 NAND2X1_49 ( .A(_199_), .B(_203_), .Y(_91__0_) );
INVX1 INVX1_54 ( .A(w_C_1_), .Y(_207_) );
OR2X2 OR2X2_23 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_208_) );
NAND2X1 NAND2X1_50 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_209_) );
NAND3X1 NAND3X1_34 ( .A(_207_), .B(_209_), .C(_208_), .Y(_210_) );
NOR2X1 NOR2X1_31 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_204_) );
AND2X2 AND2X2_24 ( .A(i_add2[1]), .B(i_add1[1]), .Y(_205_) );
OAI21X1 OAI21X1_29 ( .A(_204_), .B(_205_), .C(w_C_1_), .Y(_206_) );
NAND2X1 NAND2X1_51 ( .A(_206_), .B(_210_), .Y(_91__1_) );
INVX1 INVX1_55 ( .A(w_C_2_), .Y(_214_) );
OR2X2 OR2X2_24 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_215_) );
NAND2X1 NAND2X1_52 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_216_) );
NAND3X1 NAND3X1_35 ( .A(_214_), .B(_216_), .C(_215_), .Y(_217_) );
NOR2X1 NOR2X1_32 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_211_) );
AND2X2 AND2X2_25 ( .A(i_add2[2]), .B(i_add1[2]), .Y(_212_) );
OAI21X1 OAI21X1_30 ( .A(_211_), .B(_212_), .C(w_C_2_), .Y(_213_) );
NAND2X1 NAND2X1_53 ( .A(_213_), .B(_217_), .Y(_91__2_) );
INVX1 INVX1_56 ( .A(w_C_3_), .Y(_221_) );
OR2X2 OR2X2_25 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_222_) );
NAND2X1 NAND2X1_54 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_223_) );
NAND3X1 NAND3X1_36 ( .A(_221_), .B(_223_), .C(_222_), .Y(_224_) );
NOR2X1 NOR2X1_33 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_218_) );
AND2X2 AND2X2_26 ( .A(i_add2[3]), .B(i_add1[3]), .Y(_219_) );
OAI21X1 OAI21X1_31 ( .A(_218_), .B(_219_), .C(w_C_3_), .Y(_220_) );
NAND2X1 NAND2X1_55 ( .A(_220_), .B(_224_), .Y(_91__3_) );
BUFX2 BUFX2_21 ( .A(w_C_19_), .Y(_91__19_) );
BUFX2 BUFX2_22 ( .A(1'b0), .Y(w_C_0_) );
endmodule
