module cla_40bit ( gnd, vdd, i_add1, i_add2, o_result);

input gnd, vdd;
input [39:0] i_add1;
input [39:0] i_add2;
output [40:0] o_result;

NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_381_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_382_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_382_), .C(w_C_25_), .Y(_383_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_387_), .Y(_233__25_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(w_C_26_), .Y(_391_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_392_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_393_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_393_), .C(_392_), .Y(_394_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_388_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_389_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_388_), .B(_389_), .C(w_C_26_), .Y(_390_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_394_), .Y(_233__26_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(w_C_27_), .Y(_398_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_399_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_400_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_400_), .C(_399_), .Y(_401_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_395_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_396_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_395_), .B(_396_), .C(w_C_27_), .Y(_397_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_401_), .Y(_233__27_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(w_C_28_), .Y(_405_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_406_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_407_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_407_), .C(_406_), .Y(_408_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_402_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_403_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_403_), .C(w_C_28_), .Y(_404_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_408_), .Y(_233__28_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(w_C_29_), .Y(_412_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_413_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_414_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_414_), .C(_413_), .Y(_415_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_409_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_410_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_410_), .C(w_C_29_), .Y(_411_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_415_), .Y(_233__29_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(w_C_30_), .Y(_419_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_420_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_421_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_421_), .C(_420_), .Y(_422_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_416_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_417_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_417_), .C(w_C_30_), .Y(_418_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_422_), .Y(_233__30_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(w_C_31_), .Y(_426_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_427_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_428_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_428_), .C(_427_), .Y(_429_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_423_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_424_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_424_), .C(w_C_31_), .Y(_425_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(_429_), .Y(_233__31_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(w_C_32_), .Y(_433_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_434_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_435_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_433_), .B(_435_), .C(_434_), .Y(_436_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_430_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_431_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_431_), .C(w_C_32_), .Y(_432_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_432_), .B(_436_), .Y(_233__32_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(w_C_33_), .Y(_440_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_441_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_442_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_442_), .C(_441_), .Y(_443_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_437_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_438_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_438_), .C(w_C_33_), .Y(_439_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_443_), .Y(_233__33_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(w_C_34_), .Y(_447_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_448_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_449_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_447_), .B(_449_), .C(_448_), .Y(_450_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_444_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_445_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_445_), .C(w_C_34_), .Y(_446_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(_450_), .Y(_233__34_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(w_C_35_), .Y(_454_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_455_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_456_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_454_), .B(_456_), .C(_455_), .Y(_457_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_451_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .Y(_452_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_452_), .C(w_C_35_), .Y(_453_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(_457_), .Y(_233__35_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(w_C_36_), .Y(_461_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_462_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_463_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_463_), .C(_462_), .Y(_464_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_458_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_459_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_459_), .C(w_C_36_), .Y(_460_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_464_), .Y(_233__36_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(w_C_37_), .Y(_468_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_469_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_470_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_468_), .B(_470_), .C(_469_), .Y(_471_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_465_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_466_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_466_), .C(w_C_37_), .Y(_467_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_467_), .B(_471_), .Y(_233__37_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(w_C_38_), .Y(_475_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_476_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_477_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_477_), .C(_476_), .Y(_478_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_472_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_473_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_473_), .C(w_C_38_), .Y(_474_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_474_), .B(_478_), .Y(_233__38_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(w_C_39_), .Y(_482_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_483_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_484_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_482_), .B(_484_), .C(_483_), .Y(_485_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_479_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_480_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_480_), .C(w_C_39_), .Y(_481_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_485_), .Y(_233__39_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_489_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_490_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_491_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_491_), .C(_490_), .Y(_492_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_486_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_487_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_487_), .C(gnd), .Y(_488_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_492_), .Y(_233__0_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(w_C_1_), .Y(_496_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_497_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_498_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_498_), .C(_497_), .Y(_499_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_493_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_494_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_494_), .C(w_C_1_), .Y(_495_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_495_), .B(_499_), .Y(_233__1_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(w_C_2_), .Y(_503_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_504_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_505_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_505_), .C(_504_), .Y(_506_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_500_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_501_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_501_), .C(w_C_2_), .Y(_502_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_502_), .B(_506_), .Y(_233__2_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(w_C_3_), .Y(_510_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_511_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_512_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_510_), .B(_512_), .C(_511_), .Y(_513_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_507_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_508_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_508_), .C(w_C_3_), .Y(_509_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_509_), .B(_513_), .Y(_233__3_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .Y(_0_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(w_C_1_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[1]), .B(i_add1[1]), .Y(_1_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(i_add2[0]), .B(i_add1[0]), .C(i_add2[1]), .D(i_add1[1]), .Y(_2_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_2_), .Y(w_C_2_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_3_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_2_), .C(_3_), .Y(_4_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .C(_4_), .Y(_5_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_5_), .Y(w_C_3_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_6_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(i_add2[2]), .B(i_add1[2]), .Y(_7_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[3]), .B(i_add1[3]), .Y(_8_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_8_), .C(_4_), .Y(_9_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_9_), .Y(w_C_4_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_10_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_6_), .B(_10_), .C(_9_), .Y(_11_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .C(_11_), .Y(_12_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_12_), .Y(w_C_5_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .Y(_13_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add1[5]), .Y(_14_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_15_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_15_), .Y(_16_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_17_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_17_), .Y(_18_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_18_), .C(_11_), .Y(_19_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_14_), .C(_19_), .Y(w_C_6_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_14_), .Y(_20_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_20_), .Y(_21_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_22_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(_23_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_23_), .C(_19_), .Y(_24_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .C(_24_), .Y(_25_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(w_C_7_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .Y(_26_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add1[7]), .Y(_27_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_28_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_28_), .Y(_29_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_30_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_31_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_31_), .C(_24_), .Y(_32_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_27_), .C(_32_), .Y(w_C_8_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_27_), .Y(_33_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_33_), .Y(_34_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_35_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_35_), .Y(_36_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_36_), .C(_32_), .Y(_37_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .C(_37_), .Y(_38_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_38_), .Y(w_C_9_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .Y(_39_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add1[9]), .Y(_40_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_41_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_41_), .Y(_42_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_43_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_43_), .Y(_44_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_44_), .C(_37_), .Y(_45_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_40_), .C(_45_), .Y(w_C_10_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_40_), .Y(_46_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_46_), .Y(_47_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_48_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_48_), .Y(_49_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_49_), .C(_45_), .Y(_50_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .C(_50_), .Y(_51_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_51_), .Y(w_C_11_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .Y(_52_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add1[11]), .Y(_53_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_53_), .Y(_54_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_54_), .Y(_55_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_56_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_56_), .Y(_57_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_58_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_58_), .Y(_59_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_59_), .C(_50_), .Y(_60_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_55_), .Y(_61_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_61_), .Y(w_C_12_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_62_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_62_), .Y(_63_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_63_), .C(_60_), .Y(_64_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .C(_64_), .Y(_65_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_65_), .Y(w_C_13_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .Y(_66_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(i_add1[13]), .Y(_67_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_67_), .Y(_68_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_68_), .Y(_69_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_70_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_70_), .Y(_71_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_72_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_72_), .Y(_73_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_73_), .C(_64_), .Y(_74_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_69_), .Y(_75_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_75_), .Y(w_C_14_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_76_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_76_), .Y(_77_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_77_), .C(_74_), .Y(_78_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .C(_78_), .Y(_79_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_79_), .Y(w_C_15_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .Y(_80_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add1[15]), .Y(_81_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_81_), .Y(_82_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_82_), .Y(_83_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_84_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_84_), .Y(_85_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_86_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_86_), .Y(_87_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_87_), .C(_78_), .Y(_88_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_83_), .Y(_89_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_89_), .Y(w_C_16_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_90_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_90_), .Y(_91_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_91_), .C(_88_), .Y(_92_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .C(_92_), .Y(_93_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_93_), .Y(w_C_17_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .Y(_94_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add1[17]), .Y(_95_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_95_), .Y(_96_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_96_), .Y(_97_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_98_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_98_), .Y(_99_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_100_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(_100_), .Y(_101_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_101_), .C(_92_), .Y(_102_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_97_), .Y(_103_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_103_), .Y(w_C_18_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_104_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(_104_), .Y(_105_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_105_), .C(_102_), .Y(_106_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .C(_106_), .Y(_107_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_107_), .Y(w_C_19_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .Y(_108_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add1[19]), .Y(_109_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_109_), .Y(_110_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_110_), .Y(_111_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_112_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_112_), .Y(_113_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_114_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(_114_), .Y(_115_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_115_), .C(_106_), .Y(_116_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_111_), .Y(_117_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_117_), .Y(w_C_20_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_118_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_118_), .Y(_119_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_119_), .C(_116_), .Y(_120_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .C(_120_), .Y(_121_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_121_), .Y(w_C_21_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .Y(_122_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add1[21]), .Y(_123_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_123_), .Y(_124_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_124_), .Y(_125_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_126_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_126_), .Y(_127_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_128_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(_128_), .Y(_129_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_129_), .C(_120_), .Y(_130_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_125_), .Y(_131_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(_131_), .Y(w_C_22_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_132_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(_132_), .Y(_133_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_133_), .C(_130_), .Y(_134_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .C(_134_), .Y(_135_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(_135_), .Y(w_C_23_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .Y(_136_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add1[23]), .Y(_137_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_137_), .Y(_138_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(_138_), .Y(_139_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_140_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_140_), .Y(_141_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_142_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_142_), .Y(_143_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_143_), .C(_134_), .Y(_144_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_139_), .Y(_145_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(_145_), .Y(w_C_24_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_146_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(_146_), .Y(_147_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_147_), .C(_144_), .Y(_148_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .C(_148_), .Y(_149_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(_149_), .Y(w_C_25_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .Y(_150_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(i_add1[25]), .Y(_151_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_151_), .Y(_152_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(_152_), .Y(_153_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_154_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(_154_), .Y(_155_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_156_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(_156_), .Y(_157_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_157_), .C(_148_), .Y(_158_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_153_), .Y(_159_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(_159_), .Y(w_C_26_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_160_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(_160_), .Y(_161_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_161_), .C(_158_), .Y(_162_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .C(_162_), .Y(_163_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_163_), .Y(w_C_27_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .Y(_164_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(i_add1[27]), .Y(_165_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_165_), .Y(_166_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_166_), .Y(_167_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[26]), .B(i_add1[26]), .Y(_168_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(_168_), .Y(_169_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[27]), .B(i_add1[27]), .Y(_170_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_170_), .Y(_171_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_171_), .C(_162_), .Y(_172_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_167_), .Y(_173_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(_173_), .Y(w_C_28_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_174_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(_174_), .Y(_175_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_175_), .C(_172_), .Y(_176_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .C(_176_), .Y(_177_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(_177_), .Y(w_C_29_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .Y(_178_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(i_add1[29]), .Y(_179_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_179_), .Y(_180_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(_180_), .Y(_181_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[28]), .B(i_add1[28]), .Y(_182_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(_182_), .Y(_183_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[29]), .B(i_add1[29]), .Y(_184_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(_184_), .Y(_185_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_185_), .C(_176_), .Y(_186_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_181_), .Y(_187_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(_187_), .Y(w_C_30_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_188_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(_188_), .Y(_189_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_189_), .C(_186_), .Y(_190_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .C(_190_), .Y(_191_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(_191_), .Y(w_C_31_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_192_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[31]), .B(i_add1[31]), .Y(_193_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_191_), .C(_192_), .Y(w_C_32_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_194_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[30]), .B(i_add1[30]), .Y(_195_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(_195_), .Y(_196_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(_193_), .Y(_197_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_197_), .C(_190_), .Y(_198_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[32]), .B(i_add1[32]), .Y(_199_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(_199_), .C(_198_), .Y(_200_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_194_), .Y(w_C_33_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .Y(_201_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(i_add1[33]), .Y(_202_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_202_), .Y(_203_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_203_), .C(_200_), .Y(_204_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_201_), .B(_202_), .C(_204_), .Y(w_C_34_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .Y(_205_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(i_add1[34]), .Y(_206_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .C(w_C_34_), .Y(_207_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_206_), .C(_207_), .Y(w_C_35_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .Y(_208_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(i_add1[35]), .Y(_209_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_209_), .Y(_210_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(w_C_35_), .B(_210_), .Y(_211_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[35]), .B(i_add1[35]), .C(_211_), .Y(_212_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(_212_), .Y(w_C_36_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_213_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[36]), .B(i_add1[36]), .Y(_214_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_212_), .C(_213_), .Y(w_C_37_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_215_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(_214_), .Y(_216_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(_210_), .Y(_217_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_206_), .Y(_218_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[33]), .B(i_add1[33]), .Y(_219_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[34]), .B(i_add1[34]), .Y(_220_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_220_), .C(_204_), .Y(_221_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_209_), .Y(_222_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(_222_), .C(_221_), .Y(_223_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_213_), .C(_223_), .Y(_224_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(i_add2[37]), .B(i_add1[37]), .Y(_225_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_225_), .C(_224_), .Y(_226_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_226_), .Y(w_C_38_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_227_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[38]), .B(i_add1[38]), .Y(_228_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_228_), .C(_226_), .Y(_229_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_227_), .Y(w_C_39_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_230_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(i_add2[39]), .B(i_add1[39]), .Y(_231_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_231_), .C(_229_), .Y(_232_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_232_), .Y(w_C_40_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_233__0_), .Y(o_result[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_233__1_), .Y(o_result[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_233__2_), .Y(o_result[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_233__3_), .Y(o_result[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_233__4_), .Y(o_result[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_233__5_), .Y(o_result[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_233__6_), .Y(o_result[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_233__7_), .Y(o_result[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_233__8_), .Y(o_result[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_233__9_), .Y(o_result[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_233__10_), .Y(o_result[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_233__11_), .Y(o_result[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_233__12_), .Y(o_result[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_233__13_), .Y(o_result[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_233__14_), .Y(o_result[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_233__15_), .Y(o_result[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_233__16_), .Y(o_result[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_233__17_), .Y(o_result[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_233__18_), .Y(o_result[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_233__19_), .Y(o_result[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_233__20_), .Y(o_result[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_233__21_), .Y(o_result[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_233__22_), .Y(o_result[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_233__23_), .Y(o_result[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_233__24_), .Y(o_result[24]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_233__25_), .Y(o_result[25]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_233__26_), .Y(o_result[26]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_233__27_), .Y(o_result[27]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_233__28_), .Y(o_result[28]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_233__29_), .Y(o_result[29]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_233__30_), .Y(o_result[30]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_233__31_), .Y(o_result[31]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_233__32_), .Y(o_result[32]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_233__33_), .Y(o_result[33]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_233__34_), .Y(o_result[34]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_233__35_), .Y(o_result[35]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_233__36_), .Y(o_result[36]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_233__37_), .Y(o_result[37]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_233__38_), .Y(o_result[38]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_233__39_), .Y(o_result[39]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(w_C_40_), .Y(o_result[40]) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(w_C_4_), .Y(_237_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_238_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_239_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_239_), .C(_238_), .Y(_240_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_234_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[4]), .B(i_add1[4]), .Y(_235_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_235_), .C(w_C_4_), .Y(_236_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_240_), .Y(_233__4_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(w_C_5_), .Y(_244_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_245_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_246_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_246_), .C(_245_), .Y(_247_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_241_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[5]), .B(i_add1[5]), .Y(_242_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_242_), .C(w_C_5_), .Y(_243_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_247_), .Y(_233__5_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(w_C_6_), .Y(_251_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_252_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_253_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_251_), .B(_253_), .C(_252_), .Y(_254_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_248_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[6]), .B(i_add1[6]), .Y(_249_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_249_), .C(w_C_6_), .Y(_250_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_254_), .Y(_233__6_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(w_C_7_), .Y(_258_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_259_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_260_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_260_), .C(_259_), .Y(_261_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_255_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(i_add2[7]), .B(i_add1[7]), .Y(_256_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_256_), .C(w_C_7_), .Y(_257_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_261_), .Y(_233__7_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(w_C_8_), .Y(_265_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_266_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_267_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_267_), .C(_266_), .Y(_268_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_262_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(i_add2[8]), .B(i_add1[8]), .Y(_263_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_263_), .C(w_C_8_), .Y(_264_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_268_), .Y(_233__8_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(w_C_9_), .Y(_272_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_273_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_274_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_272_), .B(_274_), .C(_273_), .Y(_275_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_269_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(i_add2[9]), .B(i_add1[9]), .Y(_270_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_270_), .C(w_C_9_), .Y(_271_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_275_), .Y(_233__9_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(w_C_10_), .Y(_279_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_280_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_281_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_279_), .B(_281_), .C(_280_), .Y(_282_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_276_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(i_add2[10]), .B(i_add1[10]), .Y(_277_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_277_), .C(w_C_10_), .Y(_278_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_282_), .Y(_233__10_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(w_C_11_), .Y(_286_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_287_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_288_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_288_), .C(_287_), .Y(_289_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_283_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(i_add2[11]), .B(i_add1[11]), .Y(_284_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_283_), .B(_284_), .C(w_C_11_), .Y(_285_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_289_), .Y(_233__11_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(w_C_12_), .Y(_293_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_294_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_295_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_295_), .C(_294_), .Y(_296_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_290_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(i_add2[12]), .B(i_add1[12]), .Y(_291_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_291_), .C(w_C_12_), .Y(_292_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_292_), .B(_296_), .Y(_233__12_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(w_C_13_), .Y(_300_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_301_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_302_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_302_), .C(_301_), .Y(_303_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_297_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(i_add2[13]), .B(i_add1[13]), .Y(_298_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_298_), .C(w_C_13_), .Y(_299_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_303_), .Y(_233__13_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(w_C_14_), .Y(_307_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_308_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_309_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_309_), .C(_308_), .Y(_310_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_304_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(i_add2[14]), .B(i_add1[14]), .Y(_305_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_305_), .C(w_C_14_), .Y(_306_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_310_), .Y(_233__14_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(w_C_15_), .Y(_314_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_315_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_316_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_316_), .C(_315_), .Y(_317_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_311_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(i_add2[15]), .B(i_add1[15]), .Y(_312_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_312_), .C(w_C_15_), .Y(_313_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_317_), .Y(_233__15_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(w_C_16_), .Y(_321_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_322_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_323_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_323_), .C(_322_), .Y(_324_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_318_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(i_add2[16]), .B(i_add1[16]), .Y(_319_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_319_), .C(w_C_16_), .Y(_320_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_324_), .Y(_233__16_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(w_C_17_), .Y(_328_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_329_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_330_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_330_), .C(_329_), .Y(_331_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_325_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(i_add2[17]), .B(i_add1[17]), .Y(_326_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_325_), .B(_326_), .C(w_C_17_), .Y(_327_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_331_), .Y(_233__17_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(w_C_18_), .Y(_335_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_336_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_337_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_335_), .B(_337_), .C(_336_), .Y(_338_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_332_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(i_add2[18]), .B(i_add1[18]), .Y(_333_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_333_), .C(w_C_18_), .Y(_334_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_338_), .Y(_233__18_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(w_C_19_), .Y(_342_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_343_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_344_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_344_), .C(_343_), .Y(_345_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_339_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(i_add2[19]), .B(i_add1[19]), .Y(_340_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_340_), .C(w_C_19_), .Y(_341_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_345_), .Y(_233__19_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(w_C_20_), .Y(_349_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_350_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_351_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_351_), .C(_350_), .Y(_352_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_346_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(i_add2[20]), .B(i_add1[20]), .Y(_347_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_347_), .C(w_C_20_), .Y(_348_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_352_), .Y(_233__20_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(w_C_21_), .Y(_356_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_357_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_358_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_358_), .C(_357_), .Y(_359_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_353_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(i_add2[21]), .B(i_add1[21]), .Y(_354_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_354_), .C(w_C_21_), .Y(_355_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_359_), .Y(_233__21_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(w_C_22_), .Y(_363_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_364_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_365_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_365_), .C(_364_), .Y(_366_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_360_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(i_add2[22]), .B(i_add1[22]), .Y(_361_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_361_), .C(w_C_22_), .Y(_362_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_366_), .Y(_233__22_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(w_C_23_), .Y(_370_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_371_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_372_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_372_), .C(_371_), .Y(_373_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_367_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(i_add2[23]), .B(i_add1[23]), .Y(_368_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_368_), .C(w_C_23_), .Y(_369_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_373_), .Y(_233__23_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(w_C_24_), .Y(_377_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_378_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_379_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_379_), .C(_378_), .Y(_380_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_374_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(i_add2[24]), .B(i_add1[24]), .Y(_375_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_375_), .C(w_C_24_), .Y(_376_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_380_), .Y(_233__24_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(w_C_25_), .Y(_384_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_385_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(i_add2[25]), .B(i_add1[25]), .Y(_386_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_386_), .C(_385_), .Y(_387_) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(w_C_40_), .Y(_233__40_) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(w_C_0_) );
endmodule
